module conv12_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [1024-1:0] input_act,
    output logic [1024-1:0] output_act,
    output logic ready
);

logic [1024-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];
logic [7:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[519:512];
logic [7:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[527:520];
logic [7:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[535:528];
logic [7:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[543:536];
logic [7:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[551:544];
logic [7:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[559:552];
logic [7:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[567:560];
logic [7:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[575:568];
logic [7:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[583:576];
logic [7:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[591:584];
logic [7:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[599:592];
logic [7:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[607:600];
logic [7:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[615:608];
logic [7:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[623:616];
logic [7:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[631:624];
logic [7:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[639:632];
logic [7:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[647:640];
logic [7:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[655:648];
logic [7:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[663:656];
logic [7:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[671:664];
logic [7:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[679:672];
logic [7:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[687:680];
logic [7:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[695:688];
logic [7:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[703:696];
logic [7:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[711:704];
logic [7:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[719:712];
logic [7:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[727:720];
logic [7:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[735:728];
logic [7:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[743:736];
logic [7:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[751:744];
logic [7:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[759:752];
logic [7:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[767:760];
logic [7:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[775:768];
logic [7:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[783:776];
logic [7:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[791:784];
logic [7:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[799:792];
logic [7:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[807:800];
logic [7:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[815:808];
logic [7:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[823:816];
logic [7:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[831:824];
logic [7:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[839:832];
logic [7:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[847:840];
logic [7:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[855:848];
logic [7:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[863:856];
logic [7:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[871:864];
logic [7:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[879:872];
logic [7:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[887:880];
logic [7:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[895:888];
logic [7:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[903:896];
logic [7:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[911:904];
logic [7:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[919:912];
logic [7:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[927:920];
logic [7:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[935:928];
logic [7:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[943:936];
logic [7:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[951:944];
logic [7:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[959:952];
logic [7:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[967:960];
logic [7:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[975:968];
logic [7:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[983:976];
logic [7:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[991:984];
logic [7:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[999:992];
logic [7:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[1007:1000];
logic [7:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[1015:1008];
logic [7:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[1023:1016];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 15'sd 9028) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4477) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18666) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4310) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3223) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25341) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16069) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11562) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32099) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32410) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21951) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13983) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10526) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29220) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23726) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29380) * $signed(input_fmap_21[7:0]) +
	( 11'sd 578) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28172) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5902) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4330) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20966) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14056) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30882) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15238) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32466) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23396) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15215) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15246) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30054) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26178) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11452) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7084) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27349) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8618) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28898) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23072) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17267) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8452) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26169) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30623) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12044) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28594) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18489) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17484) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16657) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30022) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4553) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12404) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4841) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31256) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15976) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27195) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5911) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7482) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9884) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1528) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30982) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1701) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17812) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17644) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15075) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32676) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9300) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15281) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19894) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1571) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25779) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22924) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20341) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1712) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32078) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22482) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5550) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30328) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29066) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23454) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22063) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29132) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25264) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4417) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2372) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11092) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17728) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25630) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23797) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13416) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13747) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2490) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8841) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26875) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18628) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3751) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16756) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22506) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1819) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10967) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22145) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17651) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14122) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26697) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9562) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30884) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15889) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9064) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18287) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7628) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30990) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6446) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21206) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24056) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 15'sd 10815) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10162) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16165) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5063) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15797) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22344) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17284) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27309) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31857) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16752) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1393) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13299) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21731) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13399) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10890) * $signed(input_fmap_14[7:0]) +
	( 13'sd 4065) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8483) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14318) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13377) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26916) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11492) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7974) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13066) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27294) * $signed(input_fmap_25[7:0]) +
	( 10'sd 269) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19335) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32245) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31334) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31597) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11547) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5669) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15949) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15759) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8600) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26930) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14225) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9565) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2832) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22589) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24672) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12084) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19736) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8171) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13470) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22885) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32744) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4185) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21089) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3473) * $signed(input_fmap_53[7:0]) +
	( 10'sd 264) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31566) * $signed(input_fmap_55[7:0]) +
	( 11'sd 891) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15988) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19735) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4856) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2526) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5639) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26262) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3969) * $signed(input_fmap_63[7:0]) +
	( 14'sd 8056) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1252) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14667) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22276) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27145) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8536) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28948) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30052) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28636) * $signed(input_fmap_75[7:0]) +
	( 8'sd 102) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3440) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17971) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25750) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31929) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28101) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19884) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19883) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26143) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23981) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30050) * $signed(input_fmap_89[7:0]) +
	( 9'sd 236) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24900) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17628) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5569) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28637) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12272) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9278) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26771) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32138) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2965) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13992) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5321) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30094) * $signed(input_fmap_103[7:0]) +
	( 14'sd 8146) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7111) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32455) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28017) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21830) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8631) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10126) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22732) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12077) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6654) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25971) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8585) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17917) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10065) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31942) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10723) * $signed(input_fmap_120[7:0]) +
	( 11'sd 970) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1841) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3331) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6088) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3285) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19587) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23070) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 16'sd 32583) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7266) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17904) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14646) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8473) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24483) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7478) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14510) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2538) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26743) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1228) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22204) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3295) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22270) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17425) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9200) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15196) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24067) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6847) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2881) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26768) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15809) * $signed(input_fmap_25[7:0]) +
	( 10'sd 403) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1673) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19036) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23616) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23828) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19108) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24728) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24392) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14140) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15543) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17528) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30108) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20777) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24968) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29101) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25685) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32055) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24345) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5906) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20030) * $signed(input_fmap_49[7:0]) +
	( 11'sd 886) * $signed(input_fmap_50[7:0]) +
	( 11'sd 871) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29029) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12098) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25729) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6136) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32183) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30072) * $signed(input_fmap_57[7:0]) +
	( 11'sd 658) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17455) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6032) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2597) * $signed(input_fmap_61[7:0]) +
	( 8'sd 111) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21345) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26823) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29038) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17889) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1664) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8627) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26918) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16994) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19453) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24586) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30236) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30315) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30183) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12031) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29229) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7929) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12032) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6789) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21959) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30265) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31129) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17410) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12032) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7897) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18046) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8284) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8210) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24215) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21870) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13517) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15338) * $signed(input_fmap_94[7:0]) +
	( 9'sd 233) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24657) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30883) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22313) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12138) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12054) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13868) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32335) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10985) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11394) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18758) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9145) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19572) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6762) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32468) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30254) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18348) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2403) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12281) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6328) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17921) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8635) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11230) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1616) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5529) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23290) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4198) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8493) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30849) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13143) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14638) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6389) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 16'sd 32557) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31460) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14942) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18615) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27060) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26479) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23523) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31882) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17275) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14523) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4411) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26519) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3379) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17509) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7432) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19598) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24057) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8611) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17588) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1481) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8537) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2829) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21627) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23772) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3527) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9772) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8595) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9630) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5474) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7739) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26095) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26704) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32039) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32040) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13544) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24488) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26423) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15529) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15146) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31623) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10469) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5642) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17469) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21809) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27796) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22629) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11710) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28907) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19369) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2942) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1411) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21121) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27567) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32464) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20988) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16555) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32620) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19908) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5203) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19586) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10301) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25988) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32133) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21649) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16067) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29451) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24517) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2134) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8916) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5562) * $signed(input_fmap_82[7:0]) +
	( 8'sd 126) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15673) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11510) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17267) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11524) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16639) * $signed(input_fmap_89[7:0]) +
	( 13'sd 4078) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11495) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11202) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2896) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23014) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23385) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8990) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28044) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5295) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11018) * $signed(input_fmap_100[7:0]) +
	( 10'sd 472) * $signed(input_fmap_101[7:0]) +
	( 11'sd 554) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15504) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21050) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1617) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24223) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3425) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3996) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22130) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22462) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11593) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27129) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32047) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10105) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31759) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2792) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7397) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25661) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25587) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12564) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20643) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14633) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18477) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23013) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26138) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 16'sd 31906) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28261) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3638) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3422) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17371) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19790) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6447) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8397) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9127) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21314) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27151) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21178) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13151) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21931) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12259) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32648) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7402) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19441) * $signed(input_fmap_18[7:0]) +
	( 11'sd 682) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29328) * $signed(input_fmap_20[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17226) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19711) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13896) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3658) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22563) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28421) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17778) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27971) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25124) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24434) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31588) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25929) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9830) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7427) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23604) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1455) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3108) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21985) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27818) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30721) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2392) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19066) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29903) * $signed(input_fmap_48[7:0]) +
	( 13'sd 4027) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7366) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17478) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5917) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27563) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7326) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20113) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20161) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23123) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17972) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17362) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20579) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8193) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31631) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2158) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10480) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19995) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12780) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30060) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10524) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32625) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31474) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29690) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18634) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17178) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11829) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3754) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2962) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27605) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13741) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27365) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27695) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27352) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8830) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23329) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16264) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14763) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9461) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13292) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24311) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10822) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15133) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19012) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14389) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7261) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21279) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21591) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9757) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6623) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25247) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26440) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18808) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31362) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18415) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25598) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27109) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10274) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25676) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22536) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13617) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15950) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22480) * $signed(input_fmap_117[7:0]) +
	( 10'sd 504) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22350) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7905) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15620) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5997) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19380) * $signed(input_fmap_125[7:0]) +
	( 11'sd 896) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19031) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 16'sd 30431) * $signed(input_fmap_0[7:0]) +
	( 6'sd 19) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7383) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17710) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12513) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4152) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15982) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27272) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5127) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21692) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7820) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12101) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9756) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26654) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18886) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5824) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28646) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18052) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28956) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13921) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15146) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20426) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8655) * $signed(input_fmap_28[7:0]) +
	( 11'sd 672) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7445) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11133) * $signed(input_fmap_31[7:0]) +
	( 11'sd 856) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27491) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15387) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19542) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32082) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25078) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10978) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6210) * $signed(input_fmap_40[7:0]) +
	( 11'sd 848) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11868) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7407) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20696) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32020) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3919) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3434) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16629) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4415) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26630) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4278) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24088) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19891) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31109) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9161) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14217) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6381) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11787) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21257) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12822) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26370) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10812) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23645) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19963) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29000) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28885) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18685) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16962) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2837) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9742) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6310) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22788) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5461) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4793) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2615) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31784) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10855) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8142) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32759) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15140) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9020) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28858) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2585) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31495) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6872) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32632) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14623) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23886) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9110) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7126) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11673) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5956) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6862) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28854) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32380) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12600) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13789) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27887) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4520) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32741) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13250) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7428) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19651) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32514) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24916) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12868) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31197) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13516) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2594) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6886) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26071) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14436) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14510) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29620) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32237) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3775) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20297) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32171) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14069) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4659) * $signed(input_fmap_123[7:0]) +
	( 15'sd 16119) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1473) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1508) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 15'sd 9535) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24820) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12507) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23847) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7181) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17571) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8704) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31983) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28419) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10347) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10617) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23753) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21082) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10072) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29842) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21936) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19761) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22951) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30733) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7672) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26394) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1804) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11449) * $signed(input_fmap_28[7:0]) +
	( 10'sd 458) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13344) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22798) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32591) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10064) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12518) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5071) * $signed(input_fmap_36[7:0]) +
	( 10'sd 334) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11493) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23012) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27476) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2789) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12120) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27344) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10674) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17313) * $signed(input_fmap_47[7:0]) +
	( 9'sd 248) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6748) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3461) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10266) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2533) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12417) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6377) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28368) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13924) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9358) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22152) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18451) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23470) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21001) * $signed(input_fmap_62[7:0]) +
	( 7'sd 45) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14504) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26850) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24219) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3904) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22160) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17684) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7992) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30754) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1910) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25531) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22387) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5224) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15838) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18583) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32243) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32665) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22482) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14328) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29360) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28272) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11938) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21779) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3232) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2742) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14601) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19445) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30513) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28648) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28402) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30416) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13537) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19118) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26968) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29796) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13625) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26264) * $signed(input_fmap_100[7:0]) +
	( 11'sd 620) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31639) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27583) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16066) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6074) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21118) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25665) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30763) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_109[7:0]) +
	( 11'sd 877) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14862) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25724) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12924) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4844) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13446) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31284) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2885) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13730) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10934) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25413) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14473) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26955) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25037) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1130) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 16'sd 29319) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28196) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23533) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3098) * $signed(input_fmap_3[7:0]) +
	( 11'sd 760) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12773) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15690) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10539) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6846) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20957) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28601) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21268) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24211) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6956) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8896) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20809) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31670) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3493) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27772) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14799) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7301) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4745) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4407) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21401) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12471) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20545) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9189) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5666) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6519) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7498) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26760) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22934) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12647) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21473) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24326) * $signed(input_fmap_36[7:0]) +
	( 14'sd 8116) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7787) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13741) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22025) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17462) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21200) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25228) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16344) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3569) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22179) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27805) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18658) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10286) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19857) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1793) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18399) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2518) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24838) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7359) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16139) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5892) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4840) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13500) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23342) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30486) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3765) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26625) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17729) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6220) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22699) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30926) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17654) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3930) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2801) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23711) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11942) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9636) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25918) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24750) * $signed(input_fmap_84[7:0]) +
	( 11'sd 822) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6352) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14658) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27075) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25426) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29464) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19778) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16819) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6836) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1743) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14696) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17446) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2870) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5543) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16152) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31418) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22435) * $signed(input_fmap_102[7:0]) +
	( 11'sd 557) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3243) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28333) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_106[7:0]) +
	( 10'sd 478) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25355) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28927) * $signed(input_fmap_109[7:0]) +
	( 11'sd 888) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29617) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17762) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5268) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16449) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26879) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5919) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3782) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30160) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11326) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17235) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10641) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26256) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3320) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 14'sd 4767) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25338) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17172) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27032) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28123) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26056) * $signed(input_fmap_5[7:0]) +
	( 11'sd 828) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10093) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3820) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14584) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21248) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17792) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32392) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1182) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4737) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10215) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14025) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5138) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4815) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5612) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11215) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15433) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20851) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32081) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17989) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22273) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5579) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5113) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24835) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28027) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29508) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4514) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5745) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29239) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30854) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1540) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20557) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5156) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21275) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25944) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15137) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17456) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26155) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11375) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21389) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24905) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20131) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8685) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32188) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18628) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17441) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11382) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9233) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12273) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4270) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30790) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24402) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8810) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15627) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31395) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29172) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31189) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6426) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16861) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31928) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3505) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12053) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_80[7:0]) +
	( 11'sd 621) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28326) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26817) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27860) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20547) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5682) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13577) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3002) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8634) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21941) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14416) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25485) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28428) * $signed(input_fmap_94[7:0]) +
	( 8'sd 106) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4832) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29545) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3037) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6649) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28119) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31101) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13074) * $signed(input_fmap_102[7:0]) +
	( 10'sd 505) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17434) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8701) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13487) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12202) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29481) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31877) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28842) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27076) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8682) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11218) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5855) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8243) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12358) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18887) * $signed(input_fmap_120[7:0]) +
	( 14'sd 8064) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22149) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22443) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18359) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23131) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1767) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 16'sd 22510) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23857) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9398) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13824) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1078) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11023) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2339) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2973) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24664) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26395) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31300) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17659) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10640) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29988) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5931) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4931) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9472) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30335) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7870) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15794) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29260) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16735) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30630) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26734) * $signed(input_fmap_26[7:0]) +
	( 8'sd 99) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31193) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24884) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10914) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17500) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12289) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13235) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15602) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18590) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21500) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5679) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1181) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18888) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10575) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10014) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4434) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16504) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13965) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12158) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1818) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1330) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27606) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15697) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25756) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16679) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5060) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21589) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26172) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6261) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24731) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2209) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30987) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20237) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25865) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26713) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10959) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15471) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8285) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7601) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26711) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32387) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8050) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22631) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6325) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24359) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23986) * $signed(input_fmap_77[7:0]) +
	( 10'sd 411) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26908) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1513) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27122) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7210) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32606) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22359) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5214) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31594) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5502) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17234) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4796) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1242) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25331) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_92[7:0]) +
	( 10'sd 453) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1647) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6282) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19178) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29018) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10263) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6527) * $signed(input_fmap_101[7:0]) +
	( 10'sd 463) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24430) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18718) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12116) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16883) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28438) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27635) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10162) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2626) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18350) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29851) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7670) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1686) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17753) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8652) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12324) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2203) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8311) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4571) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17652) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28018) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16277) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4466) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28235) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 16'sd 25450) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25141) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6276) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28948) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5023) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11511) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14693) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31174) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32000) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5017) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12937) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5592) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18631) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13183) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25108) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32161) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18413) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28905) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29535) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29143) * $signed(input_fmap_20[7:0]) +
	( 11'sd 759) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6529) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4640) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2516) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5838) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7967) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9209) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26995) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9704) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9013) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18402) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32393) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7571) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5964) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7287) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15895) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24092) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28687) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10826) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11812) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9309) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11419) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24240) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4138) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4528) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3545) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9091) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26579) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8684) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5121) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29869) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23012) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31850) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16943) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27092) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4821) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5011) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5436) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29976) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6131) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3922) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17630) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28501) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21338) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4273) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19888) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19822) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25752) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2907) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14742) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31415) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13431) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22813) * $signed(input_fmap_83[7:0]) +
	( 10'sd 284) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28635) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9874) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6406) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3844) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18609) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28196) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10974) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24433) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3784) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7149) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13037) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4752) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25130) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29548) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3162) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32728) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25798) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25288) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27387) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19781) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22883) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8594) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19496) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30938) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28182) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21157) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16359) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4168) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31107) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2262) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14168) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21886) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7814) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20871) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26017) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4716) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25070) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21778) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31065) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31919) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 15'sd 13011) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24389) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27517) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26020) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14321) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16572) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32551) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31279) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19946) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2312) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12977) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31395) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11342) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30672) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16294) * $signed(input_fmap_14[7:0]) +
	( 11'sd 828) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13940) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22205) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27869) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11335) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12642) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10920) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26974) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15461) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14789) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10266) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19934) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12697) * $signed(input_fmap_30[7:0]) +
	( 10'sd 276) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9993) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13185) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10363) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17269) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25360) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31800) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4544) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11290) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5398) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24828) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32231) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18573) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21839) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32462) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11192) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1733) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31501) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27436) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6774) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30637) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3646) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10603) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27285) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19917) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2083) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3033) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2512) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16590) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5133) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13991) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16919) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1414) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15358) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21500) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11450) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5619) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31050) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16272) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31776) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20569) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18413) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32501) * $signed(input_fmap_80[7:0]) +
	( 10'sd 502) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22113) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29814) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19634) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6464) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26604) * $signed(input_fmap_88[7:0]) +
	( 9'sd 181) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12437) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13387) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20667) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25770) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25837) * $signed(input_fmap_95[7:0]) +
	( 11'sd 567) * $signed(input_fmap_96[7:0]) +
	( 10'sd 507) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1246) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7893) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3501) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3832) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27361) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20297) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28630) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29773) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6452) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8687) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11029) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29602) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30835) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2611) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7111) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7650) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22649) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5515) * $signed(input_fmap_118[7:0]) +
	( 14'sd 8036) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21119) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6156) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22326) * $signed(input_fmap_122[7:0]) +
	( 2'sd 1) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25477) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14217) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 10'sd 401) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17009) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7881) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15166) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30569) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14264) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22344) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7469) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13728) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28655) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18255) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26987) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19705) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14967) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9132) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23298) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19606) * $signed(input_fmap_17[7:0]) +
	( 11'sd 926) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14513) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18591) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24539) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19665) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5551) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7033) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14121) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16914) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18477) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23218) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16995) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29841) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6564) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9984) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6991) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30398) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16676) * $signed(input_fmap_35[7:0]) +
	( 11'sd 547) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11982) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17198) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1492) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27523) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29007) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6958) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22025) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3500) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30171) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3723) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1090) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22599) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4903) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22049) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32403) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31104) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31312) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26627) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26684) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29513) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23233) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8714) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23496) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21187) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14352) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5675) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4720) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17624) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3083) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18085) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17933) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7504) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30898) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20678) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25406) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25333) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20648) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13223) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18695) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6198) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13341) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12260) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14046) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19734) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28704) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5245) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31962) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15047) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3297) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29112) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26667) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30156) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27698) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26067) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24297) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17928) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30669) * $signed(input_fmap_99[7:0]) +
	( 11'sd 1019) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9470) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16964) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3896) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5353) * $signed(input_fmap_104[7:0]) +
	( 11'sd 955) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2537) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9260) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1576) * $signed(input_fmap_109[7:0]) +
	( 9'sd 195) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27858) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30120) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31985) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27164) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16992) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_117[7:0]) +
	( 13'sd 4073) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_119[7:0]) +
	( 14'sd 8133) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31553) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18942) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23568) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29919) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1894) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27904) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3924) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 15'sd 10417) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8261) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13864) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17275) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25051) * $signed(input_fmap_8[7:0]) +
	( 8'sd 101) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23058) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21138) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28497) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16455) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10366) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8799) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19759) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27179) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8567) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6471) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12193) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13889) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30264) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13801) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15255) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12042) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31872) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12099) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31641) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3436) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8219) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28358) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25815) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10522) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1526) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13274) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6751) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23146) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26761) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1182) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13551) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11360) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31246) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19736) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26717) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31241) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3329) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12628) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6226) * $signed(input_fmap_53[7:0]) +
	( 10'sd 326) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14592) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9123) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26655) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1718) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19402) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30589) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24617) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3989) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17923) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24464) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28622) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7357) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13531) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9022) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6289) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31160) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13783) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29607) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23102) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6055) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12733) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23345) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30075) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4924) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18590) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13528) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20390) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2420) * $signed(input_fmap_84[7:0]) +
	( 11'sd 977) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21143) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7892) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32424) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9713) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31965) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23109) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29575) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19736) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21404) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22428) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13650) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20587) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25308) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13675) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2884) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3049) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21518) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21700) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17069) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18982) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27987) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3028) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30396) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21644) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2898) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22218) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3113) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6832) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8418) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25218) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12754) * $signed(input_fmap_122[7:0]) +
	( 10'sd 271) * $signed(input_fmap_123[7:0]) +
	( 15'sd 16322) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32645) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 12'sd 1500) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21608) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18026) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20611) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4597) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2909) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12309) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20419) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5610) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6321) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2466) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21041) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29258) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10747) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13288) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5364) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10147) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7697) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9582) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3377) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19234) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19143) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1715) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18921) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5506) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7303) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21864) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27011) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2073) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8333) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17678) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4933) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18305) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15713) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7928) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28377) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29707) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9984) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4126) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16290) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1642) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9065) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14001) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21583) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8912) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21205) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21818) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25105) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11043) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23492) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30659) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21878) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32628) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13258) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28060) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30875) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21056) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11683) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7607) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30646) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3049) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26633) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12228) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16354) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15006) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16942) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2438) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19377) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32078) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8143) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25075) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1955) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28626) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15984) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22768) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2450) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32508) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26959) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16614) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7544) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3329) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12011) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14315) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21973) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18460) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31821) * $signed(input_fmap_100[7:0]) +
	( 9'sd 180) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29373) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2139) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15436) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22232) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22726) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18180) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16907) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16842) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9682) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14915) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25467) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18114) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22432) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11217) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9302) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15307) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19533) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5298) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28878) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17709) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15868) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11622) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 16'sd 26373) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21320) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3666) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7978) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24820) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26291) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30095) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14556) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17912) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8206) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14240) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7552) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5443) * $signed(input_fmap_13[7:0]) +
	( 11'sd 626) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30739) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18790) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21866) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25478) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1370) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28203) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11831) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31257) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9649) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24256) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31889) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14576) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11517) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16628) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30058) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18036) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14086) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17332) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25939) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3793) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21787) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2742) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25782) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24060) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11030) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24686) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13993) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13031) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3467) * $signed(input_fmap_47[7:0]) +
	( 6'sd 28) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7570) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7079) * $signed(input_fmap_50[7:0]) +
	( 14'sd 8169) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8969) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5975) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25103) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7861) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32653) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10475) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13831) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18888) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23450) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6230) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28146) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20167) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19456) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9742) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29517) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32401) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_71[7:0]) +
	( 8'sd 78) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4616) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31371) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10559) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3250) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12290) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24613) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19029) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2818) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13199) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11880) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16117) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31249) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5269) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30342) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1413) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7019) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26608) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8261) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26614) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14555) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17766) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23918) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30503) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1773) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3084) * $signed(input_fmap_98[7:0]) +
	( 11'sd 758) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10869) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2053) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5020) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10744) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29409) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2359) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15784) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4832) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16283) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22861) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12655) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11049) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9397) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25732) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15231) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32200) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28716) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1987) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19966) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15170) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31056) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32757) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8945) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11990) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6443) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 15'sd 9072) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20566) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27081) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21246) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11531) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17126) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22523) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29714) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19909) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6133) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6265) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19998) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9656) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25070) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29625) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23259) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31601) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20511) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5673) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13938) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26758) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21128) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7546) * $signed(input_fmap_28[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5851) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13138) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15663) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4366) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18092) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3769) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14996) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21133) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10171) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12362) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20479) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11777) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26436) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29507) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10304) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22493) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6721) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12489) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13302) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5485) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27197) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22591) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4193) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12263) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1695) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1390) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25951) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25561) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7757) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32564) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5536) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20596) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14406) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25668) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6475) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19340) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22318) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25335) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20859) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19628) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20654) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13024) * $signed(input_fmap_72[7:0]) +
	( 13'sd 4068) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1894) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2510) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31917) * $signed(input_fmap_76[7:0]) +
	( 8'sd 87) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21131) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9293) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28955) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1072) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17143) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31497) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23842) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4755) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13951) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6072) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28319) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14765) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19270) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27352) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3823) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31825) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12328) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5834) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24080) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21333) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5685) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3415) * $signed(input_fmap_99[7:0]) +
	( 9'sd 195) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20423) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21685) * $signed(input_fmap_104[7:0]) +
	( 11'sd 595) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28874) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16261) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4855) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17388) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14168) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27037) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14565) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19034) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20100) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11541) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18826) * $signed(input_fmap_119[7:0]) +
	( 9'sd 180) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11933) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10417) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17382) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15162) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28376) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 16'sd 19080) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30010) * $signed(input_fmap_2[7:0]) +
	( 15'sd 16098) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28122) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29060) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29147) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27742) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2422) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14355) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25475) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7751) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1237) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14622) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20681) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14946) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12470) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27290) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24019) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15481) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5281) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1403) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4732) * $signed(input_fmap_25[7:0]) +
	( 14'sd 8115) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14745) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27088) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8712) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28543) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3529) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19026) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3405) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9064) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29895) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11841) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27943) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25946) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18358) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3339) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18506) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24558) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13284) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9519) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10353) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22306) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17727) * $signed(input_fmap_49[7:0]) +
	( 11'sd 621) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18108) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13888) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25680) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13369) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12306) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9356) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20671) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10094) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15735) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13222) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24297) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27865) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1998) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21930) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14818) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1851) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7118) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25262) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18651) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21834) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11690) * $signed(input_fmap_71[7:0]) +
	( 10'sd 273) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2384) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7795) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7347) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9296) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9371) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12421) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12765) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3883) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25029) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3137) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28235) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6539) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26252) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26796) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25879) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23893) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31556) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12158) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2821) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28005) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22156) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14472) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2937) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20608) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1848) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_105[7:0]) +
	( 10'sd 320) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29154) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25269) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7004) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13554) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20206) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19803) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13727) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30937) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29108) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13703) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14708) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13130) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5996) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30511) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31236) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26956) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32457) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24838) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9852) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27217) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 16'sd 21042) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17674) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31258) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11540) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15607) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5051) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25431) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22225) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14400) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23853) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10898) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13811) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3032) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2317) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30258) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5170) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16079) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29431) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28734) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28561) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12759) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23363) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10739) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18717) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20947) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5387) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30766) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27403) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22980) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7934) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17854) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1251) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25738) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22763) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8997) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28553) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2271) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17981) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11138) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16749) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8034) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12653) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6044) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9875) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4181) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9603) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32154) * $signed(input_fmap_54[7:0]) +
	( 8'sd 109) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28212) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24916) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12112) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31314) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13065) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23291) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4531) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30313) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22321) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16203) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1839) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25954) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6857) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29058) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19024) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18724) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6257) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16322) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32520) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26353) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16533) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26600) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26647) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12865) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18316) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19394) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12062) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4661) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1207) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4533) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_92[7:0]) +
	( 10'sd 259) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7751) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9123) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26346) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3618) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13624) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7211) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26091) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8643) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5527) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28883) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27593) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17734) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11501) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27786) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5023) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5892) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26656) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5949) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9809) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23988) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23470) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17025) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28447) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5256) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9909) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20734) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 16'sd 23776) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15748) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15313) * $signed(input_fmap_2[7:0]) +
	( 14'sd 8165) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11909) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25149) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15891) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23779) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19073) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24008) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20655) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10493) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8325) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2572) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15642) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16840) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1432) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21329) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7549) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23984) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14968) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10470) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7311) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24059) * $signed(input_fmap_29[7:0]) +
	( 8'sd 122) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15986) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30774) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_33[7:0]) +
	( 10'sd 329) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10664) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8990) * $signed(input_fmap_36[7:0]) +
	( 11'sd 613) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29029) * $signed(input_fmap_39[7:0]) +
	( 14'sd 8085) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19820) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10279) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9852) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7227) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24944) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23102) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7813) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3504) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7928) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1586) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8776) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8503) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31740) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2145) * $signed(input_fmap_54[7:0]) +
	( 9'sd 189) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30728) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32158) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20395) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32498) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25309) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28400) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28705) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2466) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29786) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24501) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21000) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6730) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22118) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14316) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15661) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11016) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9040) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30362) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19398) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6463) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5144) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26795) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1949) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4622) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16976) * $signed(input_fmap_83[7:0]) +
	( 11'sd 915) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32122) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16995) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7680) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19920) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29233) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5034) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17961) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10572) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13532) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13667) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1235) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18418) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25933) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5756) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3701) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7514) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2870) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20956) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14001) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11734) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11507) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26546) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19768) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3155) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10216) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18199) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19975) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24440) * $signed(input_fmap_114[7:0]) +
	( 7'sd 62) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23078) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10091) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29937) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13028) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32465) * $signed(input_fmap_121[7:0]) +
	( 11'sd 733) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32366) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25798) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12204) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5676) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24607) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 14'sd 6572) * $signed(input_fmap_0[7:0]) +
	( 11'sd 761) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26452) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29199) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15600) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16028) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6889) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29677) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10350) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29193) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19935) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20681) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32446) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9348) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23737) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19559) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19338) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32182) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19106) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11486) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18298) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9935) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30276) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17096) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4280) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13924) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5525) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7017) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17084) * $signed(input_fmap_32[7:0]) +
	( 11'sd 981) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6026) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17558) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21026) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3883) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1672) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3692) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30105) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13775) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18623) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7307) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30565) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6665) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15815) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20738) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23168) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19511) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18707) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29060) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17712) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9417) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26550) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15556) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12999) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14411) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8639) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25995) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2191) * $signed(input_fmap_62[7:0]) +
	( 11'sd 1023) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21723) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29854) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16614) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25167) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24661) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32114) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26018) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28036) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19599) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29841) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31525) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21291) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25656) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21948) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2478) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21712) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31225) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30573) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10332) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1197) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3426) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8533) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27205) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16812) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18703) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29887) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4448) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20523) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27257) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32086) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32358) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30040) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19528) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7934) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_106[7:0]) +
	( 8'sd 103) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25432) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23613) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9734) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14420) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23261) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11567) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8435) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22799) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16722) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23586) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1373) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17794) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1189) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4925) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15771) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12865) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13608) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4542) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 15'sd 11075) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24120) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16321) * $signed(input_fmap_2[7:0]) +
	( 11'sd 1017) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31467) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29190) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14197) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24907) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28415) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23702) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24923) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30254) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14960) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1444) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30640) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32195) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18397) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2727) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29470) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6113) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12523) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6353) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7030) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32154) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27669) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18950) * $signed(input_fmap_26[7:0]) +
	( 15'sd 16328) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29382) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19124) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18142) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31063) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1290) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25637) * $signed(input_fmap_34[7:0]) +
	( 11'sd 513) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2869) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6230) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2931) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3148) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16161) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14802) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13511) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13884) * $signed(input_fmap_43[7:0]) +
	( 9'sd 143) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28576) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20307) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31606) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3481) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2876) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17754) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3558) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15426) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28727) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28069) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27400) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23035) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7432) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2573) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20441) * $signed(input_fmap_60[7:0]) +
	( 10'sd 318) * $signed(input_fmap_61[7:0]) +
	( 10'sd 272) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20169) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9094) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3559) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19820) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3572) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29468) * $signed(input_fmap_69[7:0]) +
	( 10'sd 340) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31703) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20456) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25109) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13603) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24623) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2943) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24551) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25704) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31754) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16508) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29118) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_83[7:0]) +
	( 11'sd 710) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15448) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30870) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32032) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18098) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26413) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13297) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9658) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18007) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19075) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13197) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3999) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28663) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31482) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19408) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9452) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7643) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12168) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11008) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21706) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15989) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19159) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14721) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9289) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5915) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31148) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31369) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20362) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7148) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7881) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32513) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24774) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27362) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2261) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24555) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31914) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 15'sd 14819) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22879) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2935) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12475) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26696) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22404) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27741) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23236) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25251) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31872) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7541) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12218) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18089) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16914) * $signed(input_fmap_13[7:0]) +
	( 9'sd 227) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21265) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25470) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21764) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22538) * $signed(input_fmap_18[7:0]) +
	( 11'sd 1000) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8471) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23139) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4573) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21754) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18991) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20682) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18747) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31768) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29313) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5508) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31832) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4346) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12273) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5986) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1281) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28525) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5933) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24507) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19485) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26540) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21040) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14173) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8200) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4456) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15472) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18022) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29202) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19911) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25812) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3481) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23767) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20100) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27548) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23283) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6452) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27029) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8504) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31403) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17278) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20032) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30529) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4757) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29894) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16516) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7627) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9818) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30641) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28135) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7506) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24054) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21080) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5432) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20515) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32128) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14900) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1036) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20058) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8879) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11649) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21664) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16331) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28336) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8656) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5746) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17030) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32763) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21232) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11889) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1100) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30681) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30301) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16964) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14924) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21177) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14646) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15771) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5863) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8409) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22720) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28649) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13823) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28185) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29242) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14612) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3133) * $signed(input_fmap_115[7:0]) +
	( 11'sd 854) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25664) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15652) * $signed(input_fmap_118[7:0]) +
	( 11'sd 582) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8520) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23986) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_122[7:0]) +
	( 9'sd 167) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32700) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13012) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21038) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18079) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 16'sd 20813) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5390) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2215) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6069) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18086) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15851) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27012) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16026) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16615) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26184) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1918) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8951) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31165) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22611) * $signed(input_fmap_15[7:0]) +
	( 11'sd 974) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5658) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10528) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27631) * $signed(input_fmap_19[7:0]) +
	( 11'sd 843) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32627) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12897) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30496) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10280) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2327) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13947) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32504) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20985) * $signed(input_fmap_28[7:0]) +
	( 12'sd 2038) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1103) * $signed(input_fmap_30[7:0]) +
	( 6'sd 25) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18087) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24414) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21118) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30054) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5043) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19722) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17420) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29610) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12576) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6472) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19687) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4480) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18835) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30544) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6691) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2893) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1427) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9946) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22660) * $signed(input_fmap_55[7:0]) +
	( 11'sd 845) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22567) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5352) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4879) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7934) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15876) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10753) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30042) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25711) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1126) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15007) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1080) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3751) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29568) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13997) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12710) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26029) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12823) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24088) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12650) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9325) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28880) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28632) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11944) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30770) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12292) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14726) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12173) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9789) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30255) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3677) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7195) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1844) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11740) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23718) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12345) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25762) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4224) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25641) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30121) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28743) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25539) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16678) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28359) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26069) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5393) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7890) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29655) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16620) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31443) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13424) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7203) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14850) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24086) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15990) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25212) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20004) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27959) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30030) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5821) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5636) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1797) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1070) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 16'sd 29432) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9879) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13356) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18222) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30868) * $signed(input_fmap_4[7:0]) +
	( 10'sd 373) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18002) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7524) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5657) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4528) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1785) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31818) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14992) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28598) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7512) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2626) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12357) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19880) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29561) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26270) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29592) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28227) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31755) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14661) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1717) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28933) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28079) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11059) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7840) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13856) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20047) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18812) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20908) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3374) * $signed(input_fmap_39[7:0]) +
	( 10'sd 429) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9487) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1334) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1620) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8385) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31133) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27926) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1929) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24815) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30221) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32436) * $signed(input_fmap_51[7:0]) +
	( 10'sd 482) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25424) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31541) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_55[7:0]) +
	( 12'sd 2032) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18975) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28652) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8873) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5521) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12084) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28822) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7548) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13570) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9743) * $signed(input_fmap_65[7:0]) +
	( 9'sd 254) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32091) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19975) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24281) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29984) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16967) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11263) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28480) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15655) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23333) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25285) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28305) * $signed(input_fmap_78[7:0]) +
	( 13'sd 4074) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28365) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13097) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28626) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30930) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13291) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31235) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15705) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30331) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8587) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11019) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1046) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30753) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5211) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25448) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24064) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32215) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18915) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29160) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9315) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13474) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27762) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22436) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9567) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4661) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11944) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6235) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24327) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18878) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1096) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26410) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6399) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16708) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31702) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30944) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5963) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21607) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4312) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4756) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20280) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2990) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14267) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24712) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 14'sd 7989) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9333) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16976) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27734) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32080) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15150) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12359) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15403) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19507) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19428) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18261) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23244) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30935) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22360) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26085) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13957) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7156) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5561) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8315) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8331) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27026) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12869) * $signed(input_fmap_23[7:0]) +
	( 10'sd 459) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24884) * $signed(input_fmap_25[7:0]) +
	( 7'sd 37) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9322) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7693) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20083) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26178) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28265) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5076) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9863) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13035) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4823) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15718) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12982) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6717) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19656) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10649) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13315) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24171) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31583) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18340) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22966) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2610) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7479) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4545) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3746) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27339) * $signed(input_fmap_59[7:0]) +
	( 11'sd 957) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13321) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9463) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25937) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14712) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11412) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20074) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18437) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8432) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11147) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7042) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7809) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6566) * $signed(input_fmap_74[7:0]) +
	( 11'sd 526) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5850) * $signed(input_fmap_76[7:0]) +
	( 10'sd 266) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15399) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32330) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22786) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30471) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15844) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3983) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31025) * $signed(input_fmap_85[7:0]) +
	( 10'sd 334) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27598) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26886) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1220) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17126) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25523) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8884) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3259) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24715) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7609) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9515) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28237) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15153) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10221) * $signed(input_fmap_100[7:0]) +
	( 11'sd 740) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2134) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16366) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23662) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1574) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12954) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32648) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20030) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30085) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27185) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22415) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20909) * $signed(input_fmap_112[7:0]) +
	( 10'sd 374) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26947) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17721) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11459) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16315) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21354) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15884) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21340) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13731) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12497) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22618) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27354) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5962) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11952) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 13'sd 2969) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20832) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9717) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21625) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24879) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11795) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2832) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21012) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14351) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12941) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29202) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5814) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18578) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16020) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21848) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26832) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15379) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18932) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6033) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5026) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2621) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21908) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6494) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28144) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25928) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15681) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20983) * $signed(input_fmap_30[7:0]) +
	( 11'sd 546) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5320) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6112) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1663) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7294) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12323) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19528) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24517) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7715) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2140) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21010) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20442) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1785) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17268) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14072) * $signed(input_fmap_48[7:0]) +
	( 10'sd 476) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3599) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8888) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19841) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9718) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18440) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21986) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13778) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29794) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23659) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24263) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17835) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13675) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24266) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17814) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32538) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1595) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25331) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_67[7:0]) +
	( 13'sd 4062) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26908) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16222) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21569) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9011) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26953) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23082) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21214) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11916) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4596) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21523) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26732) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20149) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16524) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16138) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29783) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20702) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15960) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3383) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17451) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18440) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_90[7:0]) +
	( 5'sd 8) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12046) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17694) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14883) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26984) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11250) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7720) * $signed(input_fmap_98[7:0]) +
	( 10'sd 358) * $signed(input_fmap_99[7:0]) +
	( 11'sd 574) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18672) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3901) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21223) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22791) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21379) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3153) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5740) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19493) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24338) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5034) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31712) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4697) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29915) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11536) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23361) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20494) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18976) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3436) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20024) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22216) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10773) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20826) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3539) * $signed(input_fmap_123[7:0]) +
	( 11'sd 986) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19188) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4716) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 16'sd 32487) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17722) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19857) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22361) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18740) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15766) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20300) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26122) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27519) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18879) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18459) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29705) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13005) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29251) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5788) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14793) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27439) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22807) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9776) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21657) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3532) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15223) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21034) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6059) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6366) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31727) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6778) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32019) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10945) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6904) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30512) * $signed(input_fmap_34[7:0]) +
	( 10'sd 487) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17221) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14444) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1091) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22780) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1038) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26067) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26988) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25227) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27938) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19416) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10176) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13616) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20648) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19984) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28033) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30523) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17791) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29783) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17854) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15102) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28095) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4966) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17064) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2662) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1430) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23312) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4901) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31544) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2146) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15660) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2412) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26396) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25817) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2774) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16900) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29605) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25954) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5539) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28837) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1454) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28596) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11635) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26787) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9306) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20469) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20263) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10774) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14530) * $signed(input_fmap_88[7:0]) +
	( 14'sd 8064) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19240) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14479) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21697) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6279) * $signed(input_fmap_94[7:0]) +
	( 11'sd 568) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19474) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21498) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18214) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6469) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10316) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25299) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7772) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10724) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22518) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22405) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25341) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22409) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25256) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3744) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7997) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5523) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19549) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5854) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10443) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16149) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_119[7:0]) +
	( 14'sd 8143) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23854) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26031) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3895) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23784) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2823) * $signed(input_fmap_125[7:0]) +
	( 10'sd 288) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5204) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 15'sd 13166) * $signed(input_fmap_0[7:0]) +
	( 10'sd 468) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4885) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27411) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31411) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24791) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7822) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28224) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28406) * $signed(input_fmap_13[7:0]) +
	( 14'sd 8058) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26210) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22618) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12057) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6288) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3727) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11031) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11131) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10002) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9611) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9272) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16944) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13703) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10807) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23734) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14987) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22868) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22178) * $signed(input_fmap_33[7:0]) +
	( 11'sd 786) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6950) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4560) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3673) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4661) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13436) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28485) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26289) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10497) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14330) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23564) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23014) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7766) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15514) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31330) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12078) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32275) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21517) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13828) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23456) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12000) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18630) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30778) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11087) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16608) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5951) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6077) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1899) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20263) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17751) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31021) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25299) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11773) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10281) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27587) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20589) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13490) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11242) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1944) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25118) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24365) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9555) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8464) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19496) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21526) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12825) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18462) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11151) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20144) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14481) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30107) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16760) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7012) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17475) * $signed(input_fmap_93[7:0]) +
	( 7'sd 50) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30793) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12707) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1467) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16648) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1228) * $signed(input_fmap_100[7:0]) +
	( 13'sd 4078) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12005) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24099) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28174) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2558) * $signed(input_fmap_106[7:0]) +
	( 9'sd 201) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30479) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12416) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3150) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5567) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29884) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16888) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15405) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9145) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10890) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32009) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7571) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11608) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9746) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21356) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27565) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23793) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1727) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21560) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25492) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4655) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 13'sd 3716) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3609) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27894) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9112) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6698) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29461) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4650) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19806) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7176) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30486) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1783) * $signed(input_fmap_10[7:0]) +
	( 12'sd 2026) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28924) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19369) * $signed(input_fmap_13[7:0]) +
	( 11'sd 806) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23022) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11793) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17466) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24335) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3400) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27721) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6764) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3010) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25589) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8084) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21849) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6920) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21528) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5854) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28031) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31112) * $signed(input_fmap_32[7:0]) +
	( 13'sd 4050) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6557) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4813) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1319) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23873) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15618) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19588) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4364) * $signed(input_fmap_41[7:0]) +
	( 7'sd 50) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32315) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23463) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31980) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23896) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14504) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10523) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29070) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25815) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21499) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26695) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14426) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14297) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6839) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32288) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12205) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24080) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28295) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21736) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10959) * $signed(input_fmap_63[7:0]) +
	( 10'sd 325) * $signed(input_fmap_64[7:0]) +
	( 10'sd 448) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30078) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19202) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27248) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17163) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17897) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10247) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15457) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24583) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3665) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8122) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2610) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11282) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17061) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19182) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30968) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11356) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22133) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13157) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20745) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10330) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9300) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18417) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17871) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7229) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27473) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14733) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21649) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7844) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24670) * $signed(input_fmap_101[7:0]) +
	( 14'sd 8014) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25611) * $signed(input_fmap_103[7:0]) +
	( 10'sd 499) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25697) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29990) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15607) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8545) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15297) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30530) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24060) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7742) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2049) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11342) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10722) * $signed(input_fmap_116[7:0]) +
	( 10'sd 491) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27623) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22900) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11697) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15446) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4842) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5300) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1498) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 15'sd 13698) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7678) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31453) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27415) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30063) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29723) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30530) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2206) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23508) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31379) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28973) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17754) * $signed(input_fmap_11[7:0]) +
	( 11'sd 849) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15072) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28300) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2780) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15807) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1317) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6048) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19047) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24690) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3606) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17634) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25382) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28293) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14066) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28170) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28159) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30532) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12638) * $signed(input_fmap_30[7:0]) +
	( 8'sd 91) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19319) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20259) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11697) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5939) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12869) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29514) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22398) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21131) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27503) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3255) * $signed(input_fmap_43[7:0]) +
	( 11'sd 907) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11327) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6030) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5868) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30992) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6499) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27968) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6193) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20731) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24692) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8860) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28135) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13891) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22230) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16794) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5116) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6822) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6118) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23700) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17480) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23363) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19014) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19096) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14438) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4765) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15599) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29341) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10237) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31532) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14224) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10274) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28333) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12622) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30756) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3063) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21724) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25665) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23813) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24273) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1424) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5939) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28910) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23814) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23339) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28195) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12829) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29278) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3849) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26432) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19169) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29602) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25824) * $signed(input_fmap_104[7:0]) +
	( 10'sd 490) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6390) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4455) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10530) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21009) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30416) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4986) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27115) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9393) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6207) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2154) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14850) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1729) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14234) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29658) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12583) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20188) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13123) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25089) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7371) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22345) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 13'sd 3110) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12417) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21983) * $signed(input_fmap_3[7:0]) +
	( 11'sd 1009) * $signed(input_fmap_4[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25275) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25109) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31545) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9566) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18597) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31482) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11857) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7076) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24433) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12994) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31529) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14837) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1602) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19847) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30518) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30065) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4846) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28887) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14650) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11166) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9968) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27520) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1170) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4729) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32558) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32325) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32603) * $signed(input_fmap_37[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26609) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23717) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10910) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30251) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27997) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9947) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4782) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13607) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13864) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15011) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12431) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11699) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29382) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31417) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19957) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11617) * $signed(input_fmap_56[7:0]) +
	( 11'sd 772) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16636) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15402) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29431) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25640) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22633) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10351) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11781) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15676) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16713) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6211) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6002) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29536) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16647) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19720) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5844) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23246) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14320) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15183) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3888) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7731) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32277) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1522) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21711) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25515) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18284) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20410) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26264) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20390) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32100) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27740) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27599) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17315) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26352) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19701) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17123) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7426) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1685) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11616) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2155) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26462) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16130) * $signed(input_fmap_106[7:0]) +
	( 11'sd 548) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3379) * $signed(input_fmap_108[7:0]) +
	( 9'sd 183) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6196) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27586) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16975) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14230) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26535) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17370) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22684) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32495) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1449) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23657) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14441) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6630) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2758) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13256) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6374) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16713) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 14'sd 5279) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6170) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28517) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5093) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9738) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7234) * $signed(input_fmap_6[7:0]) +
	( 8'sd 110) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20485) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29885) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7497) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21526) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9838) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8388) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24592) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3705) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25398) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9353) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_21[7:0]) +
	( 10'sd 323) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30139) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20240) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26037) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9948) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7833) * $signed(input_fmap_27[7:0]) +
	( 14'sd 8132) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12472) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7723) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22651) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2868) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13585) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9276) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18871) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14559) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22945) * $signed(input_fmap_39[7:0]) +
	( 11'sd 899) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2585) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17999) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31405) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19488) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13292) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27042) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7050) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28734) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29014) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8847) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14995) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3119) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4345) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24096) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28564) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7199) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24075) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8539) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29432) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4709) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2611) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1128) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24730) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31676) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17516) * $signed(input_fmap_68[7:0]) +
	( 14'sd 8136) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8456) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3219) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3342) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25383) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28165) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6585) * $signed(input_fmap_75[7:0]) +
	( 11'sd 670) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18165) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1698) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8155) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10059) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25644) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9580) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3513) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25964) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3765) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6882) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6483) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25392) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13219) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14358) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29612) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31190) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26375) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18968) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8259) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15265) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21325) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28720) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24700) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27397) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27885) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14786) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10581) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27298) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14458) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11877) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23951) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22620) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14382) * $signed(input_fmap_115[7:0]) +
	( 11'sd 765) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18855) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27456) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21218) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29975) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24188) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25343) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28951) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18169) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13001) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9170) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16551) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 16'sd 22614) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1965) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10100) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22568) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24815) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16598) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8633) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9345) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12234) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14393) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7687) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27129) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2718) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32542) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15081) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6468) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28190) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31209) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21376) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24683) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1350) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3206) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28937) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2971) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7437) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3757) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14240) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26234) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32256) * $signed(input_fmap_30[7:0]) +
	( 11'sd 646) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25560) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26759) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27784) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6772) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17974) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14612) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28536) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9795) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20799) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22380) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14868) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5145) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11454) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1946) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19037) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1073) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20939) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26939) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20279) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22336) * $signed(input_fmap_52[7:0]) +
	( 13'sd 4032) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27746) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3265) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22151) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13980) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18156) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18960) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29908) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2781) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6272) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5133) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20698) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27635) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17266) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11860) * $signed(input_fmap_70[7:0]) +
	( 5'sd 15) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9158) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30889) * $signed(input_fmap_73[7:0]) +
	( 15'sd 16215) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23217) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20996) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24795) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1515) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14052) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9166) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21423) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21863) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24244) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26140) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11342) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20587) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11151) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12109) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21002) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6041) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2889) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16107) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22327) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13707) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11870) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24484) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27052) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8667) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16666) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2846) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22417) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3995) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12943) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4739) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32029) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10205) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30859) * $signed(input_fmap_108[7:0]) +
	( 11'sd 667) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31203) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18251) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18865) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6991) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27158) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10247) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24329) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29714) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9057) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32219) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31136) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25520) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25401) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20885) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4996) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29146) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 16'sd 22316) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17979) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22248) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22860) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7888) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2791) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27894) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8901) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14118) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9435) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2161) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31860) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22202) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27147) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6429) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24346) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4996) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22437) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10275) * $signed(input_fmap_23[7:0]) +
	( 7'sd 56) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19210) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23613) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21778) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15196) * $signed(input_fmap_28[7:0]) +
	( 12'sd 2044) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19072) * $signed(input_fmap_30[7:0]) +
	( 11'sd 705) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24229) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19225) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10105) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24993) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2721) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5902) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3091) * $signed(input_fmap_40[7:0]) +
	( 14'sd 8169) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10941) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11659) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25522) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16235) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3734) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11612) * $signed(input_fmap_47[7:0]) +
	( 11'sd 631) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26420) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4246) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27003) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13183) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25311) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6744) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20418) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13045) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9385) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24998) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7115) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27159) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14638) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8240) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11220) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18543) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31560) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13282) * $signed(input_fmap_66[7:0]) +
	( 11'sd 720) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29990) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11773) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13690) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11520) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29968) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26636) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17702) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24715) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21197) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23286) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21329) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7079) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22617) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27600) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17789) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16239) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26446) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4308) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15080) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28574) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6942) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3867) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27199) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8760) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19669) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18132) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19678) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8703) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7577) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23112) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8773) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13284) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24142) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15282) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18418) * $signed(input_fmap_107[7:0]) +
	( 11'sd 977) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9172) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7522) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9342) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21190) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31479) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14014) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17762) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25336) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7220) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9480) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29181) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30372) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19859) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17766) * $signed(input_fmap_123[7:0]) +
	( 14'sd 8058) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2524) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12287) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7882) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 16'sd 21003) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31937) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9263) * $signed(input_fmap_2[7:0]) +
	( 16'sd 32290) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6881) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22514) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16644) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6680) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2541) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17710) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24408) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7781) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14306) * $signed(input_fmap_12[7:0]) +
	( 13'sd 4015) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2795) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25387) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3150) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17725) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17997) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5278) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7098) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7947) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24717) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1601) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24912) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3636) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12768) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7711) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8764) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2894) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15872) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32380) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17337) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16632) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2162) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16458) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5184) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30444) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19687) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11234) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12121) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29937) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12453) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14829) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21915) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28952) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7402) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26249) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18406) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32395) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16433) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2939) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32587) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25054) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10941) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24325) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26624) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9261) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29704) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30291) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11911) * $signed(input_fmap_64[7:0]) +
	( 11'sd 676) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5139) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5660) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30126) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31496) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29458) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24697) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27344) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29053) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2511) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26001) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11921) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2461) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28870) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1685) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30341) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7405) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28791) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30330) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10219) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26963) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7120) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30014) * $signed(input_fmap_90[7:0]) +
	( 10'sd 317) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30781) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8703) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7325) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23580) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30894) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12974) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17910) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16001) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23293) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9451) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27293) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30389) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6991) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26743) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29601) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21760) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3679) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31372) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21664) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8877) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15644) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13356) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30657) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30187) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16980) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1237) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31384) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12539) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1637) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11669) * $signed(input_fmap_123[7:0]) +
	( 10'sd 264) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29275) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4963) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19714) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 16'sd 25567) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24893) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29322) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15441) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29824) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31229) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29727) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30077) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14358) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15821) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20476) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18285) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6188) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4264) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12091) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2283) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30730) * $signed(input_fmap_17[7:0]) +
	( 9'sd 167) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19179) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19304) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22096) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11196) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19325) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11625) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24081) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7543) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1554) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2672) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24985) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28986) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1942) * $signed(input_fmap_33[7:0]) +
	( 11'sd 743) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3351) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18334) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6872) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32129) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16530) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6679) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3394) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27808) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18063) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23144) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28849) * $signed(input_fmap_49[7:0]) +
	( 11'sd 705) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9232) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4264) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32438) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28741) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18673) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27614) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12399) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5838) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11962) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1207) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29087) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13032) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15127) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14058) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14436) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10579) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29259) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4647) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26965) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10008) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8406) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22644) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30612) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9117) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11514) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32619) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4121) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8999) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24582) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6622) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10368) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17053) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12768) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16903) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16793) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22170) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25787) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30994) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14367) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24957) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24295) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28929) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4832) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11194) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18416) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2492) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20363) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21722) * $signed(input_fmap_105[7:0]) +
	( 11'sd 808) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19965) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2780) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11286) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22907) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20978) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7369) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1999) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20840) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12954) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30116) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31651) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18051) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11333) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4606) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9838) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9139) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5225) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5789) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12668) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 11'sd 771) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4385) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2967) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17254) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29071) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27908) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12186) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12914) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12629) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1923) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27061) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27656) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5746) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4116) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8213) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3469) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7899) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21069) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17624) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20417) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20439) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12907) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30175) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21612) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30539) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27369) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14754) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15859) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18333) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16231) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19382) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7297) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20090) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11152) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25221) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_36[7:0]) +
	( 10'sd 379) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11491) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29798) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1588) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18573) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25246) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22971) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16830) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26418) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25752) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23605) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23093) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10555) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5870) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22871) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27950) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12385) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1456) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5215) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21216) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5202) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7486) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27538) * $signed(input_fmap_60[7:0]) +
	( 10'sd 334) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15904) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20698) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28267) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2825) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6746) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31531) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5598) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26879) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5545) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24990) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31512) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10482) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31009) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5289) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10903) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19001) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13354) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8702) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30518) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16670) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9930) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30855) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17512) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2442) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17669) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9406) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24421) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17952) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29931) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2927) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22406) * $signed(input_fmap_96[7:0]) +
	( 10'sd 425) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18722) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13937) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1873) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23372) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23430) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18710) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5747) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7943) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17315) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25636) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32629) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10158) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17116) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1505) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3806) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8435) * $signed(input_fmap_117[7:0]) +
	( 4'sd 7) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23146) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30439) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4340) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9309) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10873) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22692) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17336) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 14'sd 6548) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18635) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16274) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27005) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17114) * $signed(input_fmap_4[7:0]) +
	( 10'sd 328) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3230) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31383) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25885) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24552) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10245) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8890) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16195) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9248) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8911) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22943) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1840) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7679) * $signed(input_fmap_20[7:0]) +
	( 11'sd 843) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32477) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11956) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18333) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3666) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24562) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23419) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3756) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19855) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15791) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21090) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7723) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23162) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30669) * $signed(input_fmap_35[7:0]) +
	( 14'sd 8086) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13390) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6193) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28740) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26136) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32140) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12617) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15641) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18280) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3534) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25347) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23829) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16959) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23561) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12234) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5792) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11323) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11828) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7930) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11217) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2132) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22720) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28090) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15827) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26533) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6060) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23333) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19978) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11142) * $signed(input_fmap_67[7:0]) +
	( 11'sd 571) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20769) * $signed(input_fmap_69[7:0]) +
	( 12'sd 2006) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30007) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30016) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16053) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30996) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17279) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4586) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13096) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28292) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13855) * $signed(input_fmap_79[7:0]) +
	( 13'sd 4057) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11607) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10375) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2798) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32121) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19984) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20509) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27374) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2374) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11978) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15896) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13085) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27038) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32612) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10875) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20108) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5508) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9199) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2615) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8746) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5437) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27878) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20271) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19210) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25728) * $signed(input_fmap_113[7:0]) +
	( 11'sd 549) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5170) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20078) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28191) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1224) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5366) * $signed(input_fmap_119[7:0]) +
	( 14'sd 8182) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18337) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7511) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21157) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24299) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26436) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12647) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18762) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 15'sd 13455) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13339) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27752) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29933) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13406) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21711) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10856) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3005) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15724) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10294) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13591) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6917) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3243) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22758) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28892) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20667) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3051) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15413) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20237) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24731) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17753) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20386) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24907) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17591) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22351) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23588) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19479) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2838) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24378) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31483) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18473) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20191) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26915) * $signed(input_fmap_35[7:0]) +
	( 11'sd 661) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5229) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29207) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23004) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5532) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23516) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4508) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28667) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6495) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7467) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32199) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24765) * $signed(input_fmap_47[7:0]) +
	( 11'sd 968) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29558) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31406) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26251) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4618) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6805) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28468) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13317) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3503) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7680) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31547) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10686) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10284) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12154) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24498) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12140) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22513) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25401) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2138) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17322) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19734) * $signed(input_fmap_69[7:0]) +
	( 13'sd 4042) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2841) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7584) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20613) * $signed(input_fmap_77[7:0]) +
	( 13'sd 4028) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14656) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22550) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18680) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1470) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2758) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28048) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7725) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28421) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24415) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22717) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28423) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24944) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8130) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21935) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14933) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10266) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20292) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5679) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26068) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18498) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29760) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12289) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10702) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20139) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26261) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18117) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18014) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4290) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28976) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21296) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16394) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13381) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12178) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2284) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19613) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28431) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3881) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8640) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27409) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5166) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28077) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 16'sd 24833) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6697) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3355) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18165) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28398) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28446) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32742) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18326) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20089) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29434) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8510) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4370) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3865) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26191) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15477) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21555) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30899) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30825) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25691) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22875) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5774) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12409) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6848) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2584) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13352) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16234) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22333) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19525) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19354) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9097) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5022) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10776) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17116) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12715) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5882) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12696) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21923) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6324) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18073) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10026) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2704) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7548) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27979) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30256) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17447) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31689) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1777) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13641) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9734) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3761) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16132) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23772) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6470) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21061) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29494) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12505) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20522) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18892) * $signed(input_fmap_69[7:0]) +
	( 8'sd 79) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14616) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5925) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5765) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10169) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13316) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25046) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6732) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9053) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24057) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29330) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15530) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15998) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4135) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7646) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22504) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22717) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4340) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13079) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17185) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3378) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10429) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10423) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29254) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17664) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28975) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25561) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9733) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2671) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23880) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1634) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27618) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20802) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16247) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11789) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6452) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28812) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6035) * $signed(input_fmap_112[7:0]) +
	( 6'sd 24) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15076) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19628) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32554) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17550) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23306) * $signed(input_fmap_118[7:0]) +
	( 15'sd 16296) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11677) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13243) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29491) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8485) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9474) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26949) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26293) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 15'sd 10758) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31604) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12844) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22427) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32314) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30266) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21514) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30308) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23367) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17062) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3382) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4583) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20003) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1776) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28245) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10142) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14232) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2714) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10059) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16674) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15123) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5738) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30852) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8759) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20534) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22736) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16870) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31427) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5760) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1764) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15792) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9237) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23998) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21333) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15775) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1167) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20886) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11320) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26986) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1328) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16950) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19491) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31984) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30812) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29582) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15838) * $signed(input_fmap_52[7:0]) +
	( 12'sd 2000) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26359) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26273) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15519) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9465) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6936) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19783) * $signed(input_fmap_59[7:0]) +
	( 11'sd 1009) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24417) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12493) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24087) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4178) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9994) * $signed(input_fmap_66[7:0]) +
	( 11'sd 722) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16262) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24431) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9497) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3548) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20524) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31125) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29335) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3942) * $signed(input_fmap_76[7:0]) +
	( 11'sd 825) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16020) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12521) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28094) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28739) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9435) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26147) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14828) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3370) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7590) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2163) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29863) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8709) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_92[7:0]) +
	( 7'sd 36) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9600) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11124) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18605) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32122) * $signed(input_fmap_98[7:0]) +
	( 13'sd 4063) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32391) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18168) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25956) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30301) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5804) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25137) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2650) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26627) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1359) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7160) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16464) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32681) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28591) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28168) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20186) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29757) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9303) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29203) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5393) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15859) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15847) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19629) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21743) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26142) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 15'sd 9597) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6855) * $signed(input_fmap_1[7:0]) +
	( 14'sd 8124) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10310) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22559) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28894) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2941) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10335) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1509) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13127) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26541) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11026) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14039) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22831) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26367) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5599) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25308) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8222) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13875) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25369) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10710) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32244) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30726) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26264) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25554) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6126) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9413) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31235) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31473) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2976) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13684) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22054) * $signed(input_fmap_36[7:0]) +
	( 11'sd 589) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19584) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18430) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25756) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14665) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19809) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13595) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6784) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23846) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3105) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2896) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9926) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6589) * $signed(input_fmap_51[7:0]) +
	( 10'sd 267) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29496) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26038) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8978) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19330) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24596) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30257) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28108) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9600) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26677) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14028) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14900) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19651) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22192) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25053) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13905) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14946) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7451) * $signed(input_fmap_70[7:0]) +
	( 8'sd 114) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14076) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11671) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14157) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24019) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12798) * $signed(input_fmap_77[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28701) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27755) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32714) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2416) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6941) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10506) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7265) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_87[7:0]) +
	( 11'sd 1018) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12033) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28437) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21119) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5997) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12738) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18118) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24431) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7766) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14565) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1908) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23954) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2110) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21427) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12493) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18702) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20560) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31442) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20029) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8224) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15979) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30618) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15429) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20997) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26898) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28859) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22026) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26431) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32764) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26049) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23475) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3317) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29948) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17547) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17223) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32406) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8358) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8149) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 16'sd 29544) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17870) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1472) * $signed(input_fmap_2[7:0]) +
	( 11'sd 936) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1703) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5178) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10412) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2968) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28689) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32208) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10786) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29681) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2784) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24907) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19719) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8937) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24808) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3590) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1258) * $signed(input_fmap_19[7:0]) +
	( 14'sd 8034) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4132) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28437) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1265) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7955) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28023) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17732) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28092) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2695) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30231) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7398) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17518) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19840) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7877) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15026) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28446) * $signed(input_fmap_35[7:0]) +
	( 11'sd 562) * $signed(input_fmap_36[7:0]) +
	( 11'sd 785) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14040) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6119) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1331) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27361) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24093) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16607) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32210) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29000) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21501) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1842) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10298) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7571) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17714) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17342) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13831) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21890) * $signed(input_fmap_55[7:0]) +
	( 11'sd 834) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22440) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32503) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27765) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20292) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32016) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6754) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5237) * $signed(input_fmap_64[7:0]) +
	( 8'sd 126) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11632) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8463) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19524) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8711) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19261) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28434) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9559) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30052) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23141) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25762) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1133) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5385) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28827) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1219) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16900) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14924) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7860) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16784) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7500) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11217) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21092) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15783) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17233) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17340) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6198) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_92[7:0]) +
	( 11'sd 831) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14369) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18326) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1648) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25362) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17172) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31808) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16391) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19927) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15052) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19130) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12132) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4672) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27821) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5436) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13277) * $signed(input_fmap_111[7:0]) +
	( 12'sd 2036) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24773) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25916) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13357) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9289) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6957) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32231) * $signed(input_fmap_119[7:0]) +
	( 10'sd 301) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21725) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20193) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16217) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29758) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29112) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22475) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 15'sd 15421) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11379) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12891) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15777) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11463) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13954) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19842) * $signed(input_fmap_7[7:0]) +
	( 11'sd 938) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31457) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29020) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30670) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7623) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31807) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20418) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17320) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15491) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23694) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21822) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17022) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7211) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8217) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4704) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21282) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24813) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25212) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29869) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29002) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18294) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19912) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21363) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30592) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17377) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7345) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12542) * $signed(input_fmap_36[7:0]) +
	( 10'sd 499) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29689) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13832) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22145) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4675) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7551) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29202) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8999) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26356) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5215) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28490) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9806) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31636) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17985) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24990) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26021) * $signed(input_fmap_55[7:0]) +
	( 10'sd 413) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13795) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20283) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19773) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28338) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10568) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29405) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16494) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31523) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26464) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5241) * $signed(input_fmap_67[7:0]) +
	( 5'sd 9) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16663) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3182) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30587) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27935) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18324) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19716) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9472) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5466) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22442) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8206) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28731) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17086) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27879) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14490) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29850) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30734) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32408) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27150) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27558) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21907) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18301) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8212) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3772) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16846) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11159) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6678) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27589) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24093) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6733) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21827) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16594) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5656) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11891) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30358) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14623) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1305) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28637) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1522) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27502) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30110) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4533) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15213) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20329) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16159) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31521) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12075) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28714) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5203) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28046) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32145) * $signed(input_fmap_123[7:0]) +
	( 11'sd 806) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26648) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14676) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17190) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 14'sd 4407) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30525) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25378) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14254) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30416) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4576) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29309) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28419) * $signed(input_fmap_9[7:0]) +
	( 10'sd 303) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26592) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19828) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13728) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27043) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12102) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7969) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12265) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20470) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19029) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9493) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12613) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22827) * $signed(input_fmap_24[7:0]) +
	( 11'sd 765) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8365) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23017) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2815) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9643) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27879) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27437) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2918) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17831) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17914) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10179) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29432) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22606) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2600) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25823) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16218) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2230) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3904) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2288) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25466) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5301) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17623) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27811) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9632) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30187) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2245) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14772) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10269) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18851) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1025) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7251) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14172) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15214) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21098) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22412) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5202) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19634) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16347) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32650) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12238) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4398) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25036) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17246) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22805) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27741) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11529) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28990) * $signed(input_fmap_77[7:0]) +
	( 7'sd 54) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12070) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26453) * $signed(input_fmap_81[7:0]) +
	( 9'sd 212) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4714) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14984) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31811) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13828) * $signed(input_fmap_87[7:0]) +
	( 10'sd 343) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23273) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31589) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12228) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30877) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15908) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24323) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5480) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13878) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18464) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11053) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13562) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29675) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13823) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12166) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_105[7:0]) +
	( 14'sd 8172) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2471) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24561) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1823) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11648) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25817) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_112[7:0]) +
	( 10'sd 461) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32434) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29098) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22495) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19970) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17087) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25452) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12389) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20298) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5903) * $signed(input_fmap_123[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30084) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6856) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 16'sd 20166) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14188) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19342) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29845) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1065) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27461) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4221) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25085) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20224) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6102) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1557) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12643) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30492) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5947) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4952) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2409) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13871) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26272) * $signed(input_fmap_20[7:0]) +
	( 9'sd 254) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20197) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2114) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31686) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2103) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21531) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21088) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14951) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13144) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9878) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6764) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12918) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12628) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22256) * $signed(input_fmap_35[7:0]) +
	( 5'sd 15) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12796) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30299) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21750) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14447) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22324) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27197) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11709) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2969) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20737) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20053) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28399) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29505) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20719) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27968) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22772) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17728) * $signed(input_fmap_53[7:0]) +
	( 11'sd 994) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12438) * $signed(input_fmap_55[7:0]) +
	( 11'sd 563) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32299) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32134) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4899) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12405) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19557) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12672) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21372) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25767) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7302) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15380) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8780) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22917) * $signed(input_fmap_71[7:0]) +
	( 10'sd 289) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18946) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11581) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14958) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16236) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24740) * $signed(input_fmap_77[7:0]) +
	( 11'sd 725) * $signed(input_fmap_78[7:0]) +
	( 11'sd 589) * $signed(input_fmap_79[7:0]) +
	( 11'sd 666) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2091) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32346) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29606) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27416) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27515) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31083) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3217) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14677) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18899) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30131) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32477) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27033) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31446) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19954) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15361) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7863) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21773) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30335) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7938) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3919) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18528) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30425) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22220) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6282) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7676) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2136) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5147) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25650) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3831) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18567) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5212) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6998) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3048) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26631) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24124) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19822) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22466) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31322) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26249) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17686) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27654) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26505) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30573) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 14'sd 7205) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3772) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29268) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31982) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1965) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24249) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29559) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28872) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11416) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4161) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20080) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3864) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13756) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30780) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3639) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30057) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21996) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18766) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24915) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32325) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10384) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19158) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7431) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23767) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10157) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6904) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20226) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13794) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15709) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27753) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11236) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27799) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19489) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20111) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9761) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6793) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2394) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6466) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15641) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7459) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12667) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32531) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1834) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15437) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28663) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18704) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32526) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24363) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9525) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11290) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21332) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21249) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18760) * $signed(input_fmap_63[7:0]) +
	( 11'sd 770) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28929) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19688) * $signed(input_fmap_66[7:0]) +
	( 7'sd 62) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24658) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10371) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3779) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25465) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10257) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10943) * $signed(input_fmap_74[7:0]) +
	( 11'sd 687) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6024) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27871) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29598) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18753) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22551) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7500) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30926) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14392) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15242) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24066) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27868) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22735) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22220) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8904) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29798) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25796) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5840) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26626) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19268) * $signed(input_fmap_98[7:0]) +
	( 11'sd 806) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29315) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8304) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21335) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24067) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2218) * $signed(input_fmap_104[7:0]) +
	( 13'sd 4021) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25955) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31427) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9892) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21562) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10607) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1989) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18084) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24369) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20519) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2323) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26813) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4913) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25008) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31140) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4551) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29586) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27115) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18786) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 14'sd 5724) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7203) * $signed(input_fmap_1[7:0]) +
	( 13'sd 4047) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20019) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22473) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14327) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22900) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7285) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22111) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15141) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1584) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18514) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9319) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4522) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28168) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31532) * $signed(input_fmap_17[7:0]) +
	( 11'sd 565) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30009) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5343) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6156) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23401) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_23[7:0]) +
	( 10'sd 473) * $signed(input_fmap_24[7:0]) +
	( 10'sd 263) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17396) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12420) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14986) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1907) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26937) * $signed(input_fmap_32[7:0]) +
	( 10'sd 362) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26101) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8687) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16295) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9740) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1078) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13059) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16587) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21209) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21704) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1207) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7612) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7190) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31940) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22403) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6174) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31313) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23992) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14102) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30897) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7348) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28735) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1355) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14012) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23075) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20867) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21135) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7349) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15162) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31399) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13724) * $signed(input_fmap_66[7:0]) +
	( 9'sd 219) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12415) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18575) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2220) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16907) * $signed(input_fmap_71[7:0]) +
	( 9'sd 237) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25210) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8203) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28677) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24934) * $signed(input_fmap_76[7:0]) +
	( 10'sd 490) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21836) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25687) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2168) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19397) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26307) * $signed(input_fmap_83[7:0]) +
	( 13'sd 4023) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1175) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12476) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16319) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31414) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3581) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14564) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8818) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9870) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28679) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1141) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12886) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10901) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3256) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26368) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28679) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20903) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6364) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13694) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5059) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32497) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20343) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11315) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25184) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5885) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15815) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1766) * $signed(input_fmap_110[7:0]) +
	( 11'sd 809) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26964) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22171) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4159) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23958) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28888) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30676) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14740) * $signed(input_fmap_118[7:0]) +
	( 10'sd 488) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28478) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3727) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20040) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13316) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30358) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9272) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 16'sd 19972) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24828) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19850) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31900) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19084) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23490) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21033) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9757) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30735) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27877) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12052) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22173) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17690) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4171) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23400) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15134) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4469) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28973) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20874) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1474) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14152) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23493) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3323) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13045) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9522) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8844) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15072) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2396) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25045) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19412) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18074) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7444) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22119) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27771) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20758) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26224) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21141) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31875) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21442) * $signed(input_fmap_40[7:0]) +
	( 14'sd 8033) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28262) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23553) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20812) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15894) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27548) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28756) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14002) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21352) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2073) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27430) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21424) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20426) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9721) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23926) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22231) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29606) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21313) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17570) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22458) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11742) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2364) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13330) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22107) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12109) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6354) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25263) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29146) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7087) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26776) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1245) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27382) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10155) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6016) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17927) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18436) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6705) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3892) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19848) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13725) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17317) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4518) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14253) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20247) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3411) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11413) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18694) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7905) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29472) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12151) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5009) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28467) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22173) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31610) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4553) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31655) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14618) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20639) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2956) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12768) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27121) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6297) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17665) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29977) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5752) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23611) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1538) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24279) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22603) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9182) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21758) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27630) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9585) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20353) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23497) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18600) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18861) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 15'sd 10705) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6428) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5930) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25827) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8334) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10722) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13375) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30517) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11812) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19421) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19829) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7046) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7688) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23136) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14623) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32443) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13681) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7679) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26805) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1818) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15057) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10260) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24014) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15499) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23629) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26553) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23379) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23587) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17072) * $signed(input_fmap_30[7:0]) +
	( 10'sd 508) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12277) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32541) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28231) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2154) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7699) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28028) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8853) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4873) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1055) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29567) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18550) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15812) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26199) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22546) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32486) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24852) * $signed(input_fmap_50[7:0]) +
	( 10'sd 438) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3080) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9229) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10236) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26595) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23628) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9536) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10040) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21414) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11339) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2629) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32436) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9276) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30488) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12098) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32694) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26678) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22293) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22678) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32621) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3183) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10043) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16596) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16731) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31534) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29390) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32524) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15940) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22219) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24937) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18370) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23150) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10035) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28126) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14228) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8252) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22341) * $signed(input_fmap_96[7:0]) +
	( 14'sd 8053) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25573) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19336) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17144) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25870) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3534) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12687) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12422) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24075) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20501) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31924) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31858) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8900) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6623) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9377) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30053) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12903) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22957) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30710) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30157) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5709) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30610) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24800) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28972) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8975) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 16'sd 24637) * $signed(input_fmap_0[7:0]) +
	( 11'sd 1010) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6525) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24537) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18889) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32189) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25940) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23380) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3586) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20399) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15338) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15325) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16618) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29269) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9339) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6031) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31140) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10179) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23876) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9864) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7452) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30303) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16984) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23558) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2574) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12109) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21527) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11106) * $signed(input_fmap_30[7:0]) +
	( 11'sd 642) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8623) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15847) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17738) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2196) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9277) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29511) * $signed(input_fmap_37[7:0]) +
	( 14'sd 8158) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7868) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8617) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7182) * $signed(input_fmap_41[7:0]) +
	( 11'sd 912) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3380) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29895) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27518) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17875) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22461) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11216) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18176) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1423) * $signed(input_fmap_52[7:0]) +
	( 9'sd 152) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7505) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15229) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7990) * $signed(input_fmap_56[7:0]) +
	( 6'sd 22) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32548) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2350) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13709) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28929) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18975) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1770) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30958) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6490) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29051) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22913) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2399) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9719) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26712) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9166) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8505) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15457) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20720) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24604) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31346) * $signed(input_fmap_77[7:0]) +
	( 11'sd 559) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6613) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7050) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18735) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1405) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7677) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8328) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24466) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21948) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19438) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10176) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2893) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27592) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24231) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7714) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16324) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16817) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26509) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25772) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28994) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25411) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27776) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19441) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2974) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32596) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27410) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21746) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27855) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20138) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10344) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16380) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14853) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20514) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25053) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23532) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10754) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23562) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23649) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_122[7:0]) +
	( 10'sd 467) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19451) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14726) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13369) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 16'sd 21686) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17467) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9896) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13424) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18639) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19947) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28137) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15023) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28868) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30869) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7779) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26385) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8675) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20209) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23524) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10837) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13994) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32343) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26010) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7024) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25182) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20395) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8349) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23799) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14909) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31730) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19333) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21274) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9092) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26089) * $signed(input_fmap_33[7:0]) +
	( 10'sd 440) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30962) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24650) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16368) * $signed(input_fmap_37[7:0]) +
	( 8'sd 117) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10916) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25315) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27381) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14048) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29867) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5452) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5022) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16712) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16666) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21571) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3241) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32653) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23029) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13740) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5791) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22311) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10913) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23791) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32171) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22777) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28832) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17037) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6649) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29446) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14653) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3161) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11559) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24209) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18004) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9412) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6308) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31037) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6645) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22226) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23743) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27588) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9019) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19061) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26085) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6128) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5414) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17020) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8235) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29036) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28086) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13538) * $signed(input_fmap_87[7:0]) +
	( 11'sd 966) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21239) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32236) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18772) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29457) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10556) * $signed(input_fmap_94[7:0]) +
	( 11'sd 573) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5933) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1454) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21129) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29726) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20295) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24909) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12346) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5438) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21951) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29263) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25358) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29348) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8796) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17459) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12387) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6463) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23514) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15384) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12659) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11047) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25726) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26619) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12698) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2994) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10901) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4223) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24640) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24912) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22563) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 16'sd 22435) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1449) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9354) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2645) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14912) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20554) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2745) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11610) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26961) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12233) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31340) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12498) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20329) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19961) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24070) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32009) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9670) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22686) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23548) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21120) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10530) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12894) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15534) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8296) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1561) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13846) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3525) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24099) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30679) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15549) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17328) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15574) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24051) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24491) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12411) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21492) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29689) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29510) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2319) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27635) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5802) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10370) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28171) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18776) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31887) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18985) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2804) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17169) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21019) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30268) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7766) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4993) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29659) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1842) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19414) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15621) * $signed(input_fmap_73[7:0]) +
	( 10'sd 374) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20587) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29711) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5986) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3112) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16429) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28194) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18579) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27433) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18203) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13321) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9914) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7466) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23575) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12328) * $signed(input_fmap_92[7:0]) +
	( 11'sd 687) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13402) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21803) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16950) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23664) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7819) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1392) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11130) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23149) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3374) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22088) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31877) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19893) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25976) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26265) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13282) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16024) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17796) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31908) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21469) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3440) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18082) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7839) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_124[7:0]) +
	( 13'sd 4025) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4623) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3101) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 12'sd 1884) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1837) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24519) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17634) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11626) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17352) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15952) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8521) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3451) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29528) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28074) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23706) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17915) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24277) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10083) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20595) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31208) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19079) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11114) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27699) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7760) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25654) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24667) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11835) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30771) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23212) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22596) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7302) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9597) * $signed(input_fmap_29[7:0]) +
	( 11'sd 723) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18157) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20087) * $signed(input_fmap_32[7:0]) +
	( 13'sd 4092) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29726) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_35[7:0]) +
	( 9'sd 200) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30108) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13145) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12216) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11090) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3671) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1628) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11438) * $signed(input_fmap_44[7:0]) +
	( 14'sd 8172) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24657) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26598) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14310) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16844) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24813) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9932) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31488) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29820) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13028) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30906) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18002) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7724) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30242) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9226) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16446) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31561) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13324) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29787) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15043) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10055) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3207) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20751) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30087) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17534) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32541) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7227) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16146) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2708) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27098) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31910) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28197) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18677) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4701) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14827) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12149) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24588) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10986) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24976) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4411) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21349) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13417) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8921) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22208) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16649) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25439) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8483) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3540) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12489) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2480) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2104) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29052) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26588) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24022) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18966) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5091) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12099) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14328) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21005) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12845) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13607) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19886) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25444) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22345) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13641) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32193) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25351) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18710) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18410) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5275) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17391) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25123) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3986) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 14'sd 6544) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20264) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20563) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12773) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11139) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32192) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5485) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19040) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1559) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21669) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26977) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30107) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18844) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22513) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28218) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12889) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15408) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12341) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20106) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14523) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2103) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13338) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24755) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14231) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14732) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8684) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22879) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23430) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23177) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23180) * $signed(input_fmap_40[7:0]) +
	( 10'sd 503) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26702) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5451) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3089) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11808) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23021) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22452) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5851) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24805) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6674) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15093) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20957) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5690) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15179) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11497) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14855) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25670) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15824) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11774) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10585) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1389) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21203) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8599) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18264) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9246) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6329) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24503) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11528) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3180) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17774) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29338) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3057) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26224) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7188) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30219) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9715) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9653) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24551) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17937) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4688) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29303) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29962) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24791) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7923) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23369) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17051) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24085) * $signed(input_fmap_94[7:0]) +
	( 12'sd 2016) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9825) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22976) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26684) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3664) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7596) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3808) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31419) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7468) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3034) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7333) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11081) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12898) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32455) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6843) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13351) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13314) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1024) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26029) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9679) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10211) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21287) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27400) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5809) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5147) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32249) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12545) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5681) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9365) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21949) * $signed(input_fmap_126[7:0]) +
	( 10'sd 341) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 16'sd 26821) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13473) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6823) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25313) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23472) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9583) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5385) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27644) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15460) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7910) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25754) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24913) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15084) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4642) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28498) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_16[7:0]) +
	( 10'sd 308) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1258) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29566) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23274) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25827) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31553) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15734) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27850) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23942) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18630) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8324) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18440) * $signed(input_fmap_29[7:0]) +
	( 9'sd 177) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14883) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18548) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22013) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10040) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9139) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10980) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15279) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21522) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13255) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25437) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7698) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12558) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9315) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32761) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28667) * $signed(input_fmap_45[7:0]) +
	( 11'sd 761) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13714) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12638) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28828) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27145) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17297) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16993) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23651) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19045) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8765) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32172) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1073) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19343) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17254) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4413) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23835) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13552) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20355) * $signed(input_fmap_66[7:0]) +
	( 13'sd 4025) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4442) * $signed(input_fmap_68[7:0]) +
	( 11'sd 525) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30213) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31122) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26743) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24068) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16412) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25244) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15390) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11753) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12327) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18026) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10083) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14570) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24261) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27877) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29545) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6597) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2383) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29152) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30520) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22092) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19398) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1066) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10254) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2333) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18681) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26234) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27641) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22488) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5711) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8694) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8412) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2914) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5349) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24141) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23255) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3764) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20822) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3177) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10795) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32574) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13314) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24094) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15235) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11783) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26134) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7473) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7988) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10248) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13615) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1137) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6013) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 15'sd 14706) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12515) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14982) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27336) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27002) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13454) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10218) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1075) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31968) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22445) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8420) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4360) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10809) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7932) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27781) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31786) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25409) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22390) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5504) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11211) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5185) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9520) * $signed(input_fmap_24[7:0]) +
	( 10'sd 401) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7967) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22479) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27394) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7535) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6958) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32377) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28315) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31957) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20934) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5819) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21199) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30145) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30641) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15894) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11120) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13690) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21230) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1284) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15090) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15934) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12748) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16835) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19415) * $signed(input_fmap_52[7:0]) +
	( 11'sd 856) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31178) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26708) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23761) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10822) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27222) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26321) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23842) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4514) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8519) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22885) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16000) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24823) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29643) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31696) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1451) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11070) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17202) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29677) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20334) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24528) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17572) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23083) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6496) * $signed(input_fmap_79[7:0]) +
	( 11'sd 642) * $signed(input_fmap_80[7:0]) +
	( 9'sd 173) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14326) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26886) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32071) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1172) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17379) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26745) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22244) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19556) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23181) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28824) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15658) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16784) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6185) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31346) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7205) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28385) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21879) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4209) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12824) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1551) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14108) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6118) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20476) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3080) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15215) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26377) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8891) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3303) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22325) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21106) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10906) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29505) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7534) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25378) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7331) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9519) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8111) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30191) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16842) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7054) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23442) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3608) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 15'sd 12480) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32277) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22742) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15562) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10676) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5294) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31975) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5546) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9007) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8725) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22742) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21051) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2274) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15951) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7724) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31933) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17684) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11992) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23057) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14512) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13937) * $signed(input_fmap_22[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32467) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7577) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12504) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26956) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23644) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1460) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26642) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16344) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21082) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24915) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20831) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11325) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20982) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22225) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32737) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32116) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15245) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28488) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29693) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31514) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31758) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21568) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_50[7:0]) +
	( 11'sd 809) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8864) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15958) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27568) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29187) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10260) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20144) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18654) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25521) * $signed(input_fmap_61[7:0]) +
	( 11'sd 636) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26268) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24191) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21586) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29721) * $signed(input_fmap_67[7:0]) +
	( 10'sd 329) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1902) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27453) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25231) * $signed(input_fmap_71[7:0]) +
	( 9'sd 206) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11584) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30741) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16417) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23468) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21267) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28118) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13443) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27777) * $signed(input_fmap_87[7:0]) +
	( 11'sd 800) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5208) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1674) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18906) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16651) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26997) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19085) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15127) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19040) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19646) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21990) * $signed(input_fmap_98[7:0]) +
	( 11'sd 711) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27514) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28083) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24279) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15798) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8571) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25306) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25656) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3753) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32651) * $signed(input_fmap_112[7:0]) +
	( 11'sd 852) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18677) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20792) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15714) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16465) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6941) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1487) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19338) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12939) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2755) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9386) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28308) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 16'sd 16792) * $signed(input_fmap_0[7:0]) +
	( 14'sd 8064) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18614) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10810) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25486) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13501) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14439) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4156) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7950) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1444) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16340) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16385) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13943) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19355) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20694) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7519) * $signed(input_fmap_17[7:0]) +
	( 11'sd 564) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14928) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29428) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28371) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32550) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10770) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31320) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30585) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23505) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7329) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23177) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19433) * $signed(input_fmap_30[7:0]) +
	( 9'sd 236) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10617) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24677) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13136) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12290) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9565) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10053) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14360) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2281) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31354) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32238) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1045) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9788) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21209) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22495) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23999) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9151) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3182) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32336) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11777) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5254) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18334) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12927) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29657) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4121) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20155) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14493) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11794) * $signed(input_fmap_61[7:0]) +
	( 14'sd 8144) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13682) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9363) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12909) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25934) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28186) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18047) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29816) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26580) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9257) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25667) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13013) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13960) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4542) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19916) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7529) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3717) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29539) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29105) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3615) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12913) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11370) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16531) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13529) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10784) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27015) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27943) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2257) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27320) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18966) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16820) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31415) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28981) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2963) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3415) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22420) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29220) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13402) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16521) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7698) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27758) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10302) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3260) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10793) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14643) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4121) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24171) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7044) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30101) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22290) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1981) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26239) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12970) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31865) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19910) * $signed(input_fmap_125[7:0]) +
	( 10'sd 458) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3951) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 16'sd 30642) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7200) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2880) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14942) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3875) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23408) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17931) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5600) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18712) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16228) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17886) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5262) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27902) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32731) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27542) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31068) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14755) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17078) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12518) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26344) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21737) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23975) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31129) * $signed(input_fmap_26[7:0]) +
	( 7'sd 46) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19688) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20425) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19666) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17544) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2624) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19298) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19176) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13649) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8692) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26800) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8885) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2879) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26405) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2675) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9173) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28298) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12903) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6645) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19548) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5488) * $signed(input_fmap_50[7:0]) +
	( 10'sd 269) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8624) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19849) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17024) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9672) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22088) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16139) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_58[7:0]) +
	( 11'sd 1008) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3842) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22347) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11548) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9789) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13512) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3563) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26269) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16668) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2313) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19517) * $signed(input_fmap_69[7:0]) +
	( 11'sd 825) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32566) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6048) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8723) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24125) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26050) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1899) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26100) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5389) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19635) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1763) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10628) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25778) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27727) * $signed(input_fmap_86[7:0]) +
	( 10'sd 295) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26217) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6396) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21227) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5296) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18012) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22490) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22276) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25762) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12592) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7606) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21241) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16285) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9556) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14173) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23908) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21834) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21563) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17024) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27535) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24578) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17015) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32084) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13785) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11346) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11655) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8619) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13799) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20285) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2313) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24997) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29880) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9287) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16997) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25597) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 16'sd 24450) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24772) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18036) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13706) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14364) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15462) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6005) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12570) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15327) * $signed(input_fmap_8[7:0]) +
	( 10'sd 440) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5658) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6273) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19915) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10341) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4463) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1315) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18842) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17783) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18387) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25531) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8814) * $signed(input_fmap_22[7:0]) +
	( 9'sd 131) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23547) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18841) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20121) * $signed(input_fmap_27[7:0]) +
	( 11'sd 1013) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25466) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10607) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3434) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28113) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10832) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6983) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8551) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25350) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16561) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16945) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20360) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6016) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22034) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7359) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23230) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3737) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21867) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10800) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22439) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30867) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8924) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8791) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2518) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29320) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17157) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13939) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2534) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5030) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4521) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16735) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25518) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16538) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11910) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21247) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29069) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6363) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32714) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25277) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27840) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14916) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10384) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20506) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30393) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13011) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32458) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12818) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2332) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5301) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22700) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2719) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23111) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22915) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12667) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17922) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13858) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5095) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26396) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19510) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12151) * $signed(input_fmap_98[7:0]) +
	( 11'sd 703) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13596) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11780) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10550) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16101) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24149) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9040) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2280) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25592) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2401) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14933) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22157) * $signed(input_fmap_114[7:0]) +
	( 13'sd 4089) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10968) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3362) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24133) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15698) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10508) * $signed(input_fmap_122[7:0]) +
	( 11'sd 953) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18442) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7258) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24129) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22786) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 15'sd 12848) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8560) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20467) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27384) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30617) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1188) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16029) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26004) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22458) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3930) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18576) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15521) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10133) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12917) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2682) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6538) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14121) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4963) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4231) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31384) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11660) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13752) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5190) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25660) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25304) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14666) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29160) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24423) * $signed(input_fmap_34[7:0]) +
	( 11'sd 962) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18379) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10052) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20986) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29871) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8564) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12843) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24124) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8740) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29126) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10362) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10646) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7643) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20961) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4685) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12824) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12064) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8993) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19215) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29718) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16713) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11687) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19256) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1678) * $signed(input_fmap_65[7:0]) +
	( 9'sd 244) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23473) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15229) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22396) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21609) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14601) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4640) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31239) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3769) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3423) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27156) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22260) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10798) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5978) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18487) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7517) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18654) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17769) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16751) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6738) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30243) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6914) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11552) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22209) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13424) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17899) * $signed(input_fmap_93[7:0]) +
	( 11'sd 544) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24715) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15369) * $signed(input_fmap_97[7:0]) +
	( 11'sd 555) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29091) * $signed(input_fmap_99[7:0]) +
	( 11'sd 532) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25489) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3537) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10402) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1578) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28673) * $signed(input_fmap_105[7:0]) +
	( 11'sd 665) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15833) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9860) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18986) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10266) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1676) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25461) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6953) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2179) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11647) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10870) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30631) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14127) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14865) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2694) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20614) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9764) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15671) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31081) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9932) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 14'sd 6099) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12611) * $signed(input_fmap_1[7:0]) +
	( 11'sd 808) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32007) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30588) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9013) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6210) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1099) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28187) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25307) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15285) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13250) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7197) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22741) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29565) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1991) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1341) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13074) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2905) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23205) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14421) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4963) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30854) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25019) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3374) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13475) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12585) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14090) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21256) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6652) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30024) * $signed(input_fmap_37[7:0]) +
	( 14'sd 8112) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10980) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31075) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17992) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27267) * $signed(input_fmap_43[7:0]) +
	( 10'sd 311) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16502) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8272) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13162) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29583) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29396) * $signed(input_fmap_51[7:0]) +
	( 10'sd 342) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23686) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14993) * $signed(input_fmap_54[7:0]) +
	( 10'sd 295) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7965) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22528) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23149) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24351) * $signed(input_fmap_59[7:0]) +
	( 10'sd 448) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16000) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32740) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20425) * $signed(input_fmap_63[7:0]) +
	( 11'sd 943) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8894) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28337) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12504) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26292) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15432) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21672) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8654) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1907) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17226) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22609) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28538) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19080) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7060) * $signed(input_fmap_79[7:0]) +
	( 11'sd 587) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3576) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14820) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29579) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15678) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6195) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15425) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26622) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26538) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27535) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27565) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7031) * $signed(input_fmap_91[7:0]) +
	( 14'sd 8005) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1693) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4097) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10952) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25087) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18499) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9585) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31351) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10526) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28817) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10191) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17289) * $signed(input_fmap_105[7:0]) +
	( 11'sd 915) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17350) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28076) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20242) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30286) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29549) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28946) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17372) * $signed(input_fmap_113[7:0]) +
	( 11'sd 651) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29478) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13489) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12447) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24818) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10034) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2676) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27133) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1870) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11789) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31629) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32743) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3205) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15682) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 9'sd 203) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10659) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13019) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4496) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26888) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22045) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22819) * $signed(input_fmap_7[7:0]) +
	( 13'sd 4056) * $signed(input_fmap_8[7:0]) +
	( 9'sd 172) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10397) * $signed(input_fmap_10[7:0]) +
	( 15'sd 16304) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28706) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9486) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23301) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7997) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2578) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31408) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10924) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9951) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29984) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3320) * $signed(input_fmap_21[7:0]) +
	( 11'sd 659) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32328) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20932) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15422) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16500) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3525) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13037) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19439) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17884) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7463) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5884) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5714) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1768) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12531) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23405) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11082) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9594) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21947) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23526) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2769) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24457) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3006) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10835) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28831) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6527) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27568) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4634) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_50[7:0]) +
	( 11'sd 820) * $signed(input_fmap_51[7:0]) +
	( 11'sd 800) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4976) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7209) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27361) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17514) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6013) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30761) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23904) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17120) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14516) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13468) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12542) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17706) * $signed(input_fmap_66[7:0]) +
	( 14'sd 8099) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3881) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30729) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25639) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11516) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13145) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16845) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20821) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20453) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13642) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22986) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24475) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10019) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9576) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23046) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22756) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12811) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21319) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4713) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5652) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4922) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29769) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28549) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10061) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27230) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13654) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15920) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17089) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6554) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27487) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25512) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10142) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29256) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12836) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32034) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14134) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15983) * $signed(input_fmap_107[7:0]) +
	( 10'sd 362) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18130) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32371) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1076) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3212) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14653) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6160) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4672) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22103) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13394) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28656) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21081) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27296) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28564) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17726) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12915) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10832) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14417) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16337) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 15'sd 14124) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15102) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31018) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_5[7:0]) +
	( 9'sd 219) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26415) * $signed(input_fmap_8[7:0]) +
	( 8'sd 69) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21295) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12235) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15031) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22960) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10199) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11454) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6274) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28236) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24030) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24143) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12418) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2760) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6308) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6299) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22774) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17436) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26093) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4417) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27519) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21394) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18784) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24766) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11036) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25271) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28190) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19505) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30972) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18299) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24483) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22326) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8254) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22615) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26832) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15979) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18608) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11838) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24276) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14995) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14412) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6939) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11467) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22743) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10659) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24550) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28316) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25579) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8903) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28917) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15157) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23517) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15443) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25548) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27243) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5474) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11922) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15938) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24785) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31190) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19368) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12915) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22306) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17813) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15827) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16003) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31519) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27272) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3889) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18412) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3384) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30142) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4995) * $signed(input_fmap_95[7:0]) +
	( 10'sd 315) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22244) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26243) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21498) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29235) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2048) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15682) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5746) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31818) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22055) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30586) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10513) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31345) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28422) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3825) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24590) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17924) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24417) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14703) * $signed(input_fmap_117[7:0]) +
	( 11'sd 546) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2717) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2056) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6172) * $signed(input_fmap_122[7:0]) +
	( 10'sd 258) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14059) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17391) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21531) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 15'sd 10793) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26072) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26481) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25779) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8624) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10432) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11141) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10952) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24606) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19734) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9514) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6977) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12599) * $signed(input_fmap_16[7:0]) +
	( 11'sd 595) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5506) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11698) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15375) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11141) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12345) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31631) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13407) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11476) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30459) * $signed(input_fmap_29[7:0]) +
	( 10'sd 511) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27583) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10805) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13935) * $signed(input_fmap_33[7:0]) +
	( 9'sd 205) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8299) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14803) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22432) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13136) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9292) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14142) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30975) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7300) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12957) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17347) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24366) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31913) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21001) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1907) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22726) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1049) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18930) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27633) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30910) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31818) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1396) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11538) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22432) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9481) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27295) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26231) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31258) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10516) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25620) * $signed(input_fmap_68[7:0]) +
	( 11'sd 1004) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27093) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13156) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24983) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2382) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3180) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20555) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11314) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18034) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2723) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9398) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23512) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21256) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_85[7:0]) +
	( 5'sd 11) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11948) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25879) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8302) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_90[7:0]) +
	( 10'sd 494) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17471) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19281) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5722) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4756) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17904) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9227) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28923) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29149) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6680) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21230) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28859) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3043) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28040) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4231) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14556) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28812) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27180) * $signed(input_fmap_109[7:0]) +
	( 12'sd 2011) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8376) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13481) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21598) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12176) * $signed(input_fmap_114[7:0]) +
	( 11'sd 697) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10040) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30674) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14220) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13421) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8748) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28321) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24212) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29466) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19630) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16948) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 13'sd 3030) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17779) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14187) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1668) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13628) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1186) * $signed(input_fmap_6[7:0]) +
	( 11'sd 742) * $signed(input_fmap_7[7:0]) +
	( 10'sd 258) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14805) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15505) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25960) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25633) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15946) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11759) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13021) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14409) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5752) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15427) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19186) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21104) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19532) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28639) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26510) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8755) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2982) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4155) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15643) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8649) * $signed(input_fmap_31[7:0]) +
	( 11'sd 777) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1234) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4327) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15046) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6955) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19391) * $signed(input_fmap_39[7:0]) +
	( 11'sd 545) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28604) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18478) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13110) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21214) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17561) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12031) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23255) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32568) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30178) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11876) * $signed(input_fmap_51[7:0]) +
	( 11'sd 533) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21659) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16398) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26897) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28544) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15694) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12700) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12574) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18625) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14791) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21298) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6763) * $signed(input_fmap_63[7:0]) +
	( 9'sd 158) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29266) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9067) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27847) * $signed(input_fmap_68[7:0]) +
	( 14'sd 8143) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12449) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14635) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1113) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8821) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6526) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26654) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10139) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30174) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1599) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16329) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23913) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29802) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24437) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27418) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30107) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26439) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16125) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23133) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9345) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32184) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24964) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18039) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5707) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29448) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3790) * $signed(input_fmap_97[7:0]) +
	( 14'sd 8150) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18842) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17074) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31021) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21473) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27095) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13154) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24726) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10815) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14039) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28555) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23743) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6230) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15968) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1485) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9255) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9253) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11900) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3459) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28510) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22215) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12197) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17088) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_122[7:0]) +
	( 11'sd 641) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24261) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2514) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17118) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 16'sd 19079) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22194) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19293) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29556) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24651) * $signed(input_fmap_4[7:0]) +
	( 8'sd 75) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9354) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24623) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31547) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1967) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2264) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24120) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10541) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14203) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17680) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15922) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31112) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20740) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12603) * $signed(input_fmap_18[7:0]) +
	( 12'sd 2010) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11285) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19899) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12385) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29738) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14758) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5227) * $signed(input_fmap_26[7:0]) +
	( 15'sd 16333) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26627) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3832) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14012) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14000) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30515) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1274) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10003) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1157) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27602) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19966) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32534) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14503) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13469) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32282) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23204) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19158) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1027) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1763) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6947) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12886) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29181) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24641) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8547) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6227) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18126) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21746) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21908) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27104) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26283) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21822) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12896) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14600) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5174) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3285) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8718) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24155) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15284) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17033) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14736) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11467) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22725) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28327) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13143) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14780) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26940) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18203) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16621) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24775) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14647) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4890) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31939) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26251) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19630) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17363) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15209) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9268) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21119) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30228) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31689) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23308) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10923) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13525) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16780) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16383) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1460) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32366) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14009) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18152) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27376) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8869) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14997) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22261) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30821) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32339) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25809) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2505) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22029) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24068) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12184) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10798) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9156) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17819) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4897) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19835) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5601) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26080) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27915) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26370) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4764) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12699) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_126[7:0]) +
	( 11'sd 667) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 16'sd 26439) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24503) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24086) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13650) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15689) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22944) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32208) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24647) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30344) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23879) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2294) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19463) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32480) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32223) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9598) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7543) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20967) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14646) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25439) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24222) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5861) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3491) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26239) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15313) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31612) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29740) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16254) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20645) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26910) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12323) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18787) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32115) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14549) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29068) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11647) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20181) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20731) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19478) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10856) * $signed(input_fmap_46[7:0]) +
	( 8'sd 125) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5462) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4551) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11254) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24238) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2111) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27564) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22418) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8273) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29519) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32757) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20216) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26462) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13540) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4843) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11509) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9801) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2614) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16926) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21447) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7625) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28598) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1954) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25924) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31755) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16108) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17749) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27966) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22137) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19211) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13627) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12996) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10022) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32252) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15323) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28511) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9205) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15028) * $signed(input_fmap_93[7:0]) +
	( 9'sd 218) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16851) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27076) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28693) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32193) * $signed(input_fmap_99[7:0]) +
	( 11'sd 867) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26038) * $signed(input_fmap_101[7:0]) +
	( 11'sd 582) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1314) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32211) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30573) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4814) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25790) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4974) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17682) * $signed(input_fmap_111[7:0]) +
	( 12'sd 2004) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22410) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17906) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19480) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12985) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21940) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3171) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1108) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25401) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22281) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6094) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19325) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1340) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 15'sd 10681) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8429) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30499) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19405) * $signed(input_fmap_4[7:0]) +
	( 7'sd 51) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15012) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14332) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12038) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17738) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31515) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20905) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10708) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10973) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26918) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22740) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4953) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16674) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11217) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15512) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11485) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13198) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6456) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25716) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21392) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17103) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26275) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14604) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21985) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26279) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11187) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29975) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8737) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9604) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31257) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12962) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15837) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2780) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17322) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19462) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9422) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13064) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13814) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23472) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28762) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2792) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14211) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28889) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27106) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30430) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10429) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14466) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32042) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11650) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17293) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11295) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13123) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10895) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23408) * $signed(input_fmap_62[7:0]) +
	( 10'sd 297) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14408) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3423) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14103) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18184) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8426) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16393) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30087) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1640) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6307) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28117) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32368) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1834) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13851) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4520) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3274) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1567) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29956) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8258) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14310) * $signed(input_fmap_83[7:0]) +
	( 14'sd 8176) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2165) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5836) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25036) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18086) * $signed(input_fmap_88[7:0]) +
	( 6'sd 27) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17403) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21075) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14046) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27155) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4772) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16821) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6928) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1610) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6849) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14662) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21314) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16643) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4204) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13176) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8492) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21693) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18922) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19447) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19729) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14690) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26373) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16870) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3449) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9484) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27528) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10690) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8737) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7044) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23456) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19574) * $signed(input_fmap_126[7:0]) +
	( 10'sd 305) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 16'sd 19201) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29918) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19217) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20747) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12663) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8716) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19491) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_7[7:0]) +
	( 11'sd 669) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29406) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4188) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6500) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13470) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10601) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26301) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32149) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17405) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23409) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24450) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28013) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14200) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11244) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31596) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6294) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28180) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8418) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23747) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26905) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27856) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22145) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13444) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29645) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23355) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12618) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26534) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4422) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14243) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15597) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8761) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16132) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27486) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23963) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13553) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28085) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28238) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24865) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2069) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19274) * $signed(input_fmap_52[7:0]) +
	( 11'sd 707) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3879) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23222) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13983) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26300) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8391) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32583) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3441) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13441) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20546) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17889) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6741) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3400) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21588) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27803) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21935) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10622) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17355) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7808) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5686) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26269) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18437) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7741) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31440) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17286) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24352) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23253) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8725) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1047) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9966) * $signed(input_fmap_87[7:0]) +
	( 10'sd 381) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13702) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26858) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12145) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3890) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16099) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2194) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28545) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23785) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6022) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32699) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9480) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7970) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32591) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11795) * $signed(input_fmap_103[7:0]) +
	( 10'sd 435) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32171) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27538) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20199) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12921) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3649) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32616) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2730) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11881) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25897) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23555) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18025) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32634) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2130) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_120[7:0]) +
	( 10'sd 476) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19857) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7213) * $signed(input_fmap_123[7:0]) +
	( 9'sd 198) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9558) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32636) * $signed(input_fmap_126[7:0]) +
	( 8'sd 76) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 16'sd 20299) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31039) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25480) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31217) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15147) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31006) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23962) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24195) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22630) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3962) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23773) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4539) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2874) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3509) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14911) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6385) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29347) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13755) * $signed(input_fmap_20[7:0]) +
	( 10'sd 419) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31422) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5385) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19405) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18744) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13751) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32640) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25179) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21288) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17131) * $signed(input_fmap_31[7:0]) +
	( 10'sd 386) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14205) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4148) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7969) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8443) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15242) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1531) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11332) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10192) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4313) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29927) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3714) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9717) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31213) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11828) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25173) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32475) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26860) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17420) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14421) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31966) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20525) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26499) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21719) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15749) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20088) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6571) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11409) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4696) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13051) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9732) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19145) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21193) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4283) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26032) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9307) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31437) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28779) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3153) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22630) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16269) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17383) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3365) * $signed(input_fmap_80[7:0]) +
	( 10'sd 479) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12445) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16967) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26512) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2890) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1502) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23625) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1782) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12583) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7428) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14724) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1599) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26757) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23375) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1250) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15073) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8832) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15690) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28186) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1813) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17549) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14216) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22807) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10062) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28151) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19970) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5074) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20166) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16719) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12838) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28350) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4136) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7294) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18852) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16692) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20771) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24227) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21690) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26394) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2583) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12466) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 12'sd 1891) * $signed(input_fmap_0[7:0]) +
	( 7'sd 57) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28891) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8917) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5065) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13028) * $signed(input_fmap_6[7:0]) +
	( 14'sd 8033) * $signed(input_fmap_7[7:0]) +
	( 11'sd 849) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27713) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11807) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9815) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29120) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3596) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23822) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23366) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30297) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12965) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1148) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2372) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9669) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24898) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24563) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22098) * $signed(input_fmap_25[7:0]) +
	( 10'sd 369) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23801) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3090) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21981) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31239) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20164) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29819) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24836) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23482) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26646) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27305) * $signed(input_fmap_36[7:0]) +
	( 10'sd 478) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2518) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29686) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11025) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1757) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20219) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4680) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25543) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14873) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2690) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15213) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9395) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24825) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2461) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3112) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21008) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19934) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24284) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8462) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12998) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10475) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4677) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17138) * $signed(input_fmap_60[7:0]) +
	( 13'sd 4055) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26036) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7579) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6986) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21620) * $signed(input_fmap_66[7:0]) +
	( 11'sd 589) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18201) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32364) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6635) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5938) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20341) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24945) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10315) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20858) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29620) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26633) * $signed(input_fmap_80[7:0]) +
	( 11'sd 1008) * $signed(input_fmap_81[7:0]) +
	( 13'sd 4012) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27554) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23128) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5945) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5629) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11925) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32452) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21461) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17018) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31630) * $signed(input_fmap_92[7:0]) +
	( 11'sd 691) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9979) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12541) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11045) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15632) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16383) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32166) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10677) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13494) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6968) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10966) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5642) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13056) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32180) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14076) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27841) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22233) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17099) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2048) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16747) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22099) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8216) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17799) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13927) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24042) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23333) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30082) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21174) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4990) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13175) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2783) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5941) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 15'sd 9521) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27559) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9183) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14364) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21519) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24181) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29450) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2274) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15527) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9996) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16508) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20370) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10214) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17909) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13583) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20789) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1060) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14059) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3753) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10458) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5322) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11253) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1945) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2812) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12519) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10944) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5717) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19078) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20149) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15461) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26011) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16493) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22900) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22664) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7724) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22350) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3401) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15564) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14512) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_42[7:0]) +
	( 11'sd 635) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7234) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2873) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1557) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11502) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9687) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8896) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28225) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23109) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19954) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25898) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_56[7:0]) +
	( 11'sd 658) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6891) * $signed(input_fmap_58[7:0]) +
	( 11'sd 595) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3938) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10399) * $signed(input_fmap_61[7:0]) +
	( 11'sd 609) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15141) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14344) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1930) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17749) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13486) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3272) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5479) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7769) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7251) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15476) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26603) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17132) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10597) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21351) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14337) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11416) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25221) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24481) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17124) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28008) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30991) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22227) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17042) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26889) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14330) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12724) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11540) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15882) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2622) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31483) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30939) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13166) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18098) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9615) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3193) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9935) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26488) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6031) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26281) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10730) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1962) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32389) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22658) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11602) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18019) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32711) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17074) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11006) * $signed(input_fmap_115[7:0]) +
	( 9'sd 169) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11446) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27434) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28402) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28688) * $signed(input_fmap_121[7:0]) +
	( 12'sd 2003) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1768) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32642) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10343) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27713) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22482) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 16'sd 30266) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13947) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5882) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11145) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6732) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21071) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10257) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19732) * $signed(input_fmap_7[7:0]) +
	( 11'sd 710) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20350) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12122) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23511) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29994) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4307) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11561) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7379) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9420) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9460) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9645) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3368) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_20[7:0]) +
	( 11'sd 720) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3119) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16937) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1162) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14570) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30806) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23104) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13487) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18778) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8307) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3387) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9008) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20824) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6637) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16884) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4819) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18352) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13655) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7810) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15001) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12276) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28978) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20061) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18080) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10890) * $signed(input_fmap_50[7:0]) +
	( 11'sd 621) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3249) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11378) * $signed(input_fmap_53[7:0]) +
	( 14'sd 8118) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4230) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3460) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30917) * $signed(input_fmap_58[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14299) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9283) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28142) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16845) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11402) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26856) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9606) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12409) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19184) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15471) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14186) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6584) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1550) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29978) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30311) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17397) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16907) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17188) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15995) * $signed(input_fmap_81[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6609) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25464) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32298) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19567) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3953) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6822) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1822) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27037) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9536) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27670) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1341) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10998) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31715) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16315) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15026) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28490) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32571) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2151) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11770) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27892) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4508) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12139) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23121) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8758) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8273) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14210) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24153) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17544) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1071) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18675) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14721) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6702) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1492) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14413) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9388) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11787) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6119) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27256) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3084) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 14'sd 6618) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5805) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29806) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19089) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3198) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15371) * $signed(input_fmap_7[7:0]) +
	( 11'sd 808) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14590) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17806) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24381) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12976) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26216) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32177) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28995) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23229) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14925) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17958) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1242) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20663) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11866) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28427) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3830) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17393) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30515) * $signed(input_fmap_27[7:0]) +
	( 12'sd 2021) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1090) * $signed(input_fmap_29[7:0]) +
	( 10'sd 393) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10778) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24543) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30286) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14597) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16486) * $signed(input_fmap_35[7:0]) +
	( 4'sd 7) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12186) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15390) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4546) * $signed(input_fmap_39[7:0]) +
	( 10'sd 442) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15771) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19823) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13879) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8935) * $signed(input_fmap_45[7:0]) +
	( 11'sd 958) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21625) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1754) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1380) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12816) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29967) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6656) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23660) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3854) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26739) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22049) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21545) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31768) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17557) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29529) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24865) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16859) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7683) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1051) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30557) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13376) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7413) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15525) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16408) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12556) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23175) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21469) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27907) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9325) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14210) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3609) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2648) * $signed(input_fmap_82[7:0]) +
	( 11'sd 794) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13377) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9356) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10469) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23827) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7038) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28536) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4816) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29389) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18223) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21288) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26399) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27980) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6332) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12874) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32614) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20783) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20842) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7378) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9972) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12859) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25282) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3456) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9134) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29687) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16645) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21571) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1500) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31265) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5056) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7304) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29668) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32417) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11393) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22191) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1704) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8075) * $signed(input_fmap_122[7:0]) +
	( 10'sd 256) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4947) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27939) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 15'sd 15410) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_1[7:0]) +
	( 14'sd 8168) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20991) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13253) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25186) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23543) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18650) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9763) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1904) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1462) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7030) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22756) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3777) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2929) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13185) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8311) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1456) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20527) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25928) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27168) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6326) * $signed(input_fmap_24[7:0]) +
	( 11'sd 862) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30970) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28397) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9611) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16519) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5919) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9807) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32602) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11708) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18624) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3099) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10824) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4907) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10299) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14482) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23392) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2228) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16065) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9538) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26132) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13053) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15302) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6464) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10897) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9597) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23388) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22439) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16897) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8250) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30224) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31155) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11679) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16687) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11394) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25444) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31236) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9185) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26002) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28234) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_69[7:0]) +
	( 9'sd 255) * $signed(input_fmap_70[7:0]) +
	( 14'sd 8051) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22720) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11229) * $signed(input_fmap_74[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31128) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29741) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1474) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17054) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6065) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16265) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18508) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32367) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11621) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30694) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20272) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29036) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15509) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21067) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12700) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9772) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2506) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12944) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11687) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8254) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17842) * $signed(input_fmap_100[7:0]) +
	( 11'sd 754) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8726) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14520) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29692) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5214) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3578) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24262) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13576) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23732) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32589) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6442) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8767) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3484) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31652) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2895) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29722) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32191) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31104) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6557) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24136) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11675) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6103) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6614) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 15'sd 8408) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26555) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17613) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15869) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22925) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18317) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13774) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15179) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16742) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4133) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5168) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19909) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_13[7:0]) +
	( 11'sd 904) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31613) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1779) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16714) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29695) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11318) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29981) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9102) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21760) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6933) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29932) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14857) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4652) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2994) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31603) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13960) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23615) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13002) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31241) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5499) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7365) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25915) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2849) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31219) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17195) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29015) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24588) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21593) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26925) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3883) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9360) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7196) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27439) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32103) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13747) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18199) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4680) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12712) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27819) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24595) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19661) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18161) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9065) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3452) * $signed(input_fmap_63[7:0]) +
	( 11'sd 617) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12785) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22430) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22092) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32638) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31853) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3364) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21907) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2254) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1588) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11588) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8245) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32351) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27560) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19206) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22855) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23508) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22131) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1385) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13547) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31401) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26001) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31001) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2911) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27152) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28616) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21404) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25838) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23249) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20225) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1743) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27995) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20316) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20874) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19568) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7607) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8949) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3485) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27915) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28872) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30046) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15789) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6501) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7182) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5898) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6545) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27139) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5533) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12211) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7431) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31558) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6168) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31087) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10502) * $signed(input_fmap_124[7:0]) +
	( 11'sd 829) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7875) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32501) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 16'sd 29768) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6111) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21903) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21824) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20402) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24022) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23284) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11819) * $signed(input_fmap_9[7:0]) +
	( 11'sd 890) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7172) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14691) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32465) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11079) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1251) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32110) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_17[7:0]) +
	( 9'sd 208) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20841) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15411) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4639) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30566) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25945) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12968) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10257) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23296) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14607) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30571) * $signed(input_fmap_28[7:0]) +
	( 12'sd 2032) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14277) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26317) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1754) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15304) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5671) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15282) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7318) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31594) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24917) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14483) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21405) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25379) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15349) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12917) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27358) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11425) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31236) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27247) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3287) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17870) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30933) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26015) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18932) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15614) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29568) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14384) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_65[7:0]) +
	( 8'sd 99) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6324) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23174) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25674) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6911) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7171) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8988) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15183) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25872) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1103) * $signed(input_fmap_76[7:0]) +
	( 11'sd 576) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29766) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26004) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28581) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2821) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20011) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21455) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7575) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9741) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15145) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23584) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1111) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11939) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30209) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6047) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25766) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9292) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32016) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28029) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7191) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21139) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1202) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12653) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25929) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7590) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27193) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19765) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15816) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18771) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17943) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25054) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12512) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23044) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10146) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5458) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13867) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24317) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27069) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21116) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3284) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21083) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23483) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31554) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9127) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 16'sd 19627) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23888) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28445) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19233) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_5[7:0]) +
	( 11'sd 543) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19402) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10245) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26275) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20360) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15459) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12376) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27433) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9503) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22003) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26443) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19666) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11494) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12198) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32164) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31760) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13941) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23357) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7640) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30530) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14051) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7145) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12983) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6621) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19112) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11692) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2493) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9540) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2747) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5571) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24694) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22716) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21671) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14799) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12136) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3368) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31484) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27006) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5063) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3773) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17578) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25585) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16836) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14111) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3675) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16204) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31396) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14469) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12645) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31355) * $signed(input_fmap_62[7:0]) +
	( 11'sd 854) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15043) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29030) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16846) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29358) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5886) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11850) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18777) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10801) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19290) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11891) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20064) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25881) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28867) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11788) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2116) * $signed(input_fmap_81[7:0]) +
	( 14'sd 8156) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6604) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1312) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18838) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27287) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22151) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14669) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31162) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9126) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10401) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8641) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8955) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11045) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29904) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29384) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27795) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10634) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27829) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11790) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21446) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15266) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24750) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27258) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7497) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31293) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11004) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30945) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3669) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26233) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31297) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29042) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13621) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17823) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8697) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8002) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17104) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11803) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1935) * $signed(input_fmap_125[7:0]) +
	( 12'sd 2025) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23687) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 15'sd 12133) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30644) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24219) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21019) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25261) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6769) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2889) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10430) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24020) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31243) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18814) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25162) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17149) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10917) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4124) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29977) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24256) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27318) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4117) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3158) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30160) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11838) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31180) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10929) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21053) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16382) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11218) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27209) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11032) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21431) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2201) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16477) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16963) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17450) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23365) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6716) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15734) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13766) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20199) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11097) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29331) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23767) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21531) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15368) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16478) * $signed(input_fmap_51[7:0]) +
	( 11'sd 961) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13956) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10459) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11381) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16529) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5644) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16032) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11474) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14243) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22625) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5121) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27175) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30005) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16480) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20400) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13103) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29723) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29232) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14619) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22197) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10224) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20778) * $signed(input_fmap_79[7:0]) +
	( 8'sd 94) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29535) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23780) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29784) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16066) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23964) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12811) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7449) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17284) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17573) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15968) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8413) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12155) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4275) * $signed(input_fmap_93[7:0]) +
	( 8'sd 83) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32301) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13749) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1989) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15680) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5460) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15617) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3291) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3364) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31429) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3301) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26329) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25994) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25457) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2844) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14744) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21984) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20220) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3234) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29152) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9116) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20826) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28395) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28976) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13332) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5270) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31111) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1432) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1592) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 15'sd 13197) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7324) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12570) * $signed(input_fmap_2[7:0]) +
	( 10'sd 391) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19464) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19893) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6126) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23001) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30121) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29792) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28877) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14494) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26158) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4497) * $signed(input_fmap_14[7:0]) +
	( 11'sd 998) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7823) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15854) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25153) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22163) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6975) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24946) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28758) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7122) * $signed(input_fmap_24[7:0]) +
	( 12'sd 2007) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29353) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23349) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24328) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14021) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8726) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16690) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7493) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32500) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20999) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28890) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3847) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4330) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30802) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10472) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13523) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22555) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6192) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8543) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9897) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6848) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6042) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14046) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24120) * $signed(input_fmap_53[7:0]) +
	( 11'sd 694) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15848) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8985) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1111) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31118) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29274) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25155) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20181) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13336) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17154) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10376) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26528) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10314) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8544) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26897) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30378) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2828) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17251) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16770) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29256) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24154) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16690) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11564) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29709) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24375) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26778) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18019) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14954) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17983) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2414) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24316) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32343) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3862) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15080) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32616) * $signed(input_fmap_93[7:0]) +
	( 11'sd 716) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20086) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28267) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26698) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24866) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22673) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23731) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5824) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12768) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23477) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23631) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26865) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23160) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31008) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10621) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21067) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16715) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17331) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8978) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8675) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22886) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11798) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28318) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28648) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23618) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25398) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9539) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3961) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23518) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23667) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24364) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 13'sd 3116) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13618) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14209) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15686) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11589) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26860) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18588) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24791) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29555) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17466) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8948) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28045) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27245) * $signed(input_fmap_14[7:0]) +
	( 14'sd 8074) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25397) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7338) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6355) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22615) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28944) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28594) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6469) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_26[7:0]) +
	( 11'sd 978) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11926) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5015) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18423) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26498) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24119) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17045) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25839) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5407) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1749) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1500) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19233) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10784) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13831) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16558) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23254) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8872) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19564) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26128) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32146) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13581) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5481) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1962) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4751) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19179) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29158) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25767) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16798) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27777) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24434) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12807) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5867) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5180) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20669) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17527) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11282) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17080) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30776) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27301) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7145) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1393) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13587) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18621) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28754) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12132) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18217) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6912) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1230) * $signed(input_fmap_83[7:0]) +
	( 11'sd 592) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30763) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19533) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32303) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3809) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16248) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26366) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9600) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2164) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19338) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14138) * $signed(input_fmap_95[7:0]) +
	( 10'sd 399) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25872) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4395) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_99[7:0]) +
	( 10'sd 368) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27473) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30192) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13637) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4828) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4600) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13118) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20189) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28477) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28068) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26221) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21833) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14451) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7591) * $signed(input_fmap_116[7:0]) +
	( 11'sd 844) * $signed(input_fmap_117[7:0]) +
	( 11'sd 849) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9113) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14899) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2459) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8092) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19985) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22410) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11952) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10696) * $signed(input_fmap_126[7:0]) +
	( 7'sd 55) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 16'sd 27160) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27810) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11132) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30083) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12270) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13978) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6332) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5817) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18947) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12217) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14142) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23117) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3770) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12195) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3889) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10120) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10026) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15321) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11173) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3574) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2424) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30451) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17179) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27312) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6017) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13303) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31033) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11341) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21287) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25307) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9207) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16373) * $signed(input_fmap_34[7:0]) +
	( 11'sd 696) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2059) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6376) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18934) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22388) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16924) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27148) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27033) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24185) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14039) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4642) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2937) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29473) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21955) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7342) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2155) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13675) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30532) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28021) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26942) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4349) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8999) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21835) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19354) * $signed(input_fmap_63[7:0]) +
	( 11'sd 709) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27386) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8883) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8283) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13652) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24777) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32266) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16195) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8034) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1728) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15370) * $signed(input_fmap_75[7:0]) +
	( 11'sd 981) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1290) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8834) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29247) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10994) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20254) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26017) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19562) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3837) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11761) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25411) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17824) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18568) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23048) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19297) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9077) * $signed(input_fmap_91[7:0]) +
	( 9'sd 178) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32681) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7851) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11818) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11524) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11814) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20413) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4558) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3018) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28659) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22638) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31857) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12749) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6840) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15695) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29402) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3951) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14364) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30690) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7017) * $signed(input_fmap_112[7:0]) +
	( 11'sd 917) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8872) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5021) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30739) * $signed(input_fmap_118[7:0]) +
	( 13'sd 4068) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18810) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3991) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32183) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10458) * $signed(input_fmap_124[7:0]) +
	( 15'sd 16293) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23561) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20293) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 16'sd 19283) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22515) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28320) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30545) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7566) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26199) * $signed(input_fmap_5[7:0]) +
	( 10'sd 424) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15539) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24074) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11361) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22437) * $signed(input_fmap_10[7:0]) +
	( 11'sd 827) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21819) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22022) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17505) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24965) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29320) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2867) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31543) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24248) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17709) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17750) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10130) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17424) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8189) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27173) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14439) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5378) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15237) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21765) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4229) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22622) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23828) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10276) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16980) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24810) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3780) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31794) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3556) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7682) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6861) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1261) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19698) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23837) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26153) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20451) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6357) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31312) * $signed(input_fmap_49[7:0]) +
	( 14'sd 8179) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1213) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22060) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15231) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12699) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30365) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25967) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2963) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12217) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1475) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26148) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11260) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12166) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14238) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28528) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14641) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3179) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6190) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10566) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32359) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24021) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14254) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26648) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24804) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_78[7:0]) +
	( 10'sd 420) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7007) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18514) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32456) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12895) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28733) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9406) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5097) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24049) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30069) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13491) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26543) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12914) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23839) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25199) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21019) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9699) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5397) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18254) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29201) * $signed(input_fmap_100[7:0]) +
	( 11'sd 660) * $signed(input_fmap_101[7:0]) +
	( 11'sd 824) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24499) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20824) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30069) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15584) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22860) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15178) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7022) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1743) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2346) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28734) * $signed(input_fmap_112[7:0]) +
	( 14'sd 8119) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11423) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3029) * $signed(input_fmap_115[7:0]) +
	( 9'sd 208) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5070) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31994) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14951) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29173) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18474) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17782) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3096) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1831) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18654) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28232) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 14'sd 7223) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5303) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22339) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28281) * $signed(input_fmap_3[7:0]) +
	( 13'sd 4064) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10686) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9123) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14449) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22483) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11182) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5749) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9627) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24333) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25317) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20030) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11563) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32762) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29781) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12869) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20991) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18852) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17377) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30234) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30132) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15791) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27554) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28752) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26027) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7244) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24889) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19167) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10518) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21524) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29823) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29509) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15944) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23330) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7493) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26511) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4659) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17546) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7539) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1403) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27969) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26503) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24410) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31685) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6233) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9722) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9545) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2552) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13965) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5700) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25192) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12693) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16477) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31410) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31932) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26099) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6842) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4746) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30825) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11039) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29866) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11162) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5666) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19762) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17761) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10208) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2465) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5935) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31051) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27331) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27019) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17258) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28508) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25625) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14693) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7367) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19335) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11065) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20654) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22207) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28654) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28363) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13747) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17008) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3804) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8906) * $signed(input_fmap_98[7:0]) +
	( 13'sd 4084) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4280) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19321) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2309) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18807) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14990) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1227) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14540) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12786) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15172) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21288) * $signed(input_fmap_109[7:0]) +
	( 8'sd 99) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21614) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18415) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23982) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16323) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21030) * $signed(input_fmap_120[7:0]) +
	( 10'sd 404) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23471) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10845) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6196) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 11'sd 600) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27287) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11487) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28407) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25849) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30243) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6442) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27085) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20526) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28520) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8437) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4967) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6748) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2434) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23827) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25592) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28050) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30420) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30200) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23321) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12507) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32151) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25480) * $signed(input_fmap_23[7:0]) +
	( 10'sd 380) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8148) * $signed(input_fmap_25[7:0]) +
	( 11'sd 738) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31377) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16076) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24712) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19978) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23135) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30067) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30378) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13805) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27362) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1880) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26853) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13052) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3865) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15314) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2441) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3406) * $signed(input_fmap_44[7:0]) +
	( 10'sd 371) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28532) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30101) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4659) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10963) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8430) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21575) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3517) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11210) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19946) * $signed(input_fmap_54[7:0]) +
	( 10'sd 258) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19273) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1546) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23714) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6929) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21691) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28545) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9864) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28896) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25681) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22592) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17442) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1216) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21401) * $signed(input_fmap_68[7:0]) +
	( 10'sd 476) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32330) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9503) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3048) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29744) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1459) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10310) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26860) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28638) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13945) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15398) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3314) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15853) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15019) * $signed(input_fmap_85[7:0]) +
	( 11'sd 811) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19432) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19778) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28958) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13565) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17770) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7467) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10908) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29249) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20908) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32712) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13511) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4702) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26522) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19453) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6740) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7751) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22963) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24129) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2244) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18247) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9269) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7707) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12332) * $signed(input_fmap_113[7:0]) +
	( 11'sd 973) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8309) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19072) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16605) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10838) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12633) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17988) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9876) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32582) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30490) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2461) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7273) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 16'sd 20745) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19074) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9136) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13194) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7170) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19420) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19116) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23677) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23806) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4268) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5629) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22580) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32508) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15368) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30840) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31946) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22410) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14387) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18993) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25560) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17723) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6947) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10349) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19301) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24720) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6553) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21229) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10820) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8453) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25874) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12555) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10040) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26749) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7013) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27492) * $signed(input_fmap_37[7:0]) +
	( 13'sd 4006) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4190) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27453) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17622) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5693) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23914) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17773) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27755) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7888) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17924) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13013) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8990) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23229) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1896) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13172) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24805) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23638) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19489) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5588) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26553) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19442) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19156) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23756) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3046) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19902) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26251) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13722) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19174) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9325) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25042) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29336) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30041) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15729) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19977) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5618) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23474) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16058) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30986) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32268) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20917) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9571) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8138) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19138) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32037) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10714) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13290) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12791) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26975) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30865) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20448) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27375) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14288) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12940) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1307) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7722) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3618) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6945) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20758) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31499) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19163) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3769) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1339) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19409) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32745) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10221) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11056) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9571) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12098) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5722) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8932) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12419) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32033) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15164) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2902) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30912) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 16'sd 16428) * $signed(input_fmap_0[7:0]) +
	( 11'sd 1008) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13801) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6726) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6273) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3316) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28762) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7263) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30828) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14274) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3608) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30962) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7514) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14671) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1487) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26625) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25650) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23864) * $signed(input_fmap_17[7:0]) +
	( 11'sd 668) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12663) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16671) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8738) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24640) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20972) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25418) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15183) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27070) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27200) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30872) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11338) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22016) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5415) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11192) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4930) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1918) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6267) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18710) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27780) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26955) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20213) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12112) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15489) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10856) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16859) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12902) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6293) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12102) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13516) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24247) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16468) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11712) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25476) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13375) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21769) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10936) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2482) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15969) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26865) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11474) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1529) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28607) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5732) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8595) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30891) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18472) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11497) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14792) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22704) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3793) * $signed(input_fmap_76[7:0]) +
	( 11'sd 910) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4761) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32465) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25700) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9884) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27021) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17103) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18557) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3887) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6189) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26861) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12658) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13456) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7033) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20403) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2481) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23834) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17238) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29611) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21450) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2830) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4705) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11592) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6645) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30236) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24343) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31945) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25518) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26391) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29311) * $signed(input_fmap_111[7:0]) +
	( 10'sd 468) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9346) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13148) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31157) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15108) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26573) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9632) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18554) * $signed(input_fmap_119[7:0]) +
	( 8'sd 122) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21796) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9360) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12981) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16620) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26047) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7094) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32155) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 16'sd 30443) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5761) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30536) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19437) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29179) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4482) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5626) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25869) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30586) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13397) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10490) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2370) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12839) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29444) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19340) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9717) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22898) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22666) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10954) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17526) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16814) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2254) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18339) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13407) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27249) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10260) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6708) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31977) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25274) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19147) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18027) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16173) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21989) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29352) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27566) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2154) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15894) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32657) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9403) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13717) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6836) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2995) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17615) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26698) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31980) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9107) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10851) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29692) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14543) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15246) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21598) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23305) * $signed(input_fmap_55[7:0]) +
	( 11'sd 942) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8371) * $signed(input_fmap_57[7:0]) +
	( 13'sd 4066) * $signed(input_fmap_58[7:0]) +
	( 14'sd 8151) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32503) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9044) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8503) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30662) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12164) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31046) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30391) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11735) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8642) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14962) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18445) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28557) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21399) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2924) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26597) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_76[7:0]) +
	( 14'sd 8125) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15089) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12510) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25434) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25964) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2706) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32026) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14622) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11952) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2257) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9036) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14964) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8674) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24798) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30179) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17555) * $signed(input_fmap_94[7:0]) +
	( 10'sd 346) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19941) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10400) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23978) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12554) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27804) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31937) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3930) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12712) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31809) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27756) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30172) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9518) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12517) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1539) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26995) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15681) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6290) * $signed(input_fmap_119[7:0]) +
	( 15'sd 16368) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17960) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21722) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4393) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4562) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27893) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 15'sd 12250) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16589) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22647) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23260) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2709) * $signed(input_fmap_4[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8933) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22748) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16121) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22920) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17063) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3606) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24831) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8235) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21564) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24603) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_17[7:0]) +
	( 11'sd 961) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9617) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30263) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12551) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18957) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1185) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29918) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14993) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29041) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20663) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23446) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2551) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10151) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30100) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29957) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16593) * $signed(input_fmap_34[7:0]) +
	( 5'sd 11) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10693) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27623) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29101) * $signed(input_fmap_38[7:0]) +
	( 10'sd 265) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15849) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13408) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14835) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8942) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30042) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6616) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24336) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18719) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14486) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22235) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11001) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18662) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2690) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16516) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12919) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18426) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5432) * $signed(input_fmap_58[7:0]) +
	( 12'sd 2002) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12797) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8485) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31601) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13277) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26121) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16898) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16854) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22999) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21837) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6103) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17364) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15326) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3416) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20864) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10582) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12423) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8905) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28481) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2480) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9187) * $signed(input_fmap_85[7:0]) +
	( 12'sd 2004) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3284) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18760) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19199) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13624) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29006) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12488) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8248) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10730) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31955) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22203) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24989) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28702) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13712) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1696) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10555) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19064) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23927) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11507) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24994) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11049) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2608) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3387) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28797) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31301) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10186) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24069) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5271) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7693) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21198) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19983) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14739) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28524) * $signed(input_fmap_123[7:0]) +
	( 14'sd 8012) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22615) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3030) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17594) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 16'sd 19859) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24342) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4689) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20452) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12083) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29233) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30223) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4140) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10158) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23105) * $signed(input_fmap_11[7:0]) +
	( 11'sd 647) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10438) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26829) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32268) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30073) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5013) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16658) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25964) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28748) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31773) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24109) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32585) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28793) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8842) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32089) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19680) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14499) * $signed(input_fmap_30[7:0]) +
	( 11'sd 528) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13896) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25395) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4789) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27791) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8480) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29157) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22155) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10478) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18058) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3077) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22421) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28687) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24713) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18666) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8845) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6253) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15105) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9245) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18187) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30204) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19238) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15910) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5105) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25259) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12854) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19484) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28460) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29601) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31607) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26936) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23753) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30550) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3902) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21860) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20610) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10233) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27212) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6189) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15092) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18916) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28465) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15276) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10142) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19462) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31053) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7025) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28564) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29201) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8781) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29057) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11939) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3817) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6249) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27060) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17134) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3963) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27009) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31723) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13650) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23164) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25975) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4968) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21042) * $signed(input_fmap_105[7:0]) +
	( 11'sd 592) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1364) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10285) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3275) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10495) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12760) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29875) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30365) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5667) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10250) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24241) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11816) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13786) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1410) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4805) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26386) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27082) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28864) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22862) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13908) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 16'sd 26933) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2844) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29016) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25220) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7825) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12987) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9155) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3094) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5985) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11885) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28940) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21441) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26530) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18762) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10541) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21935) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16699) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12873) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30420) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28787) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20719) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21449) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18248) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31882) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1896) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13802) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14624) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16586) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9762) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3143) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30940) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12184) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30522) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25583) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26168) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4327) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26771) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2101) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3323) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8331) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11518) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13527) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25852) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16898) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2640) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31751) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3063) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29961) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19166) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23955) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29854) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12299) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20722) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12076) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4296) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5186) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28553) * $signed(input_fmap_65[7:0]) +
	( 11'sd 600) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7728) * $signed(input_fmap_67[7:0]) +
	( 10'sd 473) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4235) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27363) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12532) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31301) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29764) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22390) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4975) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16637) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3561) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5519) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1350) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32361) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30141) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4539) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6831) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10471) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1772) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6202) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12100) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17587) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14834) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19169) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2410) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28350) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16332) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29195) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23389) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30201) * $signed(input_fmap_101[7:0]) +
	( 12'sd 2022) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17144) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32330) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26081) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30701) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7902) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25226) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26207) * $signed(input_fmap_111[7:0]) +
	( 9'sd 146) * $signed(input_fmap_112[7:0]) +
	( 11'sd 648) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20553) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13450) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13379) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31286) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25347) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18975) * $signed(input_fmap_120[7:0]) +
	( 10'sd 462) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27202) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2480) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17564) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12925) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24970) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 14'sd 5542) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11239) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28911) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2796) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23852) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18598) * $signed(input_fmap_7[7:0]) +
	( 14'sd 8100) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23405) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1366) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31673) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6197) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17019) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26245) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20157) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31845) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28667) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23849) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17427) * $signed(input_fmap_20[7:0]) +
	( 9'sd 200) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15682) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1154) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29791) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24660) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21832) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13178) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18948) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23287) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21170) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6000) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24585) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20761) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13335) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20951) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12662) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31760) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31647) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13339) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7715) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29438) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11914) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1359) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10870) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28697) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2423) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32030) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13291) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14695) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29528) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1465) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18166) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5784) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3148) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14044) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7553) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15136) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30638) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22270) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29569) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16104) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7206) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20075) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5704) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28686) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12179) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5920) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24467) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10572) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19842) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6687) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12194) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22684) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13109) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7660) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15192) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18174) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25205) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32093) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12534) * $signed(input_fmap_91[7:0]) +
	( 10'sd 335) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24116) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26022) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5338) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3531) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22655) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13754) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8424) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6170) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5800) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4701) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3432) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28071) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5088) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12537) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4313) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7748) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13721) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18310) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26893) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11733) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3954) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4516) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20681) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19208) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28682) * $signed(input_fmap_119[7:0]) +
	( 11'sd 911) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9011) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5289) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20979) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18916) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3135) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12926) * $signed(input_fmap_126[7:0]) +
	( 9'sd 219) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 14'sd 4538) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31911) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11054) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23673) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2081) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7122) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17031) * $signed(input_fmap_8[7:0]) +
	( 10'sd 258) * $signed(input_fmap_9[7:0]) +
	( 14'sd 8176) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13367) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1396) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25364) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12439) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17244) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16238) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4129) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14063) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21660) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9455) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32608) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20822) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22732) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25986) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19486) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20695) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30268) * $signed(input_fmap_32[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10984) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25324) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32008) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6981) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11338) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25357) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23310) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14984) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18339) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3040) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7643) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10797) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6344) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8963) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17379) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24145) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21499) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2998) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3605) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24499) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23955) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4764) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30408) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10944) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22815) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24323) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27814) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17555) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6441) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23847) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31850) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7581) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17527) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10508) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19587) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16338) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13322) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27732) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27587) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1430) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25890) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25110) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20817) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24131) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9835) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30844) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27704) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3358) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22844) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28114) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18556) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26275) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14973) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12713) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21767) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7452) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31204) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19960) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28640) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11759) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25371) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6031) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21305) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14162) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28251) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22228) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21124) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23950) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3818) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30377) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26147) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17540) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5641) * $signed(input_fmap_110[7:0]) +
	( 10'sd 304) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20447) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9270) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26227) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1964) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29698) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19434) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6599) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6652) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19403) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7617) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15750) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2431) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25918) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18881) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9418) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 12'sd 1481) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4208) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14682) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2080) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27999) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27526) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29797) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13505) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6705) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32552) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14773) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22498) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2898) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14733) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12430) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19829) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15182) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16487) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21002) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2298) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3356) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21137) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19500) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20213) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22772) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25573) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3277) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10202) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2157) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13257) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5917) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19146) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14012) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14564) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4466) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5285) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4271) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16685) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24838) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32715) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14211) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30426) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11786) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27714) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21986) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2338) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21535) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22310) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5170) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28064) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23383) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31509) * $signed(input_fmap_59[7:0]) +
	( 11'sd 1003) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26667) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16020) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10118) * $signed(input_fmap_64[7:0]) +
	( 10'sd 414) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21310) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8600) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16171) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17952) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4909) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23130) * $signed(input_fmap_71[7:0]) +
	( 11'sd 655) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19992) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8565) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32500) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23878) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22505) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22878) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26802) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15523) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14235) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24580) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24998) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2191) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20286) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20371) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19903) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23159) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4648) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29351) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13536) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2648) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32266) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29570) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15646) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24640) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15156) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31000) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14620) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13327) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17020) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28063) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19241) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17655) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28532) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11898) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1266) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4591) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4517) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19438) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24303) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29769) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18508) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30758) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9654) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7765) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13783) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28649) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7382) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24064) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2443) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 15'sd 16172) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30910) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16992) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_3[7:0]) +
	( 10'sd 349) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4888) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13565) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22952) * $signed(input_fmap_7[7:0]) +
	( 11'sd 610) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1257) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1498) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28067) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5045) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25722) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8758) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13603) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7387) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7250) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3521) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29721) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6672) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26284) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18553) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6479) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5177) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11599) * $signed(input_fmap_25[7:0]) +
	( 14'sd 8169) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21521) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24169) * $signed(input_fmap_28[7:0]) +
	( 9'sd 137) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3126) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4783) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1070) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9121) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4229) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14414) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14167) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23562) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15525) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21628) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30707) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23975) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32498) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9391) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9236) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5799) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14613) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7149) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12808) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8768) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32729) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7894) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12508) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22481) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27518) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28765) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32695) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7701) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22103) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4742) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22122) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15349) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2919) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29824) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20795) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20624) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11780) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28133) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13495) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6944) * $signed(input_fmap_75[7:0]) +
	( 11'sd 827) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20401) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6805) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22773) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16871) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26926) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16603) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6175) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30479) * $signed(input_fmap_84[7:0]) +
	( 13'sd 4017) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16453) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10916) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8639) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30221) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3931) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28790) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11647) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11994) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22213) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11110) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25731) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25616) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16461) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13659) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3909) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12759) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9096) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22906) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28360) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18779) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9305) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32495) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26077) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6524) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14370) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13118) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30103) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16909) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16266) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26561) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6043) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12943) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24724) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12689) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26409) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9905) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3450) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6197) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 16'sd 16932) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19119) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20490) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13995) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1054) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27161) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25397) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32033) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6237) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7919) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12326) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21606) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8791) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14249) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1500) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1139) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30472) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18092) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10954) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7087) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12822) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19166) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29952) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21768) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10109) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6491) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13439) * $signed(input_fmap_32[7:0]) +
	( 10'sd 429) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19289) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7210) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25046) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22625) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14027) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12204) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31061) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23296) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11689) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27801) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6412) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20268) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11798) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8872) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28523) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13555) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25013) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26316) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21028) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6402) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9922) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18445) * $signed(input_fmap_58[7:0]) +
	( 14'sd 8135) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5268) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26412) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7023) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32458) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15422) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21875) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18092) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11263) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22060) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27219) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12937) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11242) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15008) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24709) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19569) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24928) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31930) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21218) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4464) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15062) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29607) * $signed(input_fmap_84[7:0]) +
	( 9'sd 236) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26928) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16815) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29818) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17079) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21629) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11744) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26571) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26788) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18252) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21997) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32702) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19400) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32433) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18313) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12706) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29485) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11776) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7636) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10166) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24956) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20179) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1334) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24118) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8689) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10494) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18879) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1268) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14690) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8933) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23860) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3407) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19714) * $signed(input_fmap_119[7:0]) +
	( 11'sd 752) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5635) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5751) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30151) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11461) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21898) * $signed(input_fmap_126[7:0]) +
	( 11'sd 884) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 14'sd 5125) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29002) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11776) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13453) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32027) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9563) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2463) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22900) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23869) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13359) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5212) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13691) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23962) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18918) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2385) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14652) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6079) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24138) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14047) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9053) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16317) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3243) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22253) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20217) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11159) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15067) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15905) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2295) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20140) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6138) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27490) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16543) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7334) * $signed(input_fmap_33[7:0]) +
	( 8'sd 104) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15923) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32624) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14375) * $signed(input_fmap_38[7:0]) +
	( 11'sd 947) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15319) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18082) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21272) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14529) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2755) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14716) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10921) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27854) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1965) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19900) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21849) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3359) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4644) * $signed(input_fmap_57[7:0]) +
	( 10'sd 366) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4952) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3900) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8997) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28119) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4781) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29086) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11898) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28979) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1971) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7773) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32625) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15202) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7489) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31499) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29458) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6702) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8735) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6767) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17657) * $signed(input_fmap_77[7:0]) +
	( 10'sd 308) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6593) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11961) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13608) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11138) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13260) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10978) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10700) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25377) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20625) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7563) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31672) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12423) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12591) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12940) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3004) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6008) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20354) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1795) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5064) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2129) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2443) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31907) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20558) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9803) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4794) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21623) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29140) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20435) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15936) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25755) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27899) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23311) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6690) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7223) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22888) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27130) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23300) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30500) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23016) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2161) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6009) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20130) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1643) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24484) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21786) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4618) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12144) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 14'sd 5032) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6059) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15862) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14374) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5314) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1577) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8673) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3941) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10264) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12005) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29850) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31054) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30688) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24739) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30840) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30703) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20069) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27478) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30333) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15626) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14471) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12969) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31931) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21841) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8257) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32257) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3285) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30280) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17240) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21770) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12009) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32179) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18209) * $signed(input_fmap_34[7:0]) +
	( 8'sd 74) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17384) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29025) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27536) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32342) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11927) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31009) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16966) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5442) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22226) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2506) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10040) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25241) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23354) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13811) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32112) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18085) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17887) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3312) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14941) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20965) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22049) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10405) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6361) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15896) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24539) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19430) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18606) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25036) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3794) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8242) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8434) * $signed(input_fmap_76[7:0]) +
	( 10'sd 394) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30733) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10339) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21483) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25911) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13065) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2714) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3207) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26207) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17999) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7110) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20764) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5465) * $signed(input_fmap_91[7:0]) +
	( 11'sd 911) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32717) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5150) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30350) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26935) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12889) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3898) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16716) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21656) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32501) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28446) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19920) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28506) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19921) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11619) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14623) * $signed(input_fmap_109[7:0]) +
	( 11'sd 981) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21812) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10527) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28823) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29792) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12516) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6356) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_118[7:0]) +
	( 10'sd 288) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1255) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2936) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15888) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8432) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5004) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6476) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22650) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 16'sd 20624) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22349) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3279) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14941) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19404) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10301) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20128) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5314) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3970) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14478) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12955) * $signed(input_fmap_10[7:0]) +
	( 15'sd 16320) * $signed(input_fmap_11[7:0]) +
	( 11'sd 966) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22542) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17397) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17871) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23607) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24918) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11549) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18820) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12964) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2351) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4584) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24655) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16316) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21714) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21502) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17013) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4587) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27808) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4562) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17626) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21275) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16388) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4805) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3040) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16201) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23056) * $signed(input_fmap_39[7:0]) +
	( 8'sd 81) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14461) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27485) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15196) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22896) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3091) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7521) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12265) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9305) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21325) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6065) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15437) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25676) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28825) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10672) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25138) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13247) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3271) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22758) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6694) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12242) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26938) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27036) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26174) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1843) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25727) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1637) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12996) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22421) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20512) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27259) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20570) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5856) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5273) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6890) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24430) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5318) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28860) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19005) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24146) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14391) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16614) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3702) * $signed(input_fmap_86[7:0]) +
	( 7'sd 55) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7175) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13902) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14584) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13214) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31234) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30141) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28230) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1516) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8612) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17201) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1641) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18615) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10284) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7565) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9541) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17277) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1059) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12997) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6521) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11689) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5417) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20208) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19173) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28802) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4591) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21608) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26210) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10758) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20441) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4531) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16699) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25089) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8487) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26871) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 11'sd 848) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26699) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23998) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13980) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30034) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6613) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9240) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17784) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13773) * $signed(input_fmap_9[7:0]) +
	( 14'sd 8030) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31126) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30691) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5445) * $signed(input_fmap_13[7:0]) +
	( 9'sd 183) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22462) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19225) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7873) * $signed(input_fmap_17[7:0]) +
	( 11'sd 634) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26682) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8689) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2190) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1310) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8879) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11321) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4581) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18810) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8352) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16756) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32411) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1373) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12936) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25944) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6153) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9169) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32645) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16939) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21422) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4806) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30538) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13105) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13352) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2694) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24817) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29576) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1073) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21075) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10044) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22624) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13805) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22877) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26458) * $signed(input_fmap_56[7:0]) +
	( 8'sd 74) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7364) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30878) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4924) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9489) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14991) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10056) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9072) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11225) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30637) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8456) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4396) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4928) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1137) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4889) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_72[7:0]) +
	( 9'sd 212) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3647) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18860) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22948) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12402) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1397) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21453) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32644) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8798) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29911) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29899) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24791) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20565) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14026) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16918) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28963) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4666) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11875) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20151) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14951) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14505) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16010) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9104) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23745) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28389) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13137) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7383) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30595) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26867) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26033) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15426) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2689) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14437) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21151) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30968) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12703) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7683) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15859) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10398) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14033) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7315) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30623) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28296) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29254) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10278) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8531) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26986) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17307) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12586) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27254) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13814) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 16'sd 17872) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24361) * $signed(input_fmap_1[7:0]) +
	( 11'sd 812) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1259) * $signed(input_fmap_3[7:0]) +
	( 14'sd 8020) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22663) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31275) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3121) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10268) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8792) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14276) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31202) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21859) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15627) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3898) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19568) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16787) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16032) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14306) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21259) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28728) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24868) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20968) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29421) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11329) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30096) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23189) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20916) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25953) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21837) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3632) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24287) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28752) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1856) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24051) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6680) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23127) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19891) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2193) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17208) * $signed(input_fmap_41[7:0]) +
	( 13'sd 4087) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24366) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13705) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2811) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23664) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14604) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11166) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26165) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21030) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18579) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26558) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2581) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12599) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12820) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25991) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18644) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13191) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11133) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3464) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4510) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7416) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1686) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19442) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11403) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12672) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1411) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14611) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19471) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7658) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22783) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17446) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2366) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32100) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16849) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5248) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32509) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20168) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31980) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7988) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27678) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27783) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6533) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9705) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24214) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10175) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_96[7:0]) +
	( 13'sd 4001) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24852) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6953) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15356) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8198) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19423) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11383) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12890) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23320) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24761) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29046) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5091) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5118) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16735) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8233) * $signed(input_fmap_111[7:0]) +
	( 11'sd 1011) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30349) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16499) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30722) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20333) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13790) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29403) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26162) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1844) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1137) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4371) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11818) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32592) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 15'sd 9705) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24544) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10900) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25752) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6188) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2198) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32167) * $signed(input_fmap_6[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29948) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4639) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28636) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13588) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6649) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29609) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24777) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6437) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21120) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10115) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25879) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26312) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13823) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26970) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22438) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14667) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12021) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11744) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6085) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28394) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21351) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9833) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13763) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10728) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8674) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5101) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1149) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7940) * $signed(input_fmap_39[7:0]) +
	( 11'sd 804) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22757) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7027) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11015) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23030) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25946) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10312) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26290) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1156) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19182) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24029) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8588) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2365) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17773) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30372) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11603) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15638) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14913) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2146) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11509) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32423) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1632) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16272) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12512) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23739) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19864) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4914) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22629) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23325) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20499) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17018) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17129) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31450) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9887) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7780) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2786) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10586) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4292) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20754) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30277) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14755) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11921) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3855) * $signed(input_fmap_89[7:0]) +
	( 11'sd 970) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2365) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19880) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17890) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15804) * $signed(input_fmap_95[7:0]) +
	( 14'sd 8062) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20173) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18655) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13935) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19089) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16191) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8514) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5335) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19046) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17466) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9749) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7087) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30248) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32398) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10385) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23937) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26706) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20590) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27331) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9971) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14379) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24275) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27934) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24972) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_120[7:0]) +
	( 6'sd 23) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5872) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13729) * $signed(input_fmap_123[7:0]) +
	( 13'sd 4060) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3570) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31480) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 16'sd 17054) * $signed(input_fmap_0[7:0]) +
	( 12'sd 2031) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6928) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7033) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13157) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6034) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26813) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14721) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12335) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2517) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28671) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6712) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30179) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17544) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17041) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23528) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1920) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3964) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15896) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25999) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21124) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32437) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15738) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7485) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10420) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8556) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28319) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28360) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13070) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4335) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30574) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18694) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32285) * $signed(input_fmap_34[7:0]) +
	( 11'sd 711) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8713) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16660) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19207) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20193) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21605) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19245) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18419) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1041) * $signed(input_fmap_43[7:0]) +
	( 11'sd 984) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6645) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2357) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31246) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25688) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17449) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14207) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4248) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1598) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3042) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30348) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10977) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4874) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28296) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3998) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5596) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9586) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3219) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12665) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9822) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3737) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5458) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19722) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25965) * $signed(input_fmap_68[7:0]) +
	( 10'sd 378) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14138) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6802) * $signed(input_fmap_71[7:0]) +
	( 9'sd 148) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30140) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27534) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8950) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22629) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23555) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22254) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15244) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31648) * $signed(input_fmap_80[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17442) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1326) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24977) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16776) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22701) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28968) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31559) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18006) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10052) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32602) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22162) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18937) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10818) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5906) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30387) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10333) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6015) * $signed(input_fmap_100[7:0]) +
	( 8'sd 106) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10308) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25784) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14444) * $signed(input_fmap_104[7:0]) +
	( 14'sd 8155) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29532) * $signed(input_fmap_106[7:0]) +
	( 9'sd 175) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31784) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6609) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13153) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14138) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26682) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9771) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30450) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12093) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27392) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12640) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9364) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13568) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25964) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22201) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26923) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23489) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14103) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 16'sd 23229) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31340) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4855) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10966) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12957) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27469) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7850) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9530) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1781) * $signed(input_fmap_10[7:0]) +
	( 15'sd 16290) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14384) * $signed(input_fmap_12[7:0]) +
	( 11'sd 628) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15599) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30920) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31056) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12629) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_18[7:0]) +
	( 10'sd 362) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29011) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29084) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6397) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28646) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27246) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17958) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30476) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5475) * $signed(input_fmap_27[7:0]) +
	( 10'sd 450) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19459) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6768) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26752) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28070) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11524) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2866) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19948) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32265) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9674) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1439) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2415) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25624) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6487) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13672) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15675) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6842) * $signed(input_fmap_44[7:0]) +
	( 11'sd 915) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10260) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31171) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22969) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30645) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_50[7:0]) +
	( 7'sd 34) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24631) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30307) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25083) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11667) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5655) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16850) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15966) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10026) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8558) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3005) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27285) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19242) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29718) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23489) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3930) * $signed(input_fmap_70[7:0]) +
	( 10'sd 455) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5964) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13018) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16395) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27942) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16936) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28354) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8945) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14910) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32518) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12531) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21834) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10944) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29122) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9590) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29936) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19125) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3150) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32056) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24792) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5376) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31637) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27261) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18657) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5584) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3244) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15377) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31866) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5852) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10285) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7363) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5559) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8396) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11504) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11167) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17329) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2755) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21053) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6061) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24366) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2288) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21175) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4110) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5340) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17848) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2459) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15011) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27066) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13518) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20550) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 12'sd 1748) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25816) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4252) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27391) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19759) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22518) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3986) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23772) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9323) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28258) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10327) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20335) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1618) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24825) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12825) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20602) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20795) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29129) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4159) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18049) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19055) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24821) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30834) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26283) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32398) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12191) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25080) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4366) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14641) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6839) * $signed(input_fmap_35[7:0]) +
	( 11'sd 971) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7020) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9790) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31049) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14397) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14211) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1545) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11056) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11260) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11144) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30914) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4858) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24777) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29999) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22652) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22007) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8491) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21121) * $signed(input_fmap_55[7:0]) +
	( 13'sd 4013) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29910) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12563) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13980) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18929) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12819) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27295) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27794) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4466) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22694) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1881) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18604) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1394) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14186) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29899) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22286) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16016) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8508) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11391) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26084) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25800) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29119) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23134) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21427) * $signed(input_fmap_87[7:0]) +
	( 10'sd 426) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19637) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8518) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5523) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31047) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22608) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6767) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30422) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15179) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24818) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31671) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5762) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6033) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1643) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27100) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2590) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10792) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24065) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26010) * $signed(input_fmap_111[7:0]) +
	( 16'sd 16902) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22480) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2384) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26685) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13778) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13173) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32346) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19706) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28071) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25718) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4566) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20694) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10145) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28152) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 16'sd 24343) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2167) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12398) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11099) * $signed(input_fmap_4[7:0]) +
	( 14'sd 8092) * $signed(input_fmap_5[7:0]) +
	( 11'sd 548) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20377) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10931) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13051) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26021) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4156) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17043) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17385) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4484) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31712) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5561) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22566) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12308) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29572) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19267) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14518) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21020) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1035) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24513) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28855) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11162) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15480) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27596) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27698) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13494) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29079) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6826) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27268) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11078) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29424) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3521) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30451) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22409) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18683) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7675) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29496) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3294) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11006) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25024) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26265) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2258) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21925) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9252) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14394) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12277) * $signed(input_fmap_59[7:0]) +
	( 10'sd 413) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11547) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19838) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6866) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17428) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3972) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31961) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32731) * $signed(input_fmap_69[7:0]) +
	( 7'sd 62) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30780) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14887) * $signed(input_fmap_73[7:0]) +
	( 11'sd 830) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18625) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7083) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25195) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13275) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20418) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24119) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17385) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3940) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9918) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13916) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2399) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19639) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25669) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22579) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31360) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32364) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27617) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3365) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10478) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17128) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32477) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30560) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23218) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2080) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9849) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18481) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23008) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5986) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5525) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19840) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20734) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5777) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13896) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24404) * $signed(input_fmap_114[7:0]) +
	( 16'sd 29366) * $signed(input_fmap_115[7:0]) +
	( 7'sd 43) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2995) * $signed(input_fmap_117[7:0]) +
	( 14'sd 8091) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30975) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10313) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30424) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24520) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21354) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30883) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27657) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 16'sd 21165) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21160) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9642) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2893) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18930) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29861) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28540) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25069) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27876) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2700) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2544) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14926) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7867) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4363) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30703) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7164) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28758) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22648) * $signed(input_fmap_19[7:0]) +
	( 10'sd 370) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16859) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6434) * $signed(input_fmap_22[7:0]) +
	( 11'sd 631) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16191) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32530) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10343) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21727) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24122) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6177) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29572) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21382) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14621) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26062) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29293) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26075) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2610) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27105) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6944) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17447) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29114) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14912) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9375) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20989) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2525) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12138) * $signed(input_fmap_49[7:0]) +
	( 10'sd 432) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24342) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11182) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1613) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3456) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29773) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21374) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32631) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18082) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2891) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1994) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6739) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12860) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24312) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26358) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3045) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8948) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11514) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11824) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31384) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7511) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17628) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28701) * $signed(input_fmap_77[7:0]) +
	( 10'sd 446) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24758) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15056) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19161) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30999) * $signed(input_fmap_83[7:0]) +
	( 8'sd 72) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8673) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18976) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27823) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16043) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30201) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16864) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25788) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9839) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1595) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10710) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9830) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18184) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1586) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1892) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32034) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3728) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21027) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_105[7:0]) +
	( 15'sd 16265) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24581) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15529) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30311) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8653) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25889) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26113) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23653) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16128) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6361) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24374) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5457) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30164) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6874) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4580) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8684) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18525) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1415) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25851) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3075) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4258) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20128) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 16'sd 31949) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32621) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30989) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9298) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10918) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12292) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28382) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19306) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8691) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17236) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6087) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19215) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5016) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31264) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17880) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15534) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14872) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31664) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4594) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27509) * $signed(input_fmap_21[7:0]) +
	( 6'sd 19) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7117) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15168) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14766) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32352) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29183) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28894) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25565) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1716) * $signed(input_fmap_30[7:0]) +
	( 11'sd 548) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26421) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28016) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27712) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30509) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7994) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3612) * $signed(input_fmap_37[7:0]) +
	( 9'sd 202) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17825) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28822) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8897) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18789) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32589) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8464) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22359) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24441) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24617) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16412) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29140) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1828) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16360) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11696) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19204) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27295) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27193) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29982) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31211) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4461) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13093) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14470) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21468) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14903) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3043) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18424) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6331) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9755) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2113) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6531) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18837) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2095) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27522) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23200) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18492) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18875) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6940) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18164) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16094) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26470) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4362) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17530) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22557) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22755) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24859) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27559) * $signed(input_fmap_92[7:0]) +
	( 11'sd 716) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13836) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28303) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10552) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7164) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12348) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1774) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11984) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5726) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30176) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6656) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28622) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3867) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3180) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24485) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18593) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10710) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9455) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30495) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20572) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31238) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30944) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26757) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23817) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8702) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15328) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4844) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10858) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31534) * $signed(input_fmap_124[7:0]) +
	( 10'sd 500) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11395) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 16'sd 21652) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1874) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1097) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11593) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13317) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31469) * $signed(input_fmap_5[7:0]) +
	( 11'sd 812) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13934) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5188) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10416) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5883) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29055) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11120) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4669) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4577) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9194) * $signed(input_fmap_17[7:0]) +
	( 14'sd 8062) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27832) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18039) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11604) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2819) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27575) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27454) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30648) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30541) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6829) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4826) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12939) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30957) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30509) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29313) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2982) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32264) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9169) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16410) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7425) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22310) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3768) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30190) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5818) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22838) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13575) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17021) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10405) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27883) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5457) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6870) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16405) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27495) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24794) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27487) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9681) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4896) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13388) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9649) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28043) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8336) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29347) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19237) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17135) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30046) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25325) * $signed(input_fmap_67[7:0]) +
	( 7'sd 51) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20583) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9919) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9833) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21008) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27667) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21316) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8774) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2164) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5101) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23610) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19953) * $signed(input_fmap_85[7:0]) +
	( 14'sd 8005) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16523) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7024) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22765) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20775) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23135) * $signed(input_fmap_91[7:0]) +
	( 9'sd 168) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14838) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4640) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2435) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4962) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3540) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26256) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18215) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25533) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9310) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31538) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32102) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11716) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13912) * $signed(input_fmap_106[7:0]) +
	( 8'sd 111) * $signed(input_fmap_107[7:0]) +
	( 11'sd 561) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27204) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11751) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20503) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1746) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1435) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22827) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25969) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23693) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10981) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32622) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18070) * $signed(input_fmap_121[7:0]) +
	( 11'sd 915) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14268) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1468) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30085) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5047) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 15'sd 15823) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2309) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18020) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3135) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15076) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3988) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13539) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3916) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15319) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31907) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14995) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30761) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25184) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17925) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9500) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12860) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25780) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25934) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29064) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2218) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1857) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24730) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15084) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23522) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16746) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14461) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23802) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9634) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23781) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31618) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27439) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2363) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29125) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32222) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12615) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6689) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23945) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31741) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21847) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10996) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30366) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2401) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1849) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8409) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30698) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31306) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1773) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2161) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15510) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31002) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6431) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11994) * $signed(input_fmap_57[7:0]) +
	( 11'sd 689) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14093) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9764) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6194) * $signed(input_fmap_61[7:0]) +
	( 11'sd 658) * $signed(input_fmap_62[7:0]) +
	( 11'sd 930) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30246) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9076) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27901) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8561) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27212) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9369) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31230) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30266) * $signed(input_fmap_71[7:0]) +
	( 14'sd 8103) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2992) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27860) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11107) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29680) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28737) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25758) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23918) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21505) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15117) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1320) * $signed(input_fmap_83[7:0]) +
	( 9'sd 162) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6888) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21138) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11485) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15032) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3955) * $signed(input_fmap_89[7:0]) +
	( 11'sd 665) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14531) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6499) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11258) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8193) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19122) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25791) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4767) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14575) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20531) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31898) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23336) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24620) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22794) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28674) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2174) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11272) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29245) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32074) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29110) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29915) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26441) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6753) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22322) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31762) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5385) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20788) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17139) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25175) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6213) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4825) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19104) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2745) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 16'sd 31031) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2954) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10730) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21873) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8748) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3444) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22585) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5165) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30633) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7105) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25668) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18844) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30807) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8242) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31854) * $signed(input_fmap_15[7:0]) +
	( 14'sd 8005) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25021) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7804) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16519) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22999) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9920) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4335) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15959) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18219) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18376) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4403) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21886) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29779) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22396) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16400) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6781) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21918) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3906) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28411) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30226) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13177) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32680) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30554) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18293) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24438) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23350) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2561) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26334) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15917) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16644) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20055) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9383) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19337) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15933) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25353) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18838) * $signed(input_fmap_53[7:0]) +
	( 10'sd 257) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8611) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22165) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_57[7:0]) +
	( 11'sd 934) * $signed(input_fmap_58[7:0]) +
	( 11'sd 694) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8656) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16156) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18632) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24116) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4109) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19782) * $signed(input_fmap_65[7:0]) +
	( 11'sd 588) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22971) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29831) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18848) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_70[7:0]) +
	( 11'sd 747) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32562) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10194) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31518) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28998) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24094) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14040) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21129) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22965) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20685) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4556) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10903) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17994) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30376) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8503) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32304) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7159) * $signed(input_fmap_88[7:0]) +
	( 11'sd 514) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11046) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29183) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25359) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21835) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22172) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28688) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31937) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22101) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8746) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21037) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22633) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20717) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8616) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14430) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21356) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23062) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23019) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29230) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10210) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19381) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7036) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25255) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16118) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31278) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_119[7:0]) +
	( 14'sd 8122) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27515) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11045) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9397) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32603) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32195) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18590) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23735) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 13'sd 2218) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26893) * $signed(input_fmap_1[7:0]) +
	( 10'sd 298) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6860) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9810) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22960) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9394) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29817) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3929) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32757) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3598) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15007) * $signed(input_fmap_12[7:0]) +
	( 10'sd 498) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17493) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7811) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4664) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25664) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28011) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12159) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27811) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18588) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30996) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12370) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25848) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18944) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22046) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6194) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14392) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9705) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23399) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22713) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5782) * $signed(input_fmap_34[7:0]) +
	( 12'sd 2021) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24626) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17036) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18221) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25120) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30878) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4634) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4363) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13138) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18262) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21012) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30675) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12254) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22528) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6004) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16014) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12247) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12439) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28863) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11805) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8594) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31969) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10542) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11394) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12101) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13493) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31934) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10058) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1870) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27851) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24575) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3458) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17246) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15283) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20052) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6905) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1876) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3333) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24368) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9166) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10872) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29538) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20705) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1799) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16452) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6288) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27735) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7839) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10751) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25704) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23436) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9791) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5267) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4826) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20502) * $signed(input_fmap_101[7:0]) +
	( 13'sd 4074) * $signed(input_fmap_102[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21068) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10571) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17437) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7180) * $signed(input_fmap_109[7:0]) +
	( 9'sd 209) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12229) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21703) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11537) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10343) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15860) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7411) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7782) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28891) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6357) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7370) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1989) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9459) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14729) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2884) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21616) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21432) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 16'sd 30758) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26678) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12571) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9909) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10527) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15988) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4704) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28362) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30785) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13265) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7358) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23908) * $signed(input_fmap_12[7:0]) +
	( 15'sd 16343) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16533) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8348) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5713) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10708) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28400) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21006) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31824) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31160) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1757) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5282) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8227) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20172) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8545) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12561) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29286) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26827) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1161) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8751) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31895) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22047) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24574) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21780) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10973) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20917) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14596) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4882) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24536) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16120) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12387) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24774) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3381) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1580) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31474) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31958) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16498) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5859) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28964) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22957) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5359) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24038) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9397) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14854) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25436) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6571) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11177) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19320) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1246) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26976) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6357) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8675) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21125) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23500) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18127) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3525) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1357) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4873) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25831) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26982) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12222) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14014) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4162) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27370) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15672) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7400) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21453) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1110) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30257) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27880) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2976) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1164) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28527) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1542) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29724) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28461) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18870) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19287) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16997) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19276) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13299) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16858) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30452) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26364) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9313) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21287) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19175) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17642) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18252) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6527) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11610) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24629) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32348) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28457) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5554) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 16'sd 20397) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9214) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15804) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29876) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12078) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15815) * $signed(input_fmap_5[7:0]) +
	( 11'sd 527) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3976) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18977) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28279) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26595) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17678) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10818) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19428) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2833) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10068) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16793) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30824) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29584) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6703) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27497) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27016) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28349) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16710) * $signed(input_fmap_25[7:0]) +
	( 13'sd 4036) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11451) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18898) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12651) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5696) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27918) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31313) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30587) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13166) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7046) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20722) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8652) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32567) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9674) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3874) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24655) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12414) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30476) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20056) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5231) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12203) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7036) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9584) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22475) * $signed(input_fmap_50[7:0]) +
	( 10'sd 505) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26527) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15542) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29198) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5927) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23089) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27801) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8931) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8295) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16810) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19837) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23856) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13907) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5867) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26791) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8638) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28934) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4688) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8549) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11812) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2445) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28230) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29994) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8432) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10901) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20873) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32503) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3797) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15585) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8374) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19301) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19245) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23857) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27758) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19239) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24889) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30430) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23286) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17895) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22797) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28669) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18429) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16876) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6216) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10601) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23938) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12877) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8331) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16476) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13588) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16850) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27252) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19266) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10507) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15354) * $signed(input_fmap_116[7:0]) +
	( 10'sd 494) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17975) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5621) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14549) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18795) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7906) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12721) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13227) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3217) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20231) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28909) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 16'sd 16758) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14814) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18208) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1445) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22136) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23585) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5813) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31928) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13822) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2639) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20632) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15112) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26667) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27581) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6447) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10909) * $signed(input_fmap_16[7:0]) +
	( 9'sd 181) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7413) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27741) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8294) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26039) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22181) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16482) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16518) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13482) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28503) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22552) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28949) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1252) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27799) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16624) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19772) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13795) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26799) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5811) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9727) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12332) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32261) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2963) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2310) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13075) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17948) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20839) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28854) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16444) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13568) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12878) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30881) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21081) * $signed(input_fmap_52[7:0]) +
	( 9'sd 248) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23060) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8622) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28794) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1681) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7385) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16025) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26187) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28768) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28052) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29012) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23970) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21567) * $signed(input_fmap_70[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2518) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4286) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10266) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12430) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1208) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5372) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21542) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23198) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10090) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18242) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9824) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20464) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27713) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13729) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23724) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19742) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21192) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10574) * $signed(input_fmap_90[7:0]) +
	( 11'sd 915) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10494) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6041) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10323) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21109) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31227) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16761) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17005) * $signed(input_fmap_98[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6488) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14495) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4964) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27088) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27300) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27661) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5824) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13897) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31171) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31581) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12999) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20974) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8863) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6802) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22288) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19586) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8287) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15462) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8874) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28838) * $signed(input_fmap_120[7:0]) +
	( 11'sd 855) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24660) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20974) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6746) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28998) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15160) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8933) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 16'sd 21222) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31000) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18436) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27234) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17266) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2969) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10092) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24229) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16176) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26212) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3450) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4737) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11901) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23977) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26030) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16319) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13941) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27557) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24891) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23013) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28053) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11418) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7689) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8262) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8403) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17077) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4248) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16985) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26599) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24214) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26745) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13228) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6468) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25564) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22884) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19246) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15659) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2228) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3673) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10414) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2513) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25129) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22196) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7118) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32238) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32261) * $signed(input_fmap_47[7:0]) +
	( 10'sd 263) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32732) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9170) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3617) * $signed(input_fmap_51[7:0]) +
	( 14'sd 8012) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17739) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11002) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7484) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4620) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10094) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32129) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32722) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3410) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28087) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29294) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17670) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31312) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22700) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28720) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10323) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32585) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7655) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29855) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20218) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18570) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8717) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15945) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17356) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13358) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4656) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17458) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11955) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12712) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13807) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16394) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17368) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10000) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18022) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1825) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17081) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18736) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23431) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3616) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5989) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29725) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11831) * $signed(input_fmap_102[7:0]) +
	( 16'sd 32163) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14300) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32638) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16411) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17101) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20543) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4485) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8066) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2667) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25582) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11052) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32134) * $signed(input_fmap_117[7:0]) +
	( 11'sd 752) * $signed(input_fmap_118[7:0]) +
	( 10'sd 318) * $signed(input_fmap_119[7:0]) +
	( 11'sd 1004) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3656) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13215) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22656) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29571) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25328) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7929) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27693) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 15'sd 8570) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5318) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22228) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5780) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12208) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25801) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2629) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6880) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7006) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18215) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26311) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13618) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16369) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1282) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12493) * $signed(input_fmap_16[7:0]) +
	( 8'sd 126) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11070) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2692) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27730) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12282) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5996) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16737) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20246) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11911) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7590) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27870) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14756) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20126) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11645) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13366) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32105) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2125) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24681) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25591) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21238) * $signed(input_fmap_38[7:0]) +
	( 9'sd 253) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4815) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29616) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17876) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14380) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13277) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10924) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25851) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5011) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25245) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13667) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6899) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8434) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11453) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_53[7:0]) +
	( 10'sd 485) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10574) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22038) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27805) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8978) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9123) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2603) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14500) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10371) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2121) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21971) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15791) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19514) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11825) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6886) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30762) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3701) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6302) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13647) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1301) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14966) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13023) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21397) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19626) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14715) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24811) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14017) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3287) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22179) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22581) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31449) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31125) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23640) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19840) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16064) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14316) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28176) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30831) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4726) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15171) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12981) * $signed(input_fmap_96[7:0]) +
	( 11'sd 893) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8436) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24160) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16421) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25034) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13822) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11071) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29740) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16286) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12872) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31244) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13054) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18309) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25428) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4956) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15881) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6977) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26237) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7239) * $signed(input_fmap_118[7:0]) +
	( 15'sd 16259) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30596) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16470) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31740) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32634) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11562) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7635) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9665) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 15'sd 9510) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26183) * $signed(input_fmap_1[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26887) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6728) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12074) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29044) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1233) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20900) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9587) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27701) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5787) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32175) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9101) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26905) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27967) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12413) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23414) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6945) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7242) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12218) * $signed(input_fmap_22[7:0]) +
	( 14'sd 8150) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5264) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25390) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23400) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13240) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28738) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12685) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2410) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12876) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18763) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3075) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28143) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30806) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8432) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15780) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4916) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24388) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18669) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12737) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10487) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16274) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17684) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14375) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7970) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26510) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5280) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5055) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29658) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11270) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29754) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19620) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28359) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27592) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10112) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24788) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12008) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4198) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13156) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25195) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9561) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16037) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21908) * $signed(input_fmap_73[7:0]) +
	( 10'sd 265) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1064) * $signed(input_fmap_75[7:0]) +
	( 13'sd 4040) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27604) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3923) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9798) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32038) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15006) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12533) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1403) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28977) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9535) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10891) * $signed(input_fmap_90[7:0]) +
	( 10'sd 507) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2068) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20824) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28969) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14052) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8974) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20778) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8302) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29537) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19481) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24431) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10543) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7623) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12149) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7447) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24930) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14923) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13839) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15591) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3528) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31043) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24896) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23828) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16804) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26503) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20238) * $signed(input_fmap_119[7:0]) +
	( 10'sd 353) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26608) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19320) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31767) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3544) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9000) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6068) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20271) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 16'sd 17983) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24998) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19367) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23219) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23450) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14955) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13676) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14313) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3067) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13299) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2573) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30066) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6892) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13441) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22546) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24938) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1175) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24402) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2219) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3452) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12592) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13839) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15943) * $signed(input_fmap_28[7:0]) +
	( 13'sd 4031) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22924) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11605) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10924) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15082) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22344) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1384) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19341) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13699) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26677) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8699) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3505) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9923) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25465) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7093) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8650) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31728) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_51[7:0]) +
	( 13'sd 4090) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13704) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16541) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10506) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28680) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3454) * $signed(input_fmap_60[7:0]) +
	( 11'sd 944) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13883) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16727) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27934) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26983) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17889) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8419) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10216) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22692) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5503) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15199) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18762) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19372) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25470) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14381) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5631) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13658) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25236) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21670) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21897) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14466) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24507) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7339) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17460) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19468) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15841) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3703) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16921) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_93[7:0]) +
	( 9'sd 145) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17703) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27994) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26969) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29373) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19958) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19658) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_103[7:0]) +
	( 11'sd 673) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20058) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3713) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1089) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30159) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18123) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19718) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32331) * $signed(input_fmap_111[7:0]) +
	( 10'sd 266) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11636) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7665) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8810) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25794) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23241) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25999) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19959) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20996) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8562) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13690) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3214) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 11'sd 1002) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14154) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12700) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30571) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9798) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14585) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17726) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13277) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3946) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23651) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2723) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5000) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24206) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14962) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13833) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14290) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23940) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5062) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1456) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21877) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17017) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20684) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24724) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29919) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26900) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16581) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4950) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32015) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6969) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7621) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30171) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22527) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4409) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11513) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12674) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2310) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22284) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7355) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14905) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23971) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27610) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32275) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31110) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27813) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11662) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24808) * $signed(input_fmap_54[7:0]) +
	( 14'sd 8137) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31736) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15694) * $signed(input_fmap_57[7:0]) +
	( 10'sd 447) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15063) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32154) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8074) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26757) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13162) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17156) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29156) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12046) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25691) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23921) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1672) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30638) * $signed(input_fmap_70[7:0]) +
	( 9'sd 163) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9069) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27000) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29034) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17442) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2178) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27065) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24248) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29518) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13826) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29937) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3248) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29525) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23101) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29535) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26379) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30501) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27714) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31805) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8804) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22953) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5672) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30039) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11077) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6840) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13803) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8919) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29405) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23624) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31356) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14302) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16341) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7221) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16057) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12540) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8526) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22234) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32331) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25893) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27304) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7809) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8248) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16819) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10702) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6224) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8597) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31214) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24437) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9790) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9458) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 16'sd 24375) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18253) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16306) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12609) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14867) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26630) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7032) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21643) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22999) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13936) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24131) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27264) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3392) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23272) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26202) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19914) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25615) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23128) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11163) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9453) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11031) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1517) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10702) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6948) * $signed(input_fmap_26[7:0]) +
	( 8'sd 80) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4380) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3157) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4778) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8817) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4902) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21474) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5751) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19109) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28392) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23036) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9340) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20312) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14805) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6375) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7835) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15718) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29529) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32568) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4304) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7901) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5195) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9972) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29177) * $signed(input_fmap_52[7:0]) +
	( 11'sd 728) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3060) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23267) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17362) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23525) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5697) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31459) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27716) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28933) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22868) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16662) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25278) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1503) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23699) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18615) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32410) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24683) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27185) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6830) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4427) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31417) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29297) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24924) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25807) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5772) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10295) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28297) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18293) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4299) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21165) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27363) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26666) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32102) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20318) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6003) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8266) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8331) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30338) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8467) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1999) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22392) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21977) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4370) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7084) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16280) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17852) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26335) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15902) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26826) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20129) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15098) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13103) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2905) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29509) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26369) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3441) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4367) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18000) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6491) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14270) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6382) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29658) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31215) * $signed(input_fmap_125[7:0]) +
	( 11'sd 989) * $signed(input_fmap_126[7:0]) +
	( 11'sd 683) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 16'sd 30158) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3700) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16940) * $signed(input_fmap_2[7:0]) +
	( 13'sd 4065) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1085) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29440) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12844) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3273) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14596) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15297) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6710) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30634) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22054) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17320) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15863) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2203) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17985) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30965) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15771) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11469) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2111) * $signed(input_fmap_21[7:0]) +
	( 13'sd 4003) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12294) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18180) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11242) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30206) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26583) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5897) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15854) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15672) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13749) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16105) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12036) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24957) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16998) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5821) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22996) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20119) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22841) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1608) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16384) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31223) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16457) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11760) * $signed(input_fmap_49[7:0]) +
	( 14'sd 8058) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4322) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26879) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6798) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29659) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21256) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15370) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27229) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31334) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5634) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17413) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29789) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13540) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32302) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9746) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17096) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29901) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25554) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24106) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31458) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6543) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20024) * $signed(input_fmap_76[7:0]) +
	( 14'sd 8081) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17832) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26092) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25523) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28779) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15824) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18776) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32043) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20679) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9747) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5649) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1564) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7428) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21656) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16716) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10159) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32723) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17606) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15439) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11685) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5330) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21442) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22835) * $signed(input_fmap_100[7:0]) +
	( 11'sd 878) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4138) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24991) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12203) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5882) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28350) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27664) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5340) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30837) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21366) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24761) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26455) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24492) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26757) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27708) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1145) * $signed(input_fmap_117[7:0]) +
	( 8'sd 70) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25820) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30255) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3539) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24901) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5903) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17500) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25509) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 16'sd 29162) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15962) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2613) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24403) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20882) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23244) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7594) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3156) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26782) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7805) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21634) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2874) * $signed(input_fmap_12[7:0]) +
	( 6'sd 25) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7150) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3079) * $signed(input_fmap_15[7:0]) +
	( 10'sd 472) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16180) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16556) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29592) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18608) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16066) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13431) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18966) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15748) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22061) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23108) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10969) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8724) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7273) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7180) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26711) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12494) * $signed(input_fmap_35[7:0]) +
	( 11'sd 663) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14189) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16614) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6139) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12610) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22573) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15760) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24869) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15078) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23796) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17024) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12839) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5891) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10356) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5390) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10159) * $signed(input_fmap_56[7:0]) +
	( 10'sd 311) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15354) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17217) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32008) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28811) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19384) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10464) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16532) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15621) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14268) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15558) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20147) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26586) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31854) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27443) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6654) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5366) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20527) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32398) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19401) * $signed(input_fmap_81[7:0]) +
	( 9'sd 217) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5401) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15325) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15407) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27438) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3995) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23454) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14176) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32214) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24619) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6506) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26993) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17170) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8456) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29532) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28487) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30855) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25379) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5448) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17754) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1767) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11645) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4587) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6129) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1143) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17266) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24375) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14291) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10888) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29601) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13493) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4589) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1917) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10060) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17225) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14171) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19836) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26543) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13045) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12038) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24879) * $signed(input_fmap_126[7:0]) +
	( 9'sd 158) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 15'sd 9501) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29490) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23539) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21021) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18913) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25765) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5443) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1706) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9128) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14199) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9343) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16875) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20178) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29109) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12928) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24448) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10143) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3280) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16869) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4096) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8830) * $signed(input_fmap_21[7:0]) +
	( 10'sd 488) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14630) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2548) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29864) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2362) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27203) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20384) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6563) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8772) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9565) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32210) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20370) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29666) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25307) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8226) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25710) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16236) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10593) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6671) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13958) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14638) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4247) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30298) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24894) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1670) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7660) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24169) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19842) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30902) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25838) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4803) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17969) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29109) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30758) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25167) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19831) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28844) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16203) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13150) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15649) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32312) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12758) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5725) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31945) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9367) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15723) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23799) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27806) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10317) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19998) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7745) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31607) * $signed(input_fmap_80[7:0]) +
	( 11'sd 921) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29895) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32228) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13837) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27116) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10570) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14344) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22099) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22771) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3373) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28362) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23268) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28208) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26201) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5103) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22909) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17209) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8544) * $signed(input_fmap_102[7:0]) +
	( 11'sd 972) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8575) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27892) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30894) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32284) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1096) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32379) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23391) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29889) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31857) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8980) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18211) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32258) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26197) * $signed(input_fmap_120[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_121[7:0]) +
	( 13'sd 4019) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20365) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11607) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2176) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2205) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_127[7:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 16'sd 21033) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20741) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25335) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24143) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17047) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12318) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12837) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12041) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9379) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28038) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31474) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27125) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4418) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25259) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5714) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15380) * $signed(input_fmap_16[7:0]) +
	( 11'sd 676) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4826) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18061) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9786) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17755) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19484) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31812) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2739) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5462) * $signed(input_fmap_26[7:0]) +
	( 15'sd 16063) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23811) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27752) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15002) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29750) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1218) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21606) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21980) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14586) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17702) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25075) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15076) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13994) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16746) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22895) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21978) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8080) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12247) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27405) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16678) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6343) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19129) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20817) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16297) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28510) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6047) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7380) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21379) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13336) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27004) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26586) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7872) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19607) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15200) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19324) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27041) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13156) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2780) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7475) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_72[7:0]) +
	( 9'sd 173) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12273) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4578) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15719) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25319) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18921) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25356) * $signed(input_fmap_80[7:0]) +
	( 11'sd 894) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25072) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26066) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28675) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1173) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3358) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4357) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12362) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27568) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13361) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23997) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16395) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18390) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10898) * $signed(input_fmap_95[7:0]) +
	( 9'sd 137) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28763) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13218) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25617) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15277) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25353) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5415) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18632) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17324) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4837) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27394) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13207) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26316) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13038) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12576) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21374) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5725) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5791) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3081) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20912) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31816) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25942) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3537) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31407) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15180) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27641) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7008) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30408) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_127[7:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 16'd23080;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 16'd19266;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 16'd24591;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 16'd30231;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 15'd10405;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 11'd624;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 16'd24594;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 16'd22158;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 13'd2751;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 14'd8026;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 15'd15454;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 16'd30229;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 16'd27960;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 15'd15613;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 16'd18033;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 16'd26793;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 13'd2408;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 15'd10062;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 16'd16964;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 14'd4464;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 13'd2947;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 16'd20624;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 16'd26741;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 13'd2187;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 16'd29887;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 15'd15695;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 16'd25391;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 16'd28097;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 12'd1186;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 15'd10474;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 15'd15755;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 15'd14170;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 9'd172;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 16'd25676;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 16'd17415;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 16'd29628;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 13'd2696;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 16'd23754;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 15'd10455;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 10'd401;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 16'd27509;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 11'd642;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 12'd1616;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 16'd17650;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 16'd19970;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 14'd8087;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 16'd21939;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 16'd21987;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 13'd3555;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 16'd25647;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 16'd29285;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 16'd20867;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 16'd21711;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 15'd14935;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 15'd11173;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 15'd8775;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 16'd28172;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 16'd32168;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 16'd31227;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 16'd20869;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 16'd25749;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 14'd7783;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 16'd27482;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 15'd12494;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64 + 15'd11078;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 16'd20179;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 16'd27998;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67 + 16'd21306;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 16'd28934;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 16'd22995;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 15'd8833;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 15'd12784;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 15'd9316;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 12'd1940;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74 + 16'd24555;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 16'd21532;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 16'd22490;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 15'd13103;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 15'd13132;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79 + 16'd22977;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80 + 16'd27003;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81 + 16'd29814;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 16'd32612;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 14'd5217;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 14'd5370;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 16'd22646;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 14'd7901;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 16'd27573;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 15'd13077;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 13'd3200;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 14'd7834;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91 + 14'd4966;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 16'd26902;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 15'd15925;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 15'd13493;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 15'd9414;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 14'd7346;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97 + 16'd18621;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 16'd20223;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 4'd6;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 16'd30865;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 14'd5766;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102 + 16'd32742;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 15'd13891;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 15'd9579;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 15'd8941;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 16'd24492;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 14'd6340;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108 + 16'd27789;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 16'd32203;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 15'd16193;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 16'd16500;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 16'd21529;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113 + 16'd19967;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 16'd21314;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 16'd22674;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116 + 15'd16006;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117 + 14'd5544;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 12'd1129;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 16'd20176;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 16'd17077;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 10'd258;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 15'd15369;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 16'd22162;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124 + 15'd15924;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 13'd3910;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 15'd14912;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 16'd21695;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[21:15]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[21:15]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[21:15]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[21:15]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[21:15]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[21:15]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[21:15]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[21:15]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[21:15]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[21:15]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[21:15]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[21:15]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[21:15]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[21:15]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[21:15]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[21:15]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[21:15]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[21:15]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[21:15]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[21:15]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[21:15]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[21:15]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[21:15]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[21:15]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[21:15]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[21:15]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[21:15]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[21:15]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[21:15]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[21:15]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[21:15]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[21:15]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[21:15]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[21:15]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[21:15]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[21:15]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[21:15]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[21:15]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[21:15]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[21:15]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[21:15]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[21:15]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[21:15]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[21:15]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[21:15]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[21:15]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[21:15]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[21:15]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[21:15]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[21:15]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[21:15]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[21:15]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[21:15]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[21:15]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[21:15]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[21:15]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[21:15]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[21:15]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[21:15]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[21:15]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[21:15]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[21:15]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[21:15]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[21:15]}} :'d6) : '0;
logic [7:0] relu_64;
assign relu_64[7:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[21:15]}} :'d6) : '0;
logic [7:0] relu_65;
assign relu_65[7:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[21:15]}} :'d6) : '0;
logic [7:0] relu_66;
assign relu_66[7:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[21:15]}} :'d6) : '0;
logic [7:0] relu_67;
assign relu_67[7:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[21:15]}} :'d6) : '0;
logic [7:0] relu_68;
assign relu_68[7:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[21:15]}} :'d6) : '0;
logic [7:0] relu_69;
assign relu_69[7:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[21:15]}} :'d6) : '0;
logic [7:0] relu_70;
assign relu_70[7:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[21:15]}} :'d6) : '0;
logic [7:0] relu_71;
assign relu_71[7:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[21:15]}} :'d6) : '0;
logic [7:0] relu_72;
assign relu_72[7:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[21:15]}} :'d6) : '0;
logic [7:0] relu_73;
assign relu_73[7:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[21:15]}} :'d6) : '0;
logic [7:0] relu_74;
assign relu_74[7:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[21:15]}} :'d6) : '0;
logic [7:0] relu_75;
assign relu_75[7:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[21:15]}} :'d6) : '0;
logic [7:0] relu_76;
assign relu_76[7:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[21:15]}} :'d6) : '0;
logic [7:0] relu_77;
assign relu_77[7:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[21:15]}} :'d6) : '0;
logic [7:0] relu_78;
assign relu_78[7:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[21:15]}} :'d6) : '0;
logic [7:0] relu_79;
assign relu_79[7:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[21:15]}} :'d6) : '0;
logic [7:0] relu_80;
assign relu_80[7:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[21:15]}} :'d6) : '0;
logic [7:0] relu_81;
assign relu_81[7:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[21:15]}} :'d6) : '0;
logic [7:0] relu_82;
assign relu_82[7:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[21:15]}} :'d6) : '0;
logic [7:0] relu_83;
assign relu_83[7:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[21:15]}} :'d6) : '0;
logic [7:0] relu_84;
assign relu_84[7:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[21:15]}} :'d6) : '0;
logic [7:0] relu_85;
assign relu_85[7:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[21:15]}} :'d6) : '0;
logic [7:0] relu_86;
assign relu_86[7:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[21:15]}} :'d6) : '0;
logic [7:0] relu_87;
assign relu_87[7:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[21:15]}} :'d6) : '0;
logic [7:0] relu_88;
assign relu_88[7:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[21:15]}} :'d6) : '0;
logic [7:0] relu_89;
assign relu_89[7:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[21:15]}} :'d6) : '0;
logic [7:0] relu_90;
assign relu_90[7:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[21:15]}} :'d6) : '0;
logic [7:0] relu_91;
assign relu_91[7:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[21:15]}} :'d6) : '0;
logic [7:0] relu_92;
assign relu_92[7:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[21:15]}} :'d6) : '0;
logic [7:0] relu_93;
assign relu_93[7:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[21:15]}} :'d6) : '0;
logic [7:0] relu_94;
assign relu_94[7:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[21:15]}} :'d6) : '0;
logic [7:0] relu_95;
assign relu_95[7:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[21:15]}} :'d6) : '0;
logic [7:0] relu_96;
assign relu_96[7:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[21:15]}} :'d6) : '0;
logic [7:0] relu_97;
assign relu_97[7:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[21:15]}} :'d6) : '0;
logic [7:0] relu_98;
assign relu_98[7:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[21:15]}} :'d6) : '0;
logic [7:0] relu_99;
assign relu_99[7:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[21:15]}} :'d6) : '0;
logic [7:0] relu_100;
assign relu_100[7:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[21:15]}} :'d6) : '0;
logic [7:0] relu_101;
assign relu_101[7:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[21:15]}} :'d6) : '0;
logic [7:0] relu_102;
assign relu_102[7:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[21:15]}} :'d6) : '0;
logic [7:0] relu_103;
assign relu_103[7:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[21:15]}} :'d6) : '0;
logic [7:0] relu_104;
assign relu_104[7:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[21:15]}} :'d6) : '0;
logic [7:0] relu_105;
assign relu_105[7:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[21:15]}} :'d6) : '0;
logic [7:0] relu_106;
assign relu_106[7:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[21:15]}} :'d6) : '0;
logic [7:0] relu_107;
assign relu_107[7:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[21:15]}} :'d6) : '0;
logic [7:0] relu_108;
assign relu_108[7:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[21:15]}} :'d6) : '0;
logic [7:0] relu_109;
assign relu_109[7:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[21:15]}} :'d6) : '0;
logic [7:0] relu_110;
assign relu_110[7:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[21:15]}} :'d6) : '0;
logic [7:0] relu_111;
assign relu_111[7:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[21:15]}} :'d6) : '0;
logic [7:0] relu_112;
assign relu_112[7:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[21:15]}} :'d6) : '0;
logic [7:0] relu_113;
assign relu_113[7:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[21:15]}} :'d6) : '0;
logic [7:0] relu_114;
assign relu_114[7:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[21:15]}} :'d6) : '0;
logic [7:0] relu_115;
assign relu_115[7:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[21:15]}} :'d6) : '0;
logic [7:0] relu_116;
assign relu_116[7:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[21:15]}} :'d6) : '0;
logic [7:0] relu_117;
assign relu_117[7:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[21:15]}} :'d6) : '0;
logic [7:0] relu_118;
assign relu_118[7:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[21:15]}} :'d6) : '0;
logic [7:0] relu_119;
assign relu_119[7:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[21:15]}} :'d6) : '0;
logic [7:0] relu_120;
assign relu_120[7:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[21:15]}} :'d6) : '0;
logic [7:0] relu_121;
assign relu_121[7:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[21:15]}} :'d6) : '0;
logic [7:0] relu_122;
assign relu_122[7:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[21:15]}} :'d6) : '0;
logic [7:0] relu_123;
assign relu_123[7:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[21:15]}} :'d6) : '0;
logic [7:0] relu_124;
assign relu_124[7:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[21:15]}} :'d6) : '0;
logic [7:0] relu_125;
assign relu_125[7:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[21:15]}} :'d6) : '0;
logic [7:0] relu_126;
assign relu_126[7:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[21:15]}} :'d6) : '0;
logic [7:0] relu_127;
assign relu_127[7:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[21:15]}} :'d6) : '0;

assign output_act = {
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
