module conv9_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [2048-1:0] input_act,
    output logic [2048-1:0] output_act,
    output logic ready
);

logic [2048-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [15:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[15:0];
logic [15:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[31:16];
logic [15:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[47:32];
logic [15:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[63:48];
logic [15:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[79:64];
logic [15:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[95:80];
logic [15:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[111:96];
logic [15:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[127:112];
logic [15:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[143:128];
logic [15:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[159:144];
logic [15:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[175:160];
logic [15:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[191:176];
logic [15:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[207:192];
logic [15:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[223:208];
logic [15:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[239:224];
logic [15:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[255:240];
logic [15:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[271:256];
logic [15:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[287:272];
logic [15:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[303:288];
logic [15:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[319:304];
logic [15:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[335:320];
logic [15:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[351:336];
logic [15:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[367:352];
logic [15:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[383:368];
logic [15:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[399:384];
logic [15:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[415:400];
logic [15:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[431:416];
logic [15:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[447:432];
logic [15:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[463:448];
logic [15:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[479:464];
logic [15:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[495:480];
logic [15:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[511:496];
logic [15:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[527:512];
logic [15:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[543:528];
logic [15:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[559:544];
logic [15:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[575:560];
logic [15:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[591:576];
logic [15:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[607:592];
logic [15:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[623:608];
logic [15:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[639:624];
logic [15:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[655:640];
logic [15:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[671:656];
logic [15:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[687:672];
logic [15:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[703:688];
logic [15:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[719:704];
logic [15:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[735:720];
logic [15:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[751:736];
logic [15:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[767:752];
logic [15:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[783:768];
logic [15:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[799:784];
logic [15:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[815:800];
logic [15:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[831:816];
logic [15:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[847:832];
logic [15:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[863:848];
logic [15:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[879:864];
logic [15:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[895:880];
logic [15:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[911:896];
logic [15:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[927:912];
logic [15:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[943:928];
logic [15:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[959:944];
logic [15:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[975:960];
logic [15:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[991:976];
logic [15:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[1007:992];
logic [15:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[1023:1008];
logic [15:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[1039:1024];
logic [15:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[1055:1040];
logic [15:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[1071:1056];
logic [15:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[1087:1072];
logic [15:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[1103:1088];
logic [15:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[1119:1104];
logic [15:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[1135:1120];
logic [15:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[1151:1136];
logic [15:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[1167:1152];
logic [15:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[1183:1168];
logic [15:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[1199:1184];
logic [15:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[1215:1200];
logic [15:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[1231:1216];
logic [15:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[1247:1232];
logic [15:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[1263:1248];
logic [15:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[1279:1264];
logic [15:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[1295:1280];
logic [15:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[1311:1296];
logic [15:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[1327:1312];
logic [15:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[1343:1328];
logic [15:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[1359:1344];
logic [15:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[1375:1360];
logic [15:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[1391:1376];
logic [15:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[1407:1392];
logic [15:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[1423:1408];
logic [15:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[1439:1424];
logic [15:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[1455:1440];
logic [15:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[1471:1456];
logic [15:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[1487:1472];
logic [15:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[1503:1488];
logic [15:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[1519:1504];
logic [15:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[1535:1520];
logic [15:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[1551:1536];
logic [15:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[1567:1552];
logic [15:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[1583:1568];
logic [15:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[1599:1584];
logic [15:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[1615:1600];
logic [15:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[1631:1616];
logic [15:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[1647:1632];
logic [15:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[1663:1648];
logic [15:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[1679:1664];
logic [15:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[1695:1680];
logic [15:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[1711:1696];
logic [15:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[1727:1712];
logic [15:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[1743:1728];
logic [15:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[1759:1744];
logic [15:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[1775:1760];
logic [15:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[1791:1776];
logic [15:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[1807:1792];
logic [15:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[1823:1808];
logic [15:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[1839:1824];
logic [15:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[1855:1840];
logic [15:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[1871:1856];
logic [15:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[1887:1872];
logic [15:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[1903:1888];
logic [15:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[1919:1904];
logic [15:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[1935:1920];
logic [15:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[1951:1936];
logic [15:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[1967:1952];
logic [15:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[1983:1968];
logic [15:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[1999:1984];
logic [15:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[2015:2000];
logic [15:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[2031:2016];
logic [15:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[2047:2032];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 14'sd 5221) * $signed(input_fmap_0[15:0]) +
	( 12'sd 1889) * $signed(input_fmap_1[15:0]) +
	( 16'sd 16615) * $signed(input_fmap_2[15:0]) +
	( 10'sd 325) * $signed(input_fmap_3[15:0]) +
	( 14'sd 5426) * $signed(input_fmap_4[15:0]) +
	( 16'sd 32067) * $signed(input_fmap_5[15:0]) +
	( 12'sd 1465) * $signed(input_fmap_6[15:0]) +
	( 16'sd 17971) * $signed(input_fmap_7[15:0]) +
	( 14'sd 7263) * $signed(input_fmap_8[15:0]) +
	( 14'sd 6138) * $signed(input_fmap_9[15:0]) +
	( 15'sd 15754) * $signed(input_fmap_10[15:0]) +
	( 16'sd 26305) * $signed(input_fmap_11[15:0]) +
	( 16'sd 27660) * $signed(input_fmap_12[15:0]) +
	( 7'sd 62) * $signed(input_fmap_13[15:0]) +
	( 15'sd 16006) * $signed(input_fmap_14[15:0]) +
	( 16'sd 26604) * $signed(input_fmap_15[15:0]) +
	( 12'sd 1446) * $signed(input_fmap_16[15:0]) +
	( 14'sd 6408) * $signed(input_fmap_17[15:0]) +
	( 14'sd 4953) * $signed(input_fmap_18[15:0]) +
	( 16'sd 20766) * $signed(input_fmap_19[15:0]) +
	( 14'sd 4173) * $signed(input_fmap_20[15:0]) +
	( 12'sd 1388) * $signed(input_fmap_21[15:0]) +
	( 16'sd 19974) * $signed(input_fmap_22[15:0]) +
	( 13'sd 2185) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17278) * $signed(input_fmap_24[15:0]) +
	( 16'sd 17571) * $signed(input_fmap_25[15:0]) +
	( 15'sd 11287) * $signed(input_fmap_26[15:0]) +
	( 15'sd 14789) * $signed(input_fmap_27[15:0]) +
	( 16'sd 22769) * $signed(input_fmap_28[15:0]) +
	( 16'sd 26500) * $signed(input_fmap_29[15:0]) +
	( 15'sd 11559) * $signed(input_fmap_30[15:0]) +
	( 14'sd 6431) * $signed(input_fmap_31[15:0]) +
	( 16'sd 17893) * $signed(input_fmap_32[15:0]) +
	( 16'sd 23320) * $signed(input_fmap_33[15:0]) +
	( 15'sd 12039) * $signed(input_fmap_34[15:0]) +
	( 15'sd 8797) * $signed(input_fmap_35[15:0]) +
	( 16'sd 27712) * $signed(input_fmap_36[15:0]) +
	( 16'sd 23338) * $signed(input_fmap_37[15:0]) +
	( 16'sd 27534) * $signed(input_fmap_38[15:0]) +
	( 16'sd 29843) * $signed(input_fmap_39[15:0]) +
	( 16'sd 24160) * $signed(input_fmap_40[15:0]) +
	( 14'sd 7663) * $signed(input_fmap_41[15:0]) +
	( 12'sd 1982) * $signed(input_fmap_42[15:0]) +
	( 15'sd 16169) * $signed(input_fmap_43[15:0]) +
	( 13'sd 3651) * $signed(input_fmap_44[15:0]) +
	( 16'sd 32472) * $signed(input_fmap_45[15:0]) +
	( 15'sd 11672) * $signed(input_fmap_46[15:0]) +
	( 16'sd 25065) * $signed(input_fmap_47[15:0]) +
	( 15'sd 11870) * $signed(input_fmap_48[15:0]) +
	( 16'sd 22058) * $signed(input_fmap_49[15:0]) +
	( 16'sd 23174) * $signed(input_fmap_50[15:0]) +
	( 16'sd 26597) * $signed(input_fmap_51[15:0]) +
	( 14'sd 6011) * $signed(input_fmap_52[15:0]) +
	( 15'sd 9909) * $signed(input_fmap_53[15:0]) +
	( 16'sd 19477) * $signed(input_fmap_54[15:0]) +
	( 15'sd 11183) * $signed(input_fmap_55[15:0]) +
	( 15'sd 15412) * $signed(input_fmap_56[15:0]) +
	( 16'sd 25515) * $signed(input_fmap_57[15:0]) +
	( 16'sd 20109) * $signed(input_fmap_58[15:0]) +
	( 14'sd 7579) * $signed(input_fmap_59[15:0]) +
	( 15'sd 8339) * $signed(input_fmap_60[15:0]) +
	( 16'sd 30268) * $signed(input_fmap_61[15:0]) +
	( 16'sd 25657) * $signed(input_fmap_62[15:0]) +
	( 12'sd 1140) * $signed(input_fmap_63[15:0]) +
	( 15'sd 14598) * $signed(input_fmap_64[15:0]) +
	( 16'sd 31959) * $signed(input_fmap_65[15:0]) +
	( 15'sd 14577) * $signed(input_fmap_66[15:0]) +
	( 16'sd 31513) * $signed(input_fmap_67[15:0]) +
	( 12'sd 1249) * $signed(input_fmap_68[15:0]) +
	( 16'sd 24091) * $signed(input_fmap_69[15:0]) +
	( 15'sd 11899) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11154) * $signed(input_fmap_71[15:0]) +
	( 16'sd 26183) * $signed(input_fmap_72[15:0]) +
	( 15'sd 11365) * $signed(input_fmap_73[15:0]) +
	( 16'sd 24144) * $signed(input_fmap_74[15:0]) +
	( 13'sd 4022) * $signed(input_fmap_75[15:0]) +
	( 13'sd 3192) * $signed(input_fmap_76[15:0]) +
	( 15'sd 15112) * $signed(input_fmap_77[15:0]) +
	( 16'sd 19695) * $signed(input_fmap_78[15:0]) +
	( 12'sd 1289) * $signed(input_fmap_79[15:0]) +
	( 15'sd 13656) * $signed(input_fmap_80[15:0]) +
	( 16'sd 16500) * $signed(input_fmap_81[15:0]) +
	( 14'sd 7682) * $signed(input_fmap_82[15:0]) +
	( 16'sd 27034) * $signed(input_fmap_83[15:0]) +
	( 15'sd 8743) * $signed(input_fmap_84[15:0]) +
	( 16'sd 31208) * $signed(input_fmap_85[15:0]) +
	( 12'sd 1210) * $signed(input_fmap_86[15:0]) +
	( 16'sd 18961) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6281) * $signed(input_fmap_88[15:0]) +
	( 11'sd 796) * $signed(input_fmap_89[15:0]) +
	( 9'sd 167) * $signed(input_fmap_90[15:0]) +
	( 15'sd 8585) * $signed(input_fmap_91[15:0]) +
	( 16'sd 21752) * $signed(input_fmap_92[15:0]) +
	( 14'sd 6403) * $signed(input_fmap_93[15:0]) +
	( 15'sd 11387) * $signed(input_fmap_94[15:0]) +
	( 15'sd 15775) * $signed(input_fmap_95[15:0]) +
	( 16'sd 19415) * $signed(input_fmap_96[15:0]) +
	( 14'sd 7670) * $signed(input_fmap_97[15:0]) +
	( 15'sd 14457) * $signed(input_fmap_98[15:0]) +
	( 16'sd 16470) * $signed(input_fmap_99[15:0]) +
	( 13'sd 4085) * $signed(input_fmap_100[15:0]) +
	( 14'sd 7746) * $signed(input_fmap_101[15:0]) +
	( 15'sd 8234) * $signed(input_fmap_102[15:0]) +
	( 12'sd 1758) * $signed(input_fmap_103[15:0]) +
	( 16'sd 20629) * $signed(input_fmap_104[15:0]) +
	( 16'sd 24847) * $signed(input_fmap_105[15:0]) +
	( 15'sd 14189) * $signed(input_fmap_106[15:0]) +
	( 15'sd 13321) * $signed(input_fmap_107[15:0]) +
	( 11'sd 1006) * $signed(input_fmap_108[15:0]) +
	( 15'sd 11067) * $signed(input_fmap_109[15:0]) +
	( 16'sd 28448) * $signed(input_fmap_110[15:0]) +
	( 15'sd 15568) * $signed(input_fmap_111[15:0]) +
	( 16'sd 19508) * $signed(input_fmap_112[15:0]) +
	( 16'sd 17014) * $signed(input_fmap_113[15:0]) +
	( 12'sd 1471) * $signed(input_fmap_114[15:0]) +
	( 15'sd 10896) * $signed(input_fmap_115[15:0]) +
	( 15'sd 9594) * $signed(input_fmap_116[15:0]) +
	( 16'sd 24654) * $signed(input_fmap_117[15:0]) +
	( 16'sd 27482) * $signed(input_fmap_118[15:0]) +
	( 16'sd 18044) * $signed(input_fmap_119[15:0]) +
	( 10'sd 479) * $signed(input_fmap_120[15:0]) +
	( 16'sd 27133) * $signed(input_fmap_121[15:0]) +
	( 16'sd 18288) * $signed(input_fmap_122[15:0]) +
	( 16'sd 19174) * $signed(input_fmap_123[15:0]) +
	( 16'sd 31541) * $signed(input_fmap_124[15:0]) +
	( 14'sd 4571) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6745) * $signed(input_fmap_126[15:0]) +
	( 16'sd 31706) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 15'sd 16180) * $signed(input_fmap_0[15:0]) +
	( 16'sd 16524) * $signed(input_fmap_1[15:0]) +
	( 15'sd 9146) * $signed(input_fmap_2[15:0]) +
	( 16'sd 21406) * $signed(input_fmap_3[15:0]) +
	( 16'sd 32752) * $signed(input_fmap_4[15:0]) +
	( 16'sd 26144) * $signed(input_fmap_5[15:0]) +
	( 16'sd 29195) * $signed(input_fmap_6[15:0]) +
	( 16'sd 28129) * $signed(input_fmap_7[15:0]) +
	( 14'sd 8041) * $signed(input_fmap_8[15:0]) +
	( 15'sd 11438) * $signed(input_fmap_9[15:0]) +
	( 16'sd 24554) * $signed(input_fmap_10[15:0]) +
	( 11'sd 673) * $signed(input_fmap_11[15:0]) +
	( 13'sd 3677) * $signed(input_fmap_12[15:0]) +
	( 11'sd 604) * $signed(input_fmap_13[15:0]) +
	( 15'sd 13770) * $signed(input_fmap_14[15:0]) +
	( 16'sd 19636) * $signed(input_fmap_15[15:0]) +
	( 16'sd 21228) * $signed(input_fmap_16[15:0]) +
	( 14'sd 8042) * $signed(input_fmap_17[15:0]) +
	( 15'sd 9080) * $signed(input_fmap_18[15:0]) +
	( 15'sd 11933) * $signed(input_fmap_19[15:0]) +
	( 15'sd 10611) * $signed(input_fmap_20[15:0]) +
	( 13'sd 3106) * $signed(input_fmap_21[15:0]) +
	( 16'sd 19735) * $signed(input_fmap_22[15:0]) +
	( 16'sd 20727) * $signed(input_fmap_23[15:0]) +
	( 15'sd 11457) * $signed(input_fmap_24[15:0]) +
	( 16'sd 28832) * $signed(input_fmap_25[15:0]) +
	( 15'sd 14506) * $signed(input_fmap_26[15:0]) +
	( 16'sd 31786) * $signed(input_fmap_27[15:0]) +
	( 15'sd 12910) * $signed(input_fmap_28[15:0]) +
	( 13'sd 4059) * $signed(input_fmap_29[15:0]) +
	( 13'sd 2139) * $signed(input_fmap_30[15:0]) +
	( 16'sd 16784) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28573) * $signed(input_fmap_32[15:0]) +
	( 16'sd 29603) * $signed(input_fmap_33[15:0]) +
	( 13'sd 2598) * $signed(input_fmap_34[15:0]) +
	( 16'sd 32582) * $signed(input_fmap_35[15:0]) +
	( 15'sd 9579) * $signed(input_fmap_36[15:0]) +
	( 16'sd 27356) * $signed(input_fmap_37[15:0]) +
	( 15'sd 15543) * $signed(input_fmap_38[15:0]) +
	( 13'sd 4000) * $signed(input_fmap_39[15:0]) +
	( 16'sd 22663) * $signed(input_fmap_40[15:0]) +
	( 15'sd 10671) * $signed(input_fmap_41[15:0]) +
	( 16'sd 26654) * $signed(input_fmap_42[15:0]) +
	( 15'sd 11127) * $signed(input_fmap_43[15:0]) +
	( 14'sd 7089) * $signed(input_fmap_44[15:0]) +
	( 16'sd 32325) * $signed(input_fmap_45[15:0]) +
	( 15'sd 9023) * $signed(input_fmap_46[15:0]) +
	( 15'sd 10255) * $signed(input_fmap_47[15:0]) +
	( 16'sd 22698) * $signed(input_fmap_48[15:0]) +
	( 16'sd 31727) * $signed(input_fmap_49[15:0]) +
	( 16'sd 25126) * $signed(input_fmap_50[15:0]) +
	( 16'sd 31825) * $signed(input_fmap_51[15:0]) +
	( 16'sd 26826) * $signed(input_fmap_52[15:0]) +
	( 16'sd 18938) * $signed(input_fmap_53[15:0]) +
	( 16'sd 27592) * $signed(input_fmap_54[15:0]) +
	( 16'sd 18535) * $signed(input_fmap_55[15:0]) +
	( 16'sd 22439) * $signed(input_fmap_56[15:0]) +
	( 16'sd 32017) * $signed(input_fmap_57[15:0]) +
	( 16'sd 18249) * $signed(input_fmap_58[15:0]) +
	( 14'sd 5533) * $signed(input_fmap_59[15:0]) +
	( 15'sd 11009) * $signed(input_fmap_60[15:0]) +
	( 14'sd 7994) * $signed(input_fmap_61[15:0]) +
	( 11'sd 902) * $signed(input_fmap_62[15:0]) +
	( 13'sd 2618) * $signed(input_fmap_63[15:0]) +
	( 14'sd 4510) * $signed(input_fmap_64[15:0]) +
	( 16'sd 32690) * $signed(input_fmap_65[15:0]) +
	( 16'sd 30373) * $signed(input_fmap_66[15:0]) +
	( 15'sd 9524) * $signed(input_fmap_67[15:0]) +
	( 15'sd 13086) * $signed(input_fmap_68[15:0]) +
	( 14'sd 5445) * $signed(input_fmap_69[15:0]) +
	( 16'sd 24058) * $signed(input_fmap_70[15:0]) +
	( 13'sd 2905) * $signed(input_fmap_71[15:0]) +
	( 12'sd 1078) * $signed(input_fmap_72[15:0]) +
	( 13'sd 2396) * $signed(input_fmap_73[15:0]) +
	( 14'sd 6697) * $signed(input_fmap_74[15:0]) +
	( 13'sd 3128) * $signed(input_fmap_75[15:0]) +
	( 16'sd 27952) * $signed(input_fmap_76[15:0]) +
	( 16'sd 19956) * $signed(input_fmap_77[15:0]) +
	( 16'sd 23324) * $signed(input_fmap_78[15:0]) +
	( 16'sd 22319) * $signed(input_fmap_79[15:0]) +
	( 16'sd 22564) * $signed(input_fmap_80[15:0]) +
	( 15'sd 12848) * $signed(input_fmap_81[15:0]) +
	( 15'sd 8326) * $signed(input_fmap_82[15:0]) +
	( 16'sd 19859) * $signed(input_fmap_83[15:0]) +
	( 15'sd 14048) * $signed(input_fmap_84[15:0]) +
	( 15'sd 9534) * $signed(input_fmap_85[15:0]) +
	( 16'sd 27227) * $signed(input_fmap_86[15:0]) +
	( 16'sd 19437) * $signed(input_fmap_87[15:0]) +
	( 15'sd 10136) * $signed(input_fmap_88[15:0]) +
	( 14'sd 8117) * $signed(input_fmap_89[15:0]) +
	( 16'sd 23108) * $signed(input_fmap_90[15:0]) +
	( 16'sd 18457) * $signed(input_fmap_91[15:0]) +
	( 15'sd 15718) * $signed(input_fmap_92[15:0]) +
	( 16'sd 31320) * $signed(input_fmap_93[15:0]) +
	( 9'sd 157) * $signed(input_fmap_94[15:0]) +
	( 16'sd 26936) * $signed(input_fmap_95[15:0]) +
	( 14'sd 7202) * $signed(input_fmap_96[15:0]) +
	( 16'sd 28520) * $signed(input_fmap_97[15:0]) +
	( 15'sd 14538) * $signed(input_fmap_98[15:0]) +
	( 16'sd 26426) * $signed(input_fmap_99[15:0]) +
	( 16'sd 27392) * $signed(input_fmap_100[15:0]) +
	( 16'sd 20890) * $signed(input_fmap_101[15:0]) +
	( 16'sd 26105) * $signed(input_fmap_102[15:0]) +
	( 15'sd 14672) * $signed(input_fmap_103[15:0]) +
	( 16'sd 26488) * $signed(input_fmap_104[15:0]) +
	( 14'sd 5812) * $signed(input_fmap_105[15:0]) +
	( 16'sd 28699) * $signed(input_fmap_106[15:0]) +
	( 14'sd 5806) * $signed(input_fmap_107[15:0]) +
	( 15'sd 10669) * $signed(input_fmap_108[15:0]) +
	( 16'sd 25147) * $signed(input_fmap_109[15:0]) +
	( 16'sd 24597) * $signed(input_fmap_110[15:0]) +
	( 16'sd 32690) * $signed(input_fmap_111[15:0]) +
	( 16'sd 28419) * $signed(input_fmap_112[15:0]) +
	( 16'sd 25233) * $signed(input_fmap_113[15:0]) +
	( 14'sd 6653) * $signed(input_fmap_114[15:0]) +
	( 16'sd 26230) * $signed(input_fmap_115[15:0]) +
	( 13'sd 2759) * $signed(input_fmap_116[15:0]) +
	( 13'sd 2168) * $signed(input_fmap_117[15:0]) +
	( 14'sd 5458) * $signed(input_fmap_118[15:0]) +
	( 13'sd 2141) * $signed(input_fmap_119[15:0]) +
	( 15'sd 14466) * $signed(input_fmap_120[15:0]) +
	( 14'sd 7109) * $signed(input_fmap_121[15:0]) +
	( 16'sd 32715) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21082) * $signed(input_fmap_123[15:0]) +
	( 12'sd 1450) * $signed(input_fmap_124[15:0]) +
	( 14'sd 7696) * $signed(input_fmap_125[15:0]) +
	( 16'sd 31390) * $signed(input_fmap_126[15:0]) +
	( 15'sd 9721) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 16'sd 24132) * $signed(input_fmap_0[15:0]) +
	( 13'sd 2974) * $signed(input_fmap_1[15:0]) +
	( 16'sd 25734) * $signed(input_fmap_2[15:0]) +
	( 15'sd 11953) * $signed(input_fmap_3[15:0]) +
	( 13'sd 2628) * $signed(input_fmap_4[15:0]) +
	( 14'sd 4687) * $signed(input_fmap_5[15:0]) +
	( 16'sd 21341) * $signed(input_fmap_6[15:0]) +
	( 14'sd 6364) * $signed(input_fmap_7[15:0]) +
	( 16'sd 30658) * $signed(input_fmap_8[15:0]) +
	( 16'sd 20776) * $signed(input_fmap_9[15:0]) +
	( 16'sd 24674) * $signed(input_fmap_10[15:0]) +
	( 14'sd 7747) * $signed(input_fmap_11[15:0]) +
	( 16'sd 24928) * $signed(input_fmap_12[15:0]) +
	( 16'sd 21917) * $signed(input_fmap_13[15:0]) +
	( 16'sd 23777) * $signed(input_fmap_14[15:0]) +
	( 16'sd 29209) * $signed(input_fmap_15[15:0]) +
	( 15'sd 14316) * $signed(input_fmap_16[15:0]) +
	( 16'sd 31493) * $signed(input_fmap_17[15:0]) +
	( 16'sd 22841) * $signed(input_fmap_18[15:0]) +
	( 14'sd 5035) * $signed(input_fmap_19[15:0]) +
	( 16'sd 22657) * $signed(input_fmap_20[15:0]) +
	( 16'sd 23180) * $signed(input_fmap_21[15:0]) +
	( 16'sd 26789) * $signed(input_fmap_22[15:0]) +
	( 15'sd 15329) * $signed(input_fmap_23[15:0]) +
	( 13'sd 3033) * $signed(input_fmap_24[15:0]) +
	( 16'sd 18903) * $signed(input_fmap_25[15:0]) +
	( 13'sd 3029) * $signed(input_fmap_26[15:0]) +
	( 16'sd 19343) * $signed(input_fmap_27[15:0]) +
	( 16'sd 28522) * $signed(input_fmap_28[15:0]) +
	( 16'sd 25311) * $signed(input_fmap_29[15:0]) +
	( 16'sd 16503) * $signed(input_fmap_30[15:0]) +
	( 16'sd 20219) * $signed(input_fmap_31[15:0]) +
	( 15'sd 10265) * $signed(input_fmap_32[15:0]) +
	( 16'sd 24220) * $signed(input_fmap_33[15:0]) +
	( 15'sd 10547) * $signed(input_fmap_34[15:0]) +
	( 14'sd 4423) * $signed(input_fmap_35[15:0]) +
	( 16'sd 17000) * $signed(input_fmap_36[15:0]) +
	( 16'sd 25114) * $signed(input_fmap_37[15:0]) +
	( 13'sd 2067) * $signed(input_fmap_38[15:0]) +
	( 15'sd 10955) * $signed(input_fmap_39[15:0]) +
	( 14'sd 4375) * $signed(input_fmap_40[15:0]) +
	( 13'sd 2495) * $signed(input_fmap_41[15:0]) +
	( 12'sd 1355) * $signed(input_fmap_42[15:0]) +
	( 15'sd 9537) * $signed(input_fmap_43[15:0]) +
	( 16'sd 19968) * $signed(input_fmap_44[15:0]) +
	( 13'sd 3632) * $signed(input_fmap_45[15:0]) +
	( 16'sd 25599) * $signed(input_fmap_46[15:0]) +
	( 14'sd 5343) * $signed(input_fmap_47[15:0]) +
	( 16'sd 31393) * $signed(input_fmap_48[15:0]) +
	( 15'sd 9651) * $signed(input_fmap_49[15:0]) +
	( 12'sd 1788) * $signed(input_fmap_50[15:0]) +
	( 15'sd 11116) * $signed(input_fmap_51[15:0]) +
	( 16'sd 20217) * $signed(input_fmap_52[15:0]) +
	( 14'sd 6513) * $signed(input_fmap_53[15:0]) +
	( 15'sd 13394) * $signed(input_fmap_54[15:0]) +
	( 13'sd 3543) * $signed(input_fmap_55[15:0]) +
	( 15'sd 15709) * $signed(input_fmap_56[15:0]) +
	( 15'sd 13995) * $signed(input_fmap_57[15:0]) +
	( 15'sd 12734) * $signed(input_fmap_58[15:0]) +
	( 16'sd 23987) * $signed(input_fmap_59[15:0]) +
	( 16'sd 26109) * $signed(input_fmap_60[15:0]) +
	( 14'sd 5102) * $signed(input_fmap_61[15:0]) +
	( 14'sd 8032) * $signed(input_fmap_62[15:0]) +
	( 16'sd 22696) * $signed(input_fmap_63[15:0]) +
	( 14'sd 7948) * $signed(input_fmap_64[15:0]) +
	( 16'sd 22001) * $signed(input_fmap_65[15:0]) +
	( 16'sd 27322) * $signed(input_fmap_66[15:0]) +
	( 16'sd 21302) * $signed(input_fmap_67[15:0]) +
	( 13'sd 3404) * $signed(input_fmap_68[15:0]) +
	( 16'sd 32495) * $signed(input_fmap_69[15:0]) +
	( 15'sd 9104) * $signed(input_fmap_70[15:0]) +
	( 13'sd 3523) * $signed(input_fmap_71[15:0]) +
	( 16'sd 28400) * $signed(input_fmap_72[15:0]) +
	( 15'sd 14947) * $signed(input_fmap_73[15:0]) +
	( 16'sd 30281) * $signed(input_fmap_74[15:0]) +
	( 16'sd 30943) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19179) * $signed(input_fmap_76[15:0]) +
	( 16'sd 30535) * $signed(input_fmap_77[15:0]) +
	( 14'sd 6593) * $signed(input_fmap_78[15:0]) +
	( 15'sd 15543) * $signed(input_fmap_79[15:0]) +
	( 16'sd 17273) * $signed(input_fmap_80[15:0]) +
	( 16'sd 27037) * $signed(input_fmap_81[15:0]) +
	( 16'sd 22191) * $signed(input_fmap_82[15:0]) +
	( 15'sd 13866) * $signed(input_fmap_83[15:0]) +
	( 14'sd 6686) * $signed(input_fmap_84[15:0]) +
	( 16'sd 18126) * $signed(input_fmap_85[15:0]) +
	( 16'sd 16530) * $signed(input_fmap_86[15:0]) +
	( 16'sd 25720) * $signed(input_fmap_87[15:0]) +
	( 14'sd 5203) * $signed(input_fmap_88[15:0]) +
	( 16'sd 23633) * $signed(input_fmap_89[15:0]) +
	( 15'sd 12377) * $signed(input_fmap_90[15:0]) +
	( 14'sd 7705) * $signed(input_fmap_91[15:0]) +
	( 16'sd 30224) * $signed(input_fmap_92[15:0]) +
	( 15'sd 12563) * $signed(input_fmap_93[15:0]) +
	( 16'sd 24013) * $signed(input_fmap_94[15:0]) +
	( 14'sd 7022) * $signed(input_fmap_95[15:0]) +
	( 16'sd 29074) * $signed(input_fmap_96[15:0]) +
	( 14'sd 7162) * $signed(input_fmap_97[15:0]) +
	( 16'sd 18061) * $signed(input_fmap_98[15:0]) +
	( 15'sd 15159) * $signed(input_fmap_99[15:0]) +
	( 16'sd 21056) * $signed(input_fmap_100[15:0]) +
	( 14'sd 5190) * $signed(input_fmap_101[15:0]) +
	( 16'sd 32721) * $signed(input_fmap_102[15:0]) +
	( 14'sd 5695) * $signed(input_fmap_103[15:0]) +
	( 16'sd 27951) * $signed(input_fmap_104[15:0]) +
	( 16'sd 27466) * $signed(input_fmap_105[15:0]) +
	( 16'sd 27432) * $signed(input_fmap_106[15:0]) +
	( 14'sd 7851) * $signed(input_fmap_107[15:0]) +
	( 15'sd 14385) * $signed(input_fmap_108[15:0]) +
	( 16'sd 22774) * $signed(input_fmap_109[15:0]) +
	( 16'sd 31965) * $signed(input_fmap_110[15:0]) +
	( 14'sd 6755) * $signed(input_fmap_111[15:0]) +
	( 16'sd 27783) * $signed(input_fmap_112[15:0]) +
	( 13'sd 3501) * $signed(input_fmap_113[15:0]) +
	( 16'sd 23176) * $signed(input_fmap_114[15:0]) +
	( 16'sd 29973) * $signed(input_fmap_115[15:0]) +
	( 15'sd 9881) * $signed(input_fmap_116[15:0]) +
	( 15'sd 14681) * $signed(input_fmap_117[15:0]) +
	( 16'sd 24209) * $signed(input_fmap_118[15:0]) +
	( 16'sd 18509) * $signed(input_fmap_119[15:0]) +
	( 15'sd 8700) * $signed(input_fmap_120[15:0]) +
	( 16'sd 30290) * $signed(input_fmap_121[15:0]) +
	( 13'sd 2419) * $signed(input_fmap_122[15:0]) +
	( 16'sd 17040) * $signed(input_fmap_123[15:0]) +
	( 11'sd 776) * $signed(input_fmap_124[15:0]) +
	( 15'sd 15209) * $signed(input_fmap_125[15:0]) +
	( 15'sd 8672) * $signed(input_fmap_126[15:0]) +
	( 15'sd 9632) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 15'sd 16302) * $signed(input_fmap_0[15:0]) +
	( 15'sd 10556) * $signed(input_fmap_1[15:0]) +
	( 16'sd 28928) * $signed(input_fmap_2[15:0]) +
	( 7'sd 36) * $signed(input_fmap_3[15:0]) +
	( 15'sd 14032) * $signed(input_fmap_4[15:0]) +
	( 16'sd 25057) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2761) * $signed(input_fmap_6[15:0]) +
	( 15'sd 12352) * $signed(input_fmap_7[15:0]) +
	( 16'sd 21050) * $signed(input_fmap_8[15:0]) +
	( 16'sd 21044) * $signed(input_fmap_9[15:0]) +
	( 16'sd 27437) * $signed(input_fmap_10[15:0]) +
	( 16'sd 20058) * $signed(input_fmap_11[15:0]) +
	( 16'sd 31504) * $signed(input_fmap_12[15:0]) +
	( 15'sd 9779) * $signed(input_fmap_13[15:0]) +
	( 16'sd 32343) * $signed(input_fmap_14[15:0]) +
	( 14'sd 8008) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10947) * $signed(input_fmap_16[15:0]) +
	( 15'sd 14295) * $signed(input_fmap_17[15:0]) +
	( 13'sd 3731) * $signed(input_fmap_18[15:0]) +
	( 15'sd 11242) * $signed(input_fmap_19[15:0]) +
	( 14'sd 4608) * $signed(input_fmap_20[15:0]) +
	( 15'sd 13927) * $signed(input_fmap_21[15:0]) +
	( 16'sd 32361) * $signed(input_fmap_22[15:0]) +
	( 14'sd 6095) * $signed(input_fmap_23[15:0]) +
	( 15'sd 12885) * $signed(input_fmap_24[15:0]) +
	( 16'sd 19551) * $signed(input_fmap_25[15:0]) +
	( 16'sd 21006) * $signed(input_fmap_26[15:0]) +
	( 13'sd 3424) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24527) * $signed(input_fmap_28[15:0]) +
	( 16'sd 19642) * $signed(input_fmap_29[15:0]) +
	( 15'sd 10894) * $signed(input_fmap_30[15:0]) +
	( 15'sd 11775) * $signed(input_fmap_31[15:0]) +
	( 15'sd 8478) * $signed(input_fmap_32[15:0]) +
	( 16'sd 24637) * $signed(input_fmap_33[15:0]) +
	( 16'sd 20969) * $signed(input_fmap_34[15:0]) +
	( 16'sd 28710) * $signed(input_fmap_35[15:0]) +
	( 15'sd 9667) * $signed(input_fmap_36[15:0]) +
	( 15'sd 10266) * $signed(input_fmap_37[15:0]) +
	( 12'sd 1157) * $signed(input_fmap_38[15:0]) +
	( 16'sd 23976) * $signed(input_fmap_39[15:0]) +
	( 10'sd 370) * $signed(input_fmap_40[15:0]) +
	( 16'sd 31268) * $signed(input_fmap_41[15:0]) +
	( 13'sd 3291) * $signed(input_fmap_42[15:0]) +
	( 16'sd 19145) * $signed(input_fmap_43[15:0]) +
	( 16'sd 26135) * $signed(input_fmap_44[15:0]) +
	( 15'sd 11073) * $signed(input_fmap_45[15:0]) +
	( 15'sd 14917) * $signed(input_fmap_46[15:0]) +
	( 16'sd 21491) * $signed(input_fmap_47[15:0]) +
	( 13'sd 4030) * $signed(input_fmap_48[15:0]) +
	( 15'sd 14701) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22464) * $signed(input_fmap_50[15:0]) +
	( 15'sd 8208) * $signed(input_fmap_51[15:0]) +
	( 15'sd 12107) * $signed(input_fmap_52[15:0]) +
	( 16'sd 25549) * $signed(input_fmap_53[15:0]) +
	( 16'sd 21803) * $signed(input_fmap_54[15:0]) +
	( 10'sd 327) * $signed(input_fmap_55[15:0]) +
	( 16'sd 23733) * $signed(input_fmap_56[15:0]) +
	( 16'sd 20749) * $signed(input_fmap_57[15:0]) +
	( 12'sd 1286) * $signed(input_fmap_58[15:0]) +
	( 16'sd 18566) * $signed(input_fmap_59[15:0]) +
	( 15'sd 15150) * $signed(input_fmap_60[15:0]) +
	( 13'sd 2293) * $signed(input_fmap_61[15:0]) +
	( 16'sd 17518) * $signed(input_fmap_62[15:0]) +
	( 16'sd 21930) * $signed(input_fmap_63[15:0]) +
	( 16'sd 17495) * $signed(input_fmap_64[15:0]) +
	( 16'sd 27942) * $signed(input_fmap_65[15:0]) +
	( 16'sd 31250) * $signed(input_fmap_66[15:0]) +
	( 16'sd 25844) * $signed(input_fmap_67[15:0]) +
	( 14'sd 6089) * $signed(input_fmap_68[15:0]) +
	( 12'sd 1418) * $signed(input_fmap_69[15:0]) +
	( 16'sd 22112) * $signed(input_fmap_70[15:0]) +
	( 16'sd 19020) * $signed(input_fmap_71[15:0]) +
	( 16'sd 21012) * $signed(input_fmap_72[15:0]) +
	( 16'sd 31220) * $signed(input_fmap_73[15:0]) +
	( 16'sd 27630) * $signed(input_fmap_74[15:0]) +
	( 12'sd 1307) * $signed(input_fmap_75[15:0]) +
	( 14'sd 6201) * $signed(input_fmap_76[15:0]) +
	( 15'sd 9132) * $signed(input_fmap_77[15:0]) +
	( 16'sd 23505) * $signed(input_fmap_78[15:0]) +
	( 16'sd 22017) * $signed(input_fmap_79[15:0]) +
	( 15'sd 12223) * $signed(input_fmap_80[15:0]) +
	( 16'sd 19588) * $signed(input_fmap_81[15:0]) +
	( 12'sd 1156) * $signed(input_fmap_82[15:0]) +
	( 16'sd 26220) * $signed(input_fmap_83[15:0]) +
	( 16'sd 16573) * $signed(input_fmap_84[15:0]) +
	( 16'sd 31237) * $signed(input_fmap_85[15:0]) +
	( 16'sd 18766) * $signed(input_fmap_86[15:0]) +
	( 16'sd 27655) * $signed(input_fmap_87[15:0]) +
	( 16'sd 31282) * $signed(input_fmap_88[15:0]) +
	( 12'sd 1139) * $signed(input_fmap_89[15:0]) +
	( 15'sd 11212) * $signed(input_fmap_90[15:0]) +
	( 16'sd 28120) * $signed(input_fmap_91[15:0]) +
	( 16'sd 27848) * $signed(input_fmap_92[15:0]) +
	( 15'sd 8384) * $signed(input_fmap_93[15:0]) +
	( 13'sd 2386) * $signed(input_fmap_94[15:0]) +
	( 11'sd 517) * $signed(input_fmap_95[15:0]) +
	( 16'sd 29382) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27047) * $signed(input_fmap_97[15:0]) +
	( 16'sd 30139) * $signed(input_fmap_98[15:0]) +
	( 15'sd 10860) * $signed(input_fmap_99[15:0]) +
	( 16'sd 18574) * $signed(input_fmap_100[15:0]) +
	( 16'sd 17869) * $signed(input_fmap_101[15:0]) +
	( 16'sd 19205) * $signed(input_fmap_102[15:0]) +
	( 16'sd 20041) * $signed(input_fmap_103[15:0]) +
	( 15'sd 13662) * $signed(input_fmap_104[15:0]) +
	( 14'sd 6571) * $signed(input_fmap_105[15:0]) +
	( 16'sd 28655) * $signed(input_fmap_106[15:0]) +
	( 16'sd 17881) * $signed(input_fmap_107[15:0]) +
	( 16'sd 25814) * $signed(input_fmap_108[15:0]) +
	( 14'sd 7631) * $signed(input_fmap_109[15:0]) +
	( 15'sd 10899) * $signed(input_fmap_110[15:0]) +
	( 12'sd 1628) * $signed(input_fmap_111[15:0]) +
	( 16'sd 30377) * $signed(input_fmap_112[15:0]) +
	( 16'sd 27513) * $signed(input_fmap_113[15:0]) +
	( 15'sd 10951) * $signed(input_fmap_114[15:0]) +
	( 16'sd 20575) * $signed(input_fmap_115[15:0]) +
	( 11'sd 607) * $signed(input_fmap_116[15:0]) +
	( 16'sd 18540) * $signed(input_fmap_117[15:0]) +
	( 13'sd 2538) * $signed(input_fmap_118[15:0]) +
	( 15'sd 15383) * $signed(input_fmap_119[15:0]) +
	( 16'sd 23227) * $signed(input_fmap_120[15:0]) +
	( 16'sd 28222) * $signed(input_fmap_121[15:0]) +
	( 16'sd 30995) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21779) * $signed(input_fmap_123[15:0]) +
	( 15'sd 13149) * $signed(input_fmap_124[15:0]) +
	( 16'sd 22112) * $signed(input_fmap_125[15:0]) +
	( 15'sd 9629) * $signed(input_fmap_126[15:0]) +
	( 14'sd 6561) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 16'sd 19134) * $signed(input_fmap_0[15:0]) +
	( 15'sd 16165) * $signed(input_fmap_1[15:0]) +
	( 16'sd 19094) * $signed(input_fmap_2[15:0]) +
	( 16'sd 20389) * $signed(input_fmap_3[15:0]) +
	( 16'sd 28787) * $signed(input_fmap_4[15:0]) +
	( 16'sd 28868) * $signed(input_fmap_5[15:0]) +
	( 15'sd 9306) * $signed(input_fmap_6[15:0]) +
	( 16'sd 17421) * $signed(input_fmap_7[15:0]) +
	( 16'sd 25611) * $signed(input_fmap_8[15:0]) +
	( 16'sd 23577) * $signed(input_fmap_9[15:0]) +
	( 16'sd 22136) * $signed(input_fmap_10[15:0]) +
	( 16'sd 25066) * $signed(input_fmap_11[15:0]) +
	( 16'sd 22322) * $signed(input_fmap_12[15:0]) +
	( 16'sd 18808) * $signed(input_fmap_13[15:0]) +
	( 16'sd 22970) * $signed(input_fmap_14[15:0]) +
	( 15'sd 9879) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10235) * $signed(input_fmap_16[15:0]) +
	( 15'sd 14962) * $signed(input_fmap_17[15:0]) +
	( 16'sd 25384) * $signed(input_fmap_18[15:0]) +
	( 12'sd 1345) * $signed(input_fmap_19[15:0]) +
	( 12'sd 1379) * $signed(input_fmap_20[15:0]) +
	( 13'sd 3837) * $signed(input_fmap_21[15:0]) +
	( 16'sd 21927) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28946) * $signed(input_fmap_23[15:0]) +
	( 11'sd 624) * $signed(input_fmap_24[15:0]) +
	( 15'sd 15269) * $signed(input_fmap_25[15:0]) +
	( 16'sd 28695) * $signed(input_fmap_26[15:0]) +
	( 15'sd 10777) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24271) * $signed(input_fmap_28[15:0]) +
	( 14'sd 4127) * $signed(input_fmap_29[15:0]) +
	( 14'sd 5195) * $signed(input_fmap_30[15:0]) +
	( 12'sd 1728) * $signed(input_fmap_31[15:0]) +
	( 16'sd 24695) * $signed(input_fmap_32[15:0]) +
	( 14'sd 7732) * $signed(input_fmap_33[15:0]) +
	( 12'sd 1305) * $signed(input_fmap_34[15:0]) +
	( 16'sd 23610) * $signed(input_fmap_35[15:0]) +
	( 15'sd 9888) * $signed(input_fmap_36[15:0]) +
	( 16'sd 16567) * $signed(input_fmap_37[15:0]) +
	( 16'sd 29168) * $signed(input_fmap_38[15:0]) +
	( 16'sd 16717) * $signed(input_fmap_39[15:0]) +
	( 15'sd 16118) * $signed(input_fmap_40[15:0]) +
	( 16'sd 20829) * $signed(input_fmap_41[15:0]) +
	( 16'sd 29945) * $signed(input_fmap_42[15:0]) +
	( 15'sd 11915) * $signed(input_fmap_43[15:0]) +
	( 16'sd 20849) * $signed(input_fmap_44[15:0]) +
	( 14'sd 7448) * $signed(input_fmap_45[15:0]) +
	( 16'sd 23148) * $signed(input_fmap_46[15:0]) +
	( 16'sd 17377) * $signed(input_fmap_47[15:0]) +
	( 15'sd 10706) * $signed(input_fmap_48[15:0]) +
	( 14'sd 5581) * $signed(input_fmap_49[15:0]) +
	( 14'sd 6522) * $signed(input_fmap_50[15:0]) +
	( 14'sd 5502) * $signed(input_fmap_51[15:0]) +
	( 16'sd 28956) * $signed(input_fmap_52[15:0]) +
	( 16'sd 23675) * $signed(input_fmap_53[15:0]) +
	( 16'sd 16910) * $signed(input_fmap_54[15:0]) +
	( 16'sd 25731) * $signed(input_fmap_55[15:0]) +
	( 16'sd 26218) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17298) * $signed(input_fmap_57[15:0]) +
	( 15'sd 11863) * $signed(input_fmap_58[15:0]) +
	( 16'sd 21528) * $signed(input_fmap_59[15:0]) +
	( 16'sd 30507) * $signed(input_fmap_60[15:0]) +
	( 15'sd 9827) * $signed(input_fmap_61[15:0]) +
	( 16'sd 16679) * $signed(input_fmap_62[15:0]) +
	( 14'sd 4166) * $signed(input_fmap_63[15:0]) +
	( 15'sd 10422) * $signed(input_fmap_64[15:0]) +
	( 15'sd 12076) * $signed(input_fmap_65[15:0]) +
	( 14'sd 6929) * $signed(input_fmap_66[15:0]) +
	( 16'sd 23822) * $signed(input_fmap_67[15:0]) +
	( 16'sd 18396) * $signed(input_fmap_68[15:0]) +
	( 16'sd 24864) * $signed(input_fmap_69[15:0]) +
	( 15'sd 13972) * $signed(input_fmap_70[15:0]) +
	( 15'sd 13669) * $signed(input_fmap_71[15:0]) +
	( 12'sd 1634) * $signed(input_fmap_72[15:0]) +
	( 7'sd 45) * $signed(input_fmap_73[15:0]) +
	( 13'sd 3120) * $signed(input_fmap_74[15:0]) +
	( 15'sd 10689) * $signed(input_fmap_75[15:0]) +
	( 15'sd 12410) * $signed(input_fmap_76[15:0]) +
	( 13'sd 2064) * $signed(input_fmap_77[15:0]) +
	( 15'sd 9191) * $signed(input_fmap_78[15:0]) +
	( 14'sd 4732) * $signed(input_fmap_79[15:0]) +
	( 16'sd 17579) * $signed(input_fmap_80[15:0]) +
	( 15'sd 12861) * $signed(input_fmap_81[15:0]) +
	( 16'sd 21723) * $signed(input_fmap_82[15:0]) +
	( 15'sd 14433) * $signed(input_fmap_83[15:0]) +
	( 12'sd 1346) * $signed(input_fmap_84[15:0]) +
	( 16'sd 19825) * $signed(input_fmap_85[15:0]) +
	( 16'sd 19684) * $signed(input_fmap_86[15:0]) +
	( 12'sd 1563) * $signed(input_fmap_87[15:0]) +
	( 16'sd 30185) * $signed(input_fmap_88[15:0]) +
	( 14'sd 4489) * $signed(input_fmap_89[15:0]) +
	( 16'sd 23833) * $signed(input_fmap_90[15:0]) +
	( 16'sd 23756) * $signed(input_fmap_91[15:0]) +
	( 16'sd 30615) * $signed(input_fmap_92[15:0]) +
	( 15'sd 14475) * $signed(input_fmap_93[15:0]) +
	( 16'sd 16510) * $signed(input_fmap_94[15:0]) +
	( 16'sd 29298) * $signed(input_fmap_95[15:0]) +
	( 15'sd 11332) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27364) * $signed(input_fmap_97[15:0]) +
	( 15'sd 10760) * $signed(input_fmap_98[15:0]) +
	( 15'sd 10769) * $signed(input_fmap_99[15:0]) +
	( 15'sd 15869) * $signed(input_fmap_100[15:0]) +
	( 16'sd 24125) * $signed(input_fmap_101[15:0]) +
	( 16'sd 18650) * $signed(input_fmap_102[15:0]) +
	( 16'sd 18038) * $signed(input_fmap_103[15:0]) +
	( 16'sd 31830) * $signed(input_fmap_104[15:0]) +
	( 16'sd 21342) * $signed(input_fmap_105[15:0]) +
	( 14'sd 7421) * $signed(input_fmap_106[15:0]) +
	( 13'sd 3287) * $signed(input_fmap_107[15:0]) +
	( 15'sd 11808) * $signed(input_fmap_108[15:0]) +
	( 16'sd 17034) * $signed(input_fmap_109[15:0]) +
	( 16'sd 21861) * $signed(input_fmap_110[15:0]) +
	( 16'sd 23926) * $signed(input_fmap_111[15:0]) +
	( 15'sd 13886) * $signed(input_fmap_112[15:0]) +
	( 15'sd 14877) * $signed(input_fmap_113[15:0]) +
	( 16'sd 19413) * $signed(input_fmap_114[15:0]) +
	( 16'sd 31742) * $signed(input_fmap_115[15:0]) +
	( 14'sd 5809) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27081) * $signed(input_fmap_117[15:0]) +
	( 16'sd 32492) * $signed(input_fmap_118[15:0]) +
	( 15'sd 8750) * $signed(input_fmap_119[15:0]) +
	( 15'sd 14756) * $signed(input_fmap_120[15:0]) +
	( 16'sd 24041) * $signed(input_fmap_121[15:0]) +
	( 15'sd 13321) * $signed(input_fmap_122[15:0]) +
	( 11'sd 635) * $signed(input_fmap_123[15:0]) +
	( 14'sd 5785) * $signed(input_fmap_124[15:0]) +
	( 16'sd 23472) * $signed(input_fmap_125[15:0]) +
	( 15'sd 10023) * $signed(input_fmap_126[15:0]) +
	( 15'sd 11102) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 15'sd 10560) * $signed(input_fmap_0[15:0]) +
	( 16'sd 30565) * $signed(input_fmap_1[15:0]) +
	( 15'sd 12824) * $signed(input_fmap_2[15:0]) +
	( 16'sd 28033) * $signed(input_fmap_3[15:0]) +
	( 14'sd 5410) * $signed(input_fmap_4[15:0]) +
	( 16'sd 31941) * $signed(input_fmap_5[15:0]) +
	( 16'sd 18875) * $signed(input_fmap_6[15:0]) +
	( 16'sd 26353) * $signed(input_fmap_7[15:0]) +
	( 14'sd 6490) * $signed(input_fmap_8[15:0]) +
	( 14'sd 7132) * $signed(input_fmap_9[15:0]) +
	( 15'sd 12113) * $signed(input_fmap_10[15:0]) +
	( 16'sd 25943) * $signed(input_fmap_11[15:0]) +
	( 16'sd 19547) * $signed(input_fmap_12[15:0]) +
	( 15'sd 16225) * $signed(input_fmap_13[15:0]) +
	( 16'sd 32749) * $signed(input_fmap_14[15:0]) +
	( 15'sd 12069) * $signed(input_fmap_15[15:0]) +
	( 16'sd 20385) * $signed(input_fmap_16[15:0]) +
	( 16'sd 30530) * $signed(input_fmap_17[15:0]) +
	( 12'sd 1490) * $signed(input_fmap_18[15:0]) +
	( 16'sd 21149) * $signed(input_fmap_19[15:0]) +
	( 16'sd 17862) * $signed(input_fmap_20[15:0]) +
	( 16'sd 19442) * $signed(input_fmap_21[15:0]) +
	( 16'sd 25823) * $signed(input_fmap_22[15:0]) +
	( 16'sd 25912) * $signed(input_fmap_23[15:0]) +
	( 15'sd 16317) * $signed(input_fmap_24[15:0]) +
	( 16'sd 28936) * $signed(input_fmap_25[15:0]) +
	( 15'sd 8417) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9152) * $signed(input_fmap_27[15:0]) +
	( 16'sd 21868) * $signed(input_fmap_28[15:0]) +
	( 14'sd 6513) * $signed(input_fmap_29[15:0]) +
	( 15'sd 14186) * $signed(input_fmap_30[15:0]) +
	( 15'sd 10006) * $signed(input_fmap_31[15:0]) +
	( 16'sd 24493) * $signed(input_fmap_32[15:0]) +
	( 16'sd 17238) * $signed(input_fmap_33[15:0]) +
	( 16'sd 24765) * $signed(input_fmap_34[15:0]) +
	( 16'sd 21688) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11902) * $signed(input_fmap_36[15:0]) +
	( 15'sd 15463) * $signed(input_fmap_37[15:0]) +
	( 16'sd 31681) * $signed(input_fmap_38[15:0]) +
	( 16'sd 26805) * $signed(input_fmap_39[15:0]) +
	( 10'sd 361) * $signed(input_fmap_40[15:0]) +
	( 16'sd 25863) * $signed(input_fmap_41[15:0]) +
	( 16'sd 22170) * $signed(input_fmap_42[15:0]) +
	( 11'sd 739) * $signed(input_fmap_43[15:0]) +
	( 16'sd 25953) * $signed(input_fmap_44[15:0]) +
	( 16'sd 30822) * $signed(input_fmap_45[15:0]) +
	( 15'sd 9263) * $signed(input_fmap_46[15:0]) +
	( 16'sd 24135) * $signed(input_fmap_47[15:0]) +
	( 16'sd 32570) * $signed(input_fmap_48[15:0]) +
	( 16'sd 16408) * $signed(input_fmap_49[15:0]) +
	( 15'sd 13868) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15383) * $signed(input_fmap_51[15:0]) +
	( 16'sd 30041) * $signed(input_fmap_52[15:0]) +
	( 15'sd 8887) * $signed(input_fmap_53[15:0]) +
	( 16'sd 24543) * $signed(input_fmap_54[15:0]) +
	( 16'sd 26595) * $signed(input_fmap_55[15:0]) +
	( 16'sd 17536) * $signed(input_fmap_56[15:0]) +
	( 16'sd 18644) * $signed(input_fmap_57[15:0]) +
	( 15'sd 14019) * $signed(input_fmap_58[15:0]) +
	( 15'sd 10529) * $signed(input_fmap_59[15:0]) +
	( 15'sd 13316) * $signed(input_fmap_60[15:0]) +
	( 16'sd 18632) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3723) * $signed(input_fmap_62[15:0]) +
	( 14'sd 8128) * $signed(input_fmap_63[15:0]) +
	( 16'sd 27100) * $signed(input_fmap_64[15:0]) +
	( 16'sd 18072) * $signed(input_fmap_65[15:0]) +
	( 16'sd 17876) * $signed(input_fmap_66[15:0]) +
	( 14'sd 4170) * $signed(input_fmap_67[15:0]) +
	( 16'sd 29232) * $signed(input_fmap_68[15:0]) +
	( 15'sd 12899) * $signed(input_fmap_69[15:0]) +
	( 16'sd 30856) * $signed(input_fmap_70[15:0]) +
	( 16'sd 30291) * $signed(input_fmap_71[15:0]) +
	( 15'sd 15982) * $signed(input_fmap_72[15:0]) +
	( 15'sd 9787) * $signed(input_fmap_73[15:0]) +
	( 16'sd 32545) * $signed(input_fmap_74[15:0]) +
	( 16'sd 29002) * $signed(input_fmap_75[15:0]) +
	( 16'sd 21683) * $signed(input_fmap_76[15:0]) +
	( 16'sd 23740) * $signed(input_fmap_77[15:0]) +
	( 16'sd 25551) * $signed(input_fmap_78[15:0]) +
	( 16'sd 27877) * $signed(input_fmap_79[15:0]) +
	( 16'sd 19133) * $signed(input_fmap_80[15:0]) +
	( 16'sd 25664) * $signed(input_fmap_81[15:0]) +
	( 16'sd 26710) * $signed(input_fmap_82[15:0]) +
	( 15'sd 9230) * $signed(input_fmap_83[15:0]) +
	( 16'sd 17445) * $signed(input_fmap_84[15:0]) +
	( 15'sd 12548) * $signed(input_fmap_85[15:0]) +
	( 14'sd 7178) * $signed(input_fmap_86[15:0]) +
	( 16'sd 31451) * $signed(input_fmap_87[15:0]) +
	( 15'sd 14764) * $signed(input_fmap_88[15:0]) +
	( 14'sd 8163) * $signed(input_fmap_89[15:0]) +
	( 16'sd 24436) * $signed(input_fmap_90[15:0]) +
	( 16'sd 31416) * $signed(input_fmap_91[15:0]) +
	( 13'sd 3120) * $signed(input_fmap_92[15:0]) +
	( 15'sd 14645) * $signed(input_fmap_93[15:0]) +
	( 16'sd 28248) * $signed(input_fmap_94[15:0]) +
	( 16'sd 19280) * $signed(input_fmap_95[15:0]) +
	( 16'sd 25479) * $signed(input_fmap_96[15:0]) +
	( 16'sd 19155) * $signed(input_fmap_97[15:0]) +
	( 14'sd 5766) * $signed(input_fmap_98[15:0]) +
	( 12'sd 1380) * $signed(input_fmap_99[15:0]) +
	( 14'sd 7600) * $signed(input_fmap_100[15:0]) +
	( 13'sd 2129) * $signed(input_fmap_101[15:0]) +
	( 15'sd 13760) * $signed(input_fmap_102[15:0]) +
	( 12'sd 1344) * $signed(input_fmap_103[15:0]) +
	( 14'sd 6931) * $signed(input_fmap_104[15:0]) +
	( 15'sd 12760) * $signed(input_fmap_105[15:0]) +
	( 16'sd 30053) * $signed(input_fmap_106[15:0]) +
	( 16'sd 31661) * $signed(input_fmap_107[15:0]) +
	( 16'sd 21359) * $signed(input_fmap_108[15:0]) +
	( 16'sd 30438) * $signed(input_fmap_109[15:0]) +
	( 13'sd 2740) * $signed(input_fmap_110[15:0]) +
	( 16'sd 18223) * $signed(input_fmap_111[15:0]) +
	( 15'sd 9112) * $signed(input_fmap_112[15:0]) +
	( 16'sd 24001) * $signed(input_fmap_113[15:0]) +
	( 14'sd 4868) * $signed(input_fmap_114[15:0]) +
	( 14'sd 6525) * $signed(input_fmap_115[15:0]) +
	( 16'sd 19479) * $signed(input_fmap_116[15:0]) +
	( 15'sd 10483) * $signed(input_fmap_117[15:0]) +
	( 16'sd 31028) * $signed(input_fmap_118[15:0]) +
	( 13'sd 2606) * $signed(input_fmap_119[15:0]) +
	( 16'sd 25974) * $signed(input_fmap_120[15:0]) +
	( 14'sd 4860) * $signed(input_fmap_121[15:0]) +
	( 16'sd 26737) * $signed(input_fmap_122[15:0]) +
	( 14'sd 8014) * $signed(input_fmap_123[15:0]) +
	( 14'sd 5136) * $signed(input_fmap_124[15:0]) +
	( 14'sd 4682) * $signed(input_fmap_125[15:0]) +
	( 16'sd 17226) * $signed(input_fmap_126[15:0]) +
	( 16'sd 17715) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 15'sd 12180) * $signed(input_fmap_0[15:0]) +
	( 15'sd 12455) * $signed(input_fmap_1[15:0]) +
	( 10'sd 484) * $signed(input_fmap_2[15:0]) +
	( 10'sd 261) * $signed(input_fmap_3[15:0]) +
	( 15'sd 12221) * $signed(input_fmap_4[15:0]) +
	( 15'sd 12679) * $signed(input_fmap_5[15:0]) +
	( 16'sd 30422) * $signed(input_fmap_6[15:0]) +
	( 16'sd 25923) * $signed(input_fmap_7[15:0]) +
	( 15'sd 13343) * $signed(input_fmap_8[15:0]) +
	( 16'sd 27072) * $signed(input_fmap_9[15:0]) +
	( 13'sd 3977) * $signed(input_fmap_10[15:0]) +
	( 15'sd 12256) * $signed(input_fmap_11[15:0]) +
	( 15'sd 13600) * $signed(input_fmap_12[15:0]) +
	( 16'sd 27683) * $signed(input_fmap_13[15:0]) +
	( 15'sd 13221) * $signed(input_fmap_14[15:0]) +
	( 15'sd 9837) * $signed(input_fmap_15[15:0]) +
	( 16'sd 19114) * $signed(input_fmap_16[15:0]) +
	( 13'sd 2193) * $signed(input_fmap_17[15:0]) +
	( 16'sd 28195) * $signed(input_fmap_18[15:0]) +
	( 16'sd 17216) * $signed(input_fmap_19[15:0]) +
	( 15'sd 8320) * $signed(input_fmap_20[15:0]) +
	( 14'sd 5193) * $signed(input_fmap_21[15:0]) +
	( 16'sd 21676) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24907) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17673) * $signed(input_fmap_24[15:0]) +
	( 16'sd 28395) * $signed(input_fmap_25[15:0]) +
	( 15'sd 16326) * $signed(input_fmap_26[15:0]) +
	( 16'sd 23011) * $signed(input_fmap_27[15:0]) +
	( 16'sd 20677) * $signed(input_fmap_28[15:0]) +
	( 15'sd 10059) * $signed(input_fmap_29[15:0]) +
	( 15'sd 9277) * $signed(input_fmap_30[15:0]) +
	( 16'sd 20796) * $signed(input_fmap_31[15:0]) +
	( 14'sd 5334) * $signed(input_fmap_32[15:0]) +
	( 16'sd 16772) * $signed(input_fmap_33[15:0]) +
	( 16'sd 26136) * $signed(input_fmap_34[15:0]) +
	( 9'sd 131) * $signed(input_fmap_35[15:0]) +
	( 15'sd 12847) * $signed(input_fmap_36[15:0]) +
	( 16'sd 29865) * $signed(input_fmap_37[15:0]) +
	( 16'sd 31697) * $signed(input_fmap_38[15:0]) +
	( 16'sd 25298) * $signed(input_fmap_39[15:0]) +
	( 16'sd 27267) * $signed(input_fmap_40[15:0]) +
	( 15'sd 13492) * $signed(input_fmap_41[15:0]) +
	( 16'sd 20856) * $signed(input_fmap_42[15:0]) +
	( 15'sd 12593) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31864) * $signed(input_fmap_44[15:0]) +
	( 16'sd 29952) * $signed(input_fmap_45[15:0]) +
	( 15'sd 12909) * $signed(input_fmap_46[15:0]) +
	( 14'sd 5941) * $signed(input_fmap_47[15:0]) +
	( 14'sd 6326) * $signed(input_fmap_48[15:0]) +
	( 16'sd 27211) * $signed(input_fmap_49[15:0]) +
	( 16'sd 17037) * $signed(input_fmap_50[15:0]) +
	( 15'sd 16114) * $signed(input_fmap_51[15:0]) +
	( 16'sd 17863) * $signed(input_fmap_52[15:0]) +
	( 16'sd 23169) * $signed(input_fmap_53[15:0]) +
	( 16'sd 28533) * $signed(input_fmap_54[15:0]) +
	( 16'sd 25642) * $signed(input_fmap_55[15:0]) +
	( 16'sd 22288) * $signed(input_fmap_56[15:0]) +
	( 16'sd 29497) * $signed(input_fmap_57[15:0]) +
	( 16'sd 32020) * $signed(input_fmap_58[15:0]) +
	( 16'sd 18373) * $signed(input_fmap_59[15:0]) +
	( 15'sd 10117) * $signed(input_fmap_60[15:0]) +
	( 16'sd 17098) * $signed(input_fmap_61[15:0]) +
	( 16'sd 24014) * $signed(input_fmap_62[15:0]) +
	( 16'sd 28075) * $signed(input_fmap_63[15:0]) +
	( 16'sd 28101) * $signed(input_fmap_64[15:0]) +
	( 16'sd 21019) * $signed(input_fmap_65[15:0]) +
	( 16'sd 25162) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28591) * $signed(input_fmap_67[15:0]) +
	( 15'sd 10037) * $signed(input_fmap_68[15:0]) +
	( 15'sd 11390) * $signed(input_fmap_69[15:0]) +
	( 16'sd 19246) * $signed(input_fmap_70[15:0]) +
	( 16'sd 32470) * $signed(input_fmap_71[15:0]) +
	( 15'sd 8450) * $signed(input_fmap_72[15:0]) +
	( 14'sd 6378) * $signed(input_fmap_73[15:0]) +
	( 14'sd 6858) * $signed(input_fmap_74[15:0]) +
	( 16'sd 19965) * $signed(input_fmap_75[15:0]) +
	( 15'sd 10335) * $signed(input_fmap_76[15:0]) +
	( 12'sd 1302) * $signed(input_fmap_77[15:0]) +
	( 15'sd 14972) * $signed(input_fmap_78[15:0]) +
	( 15'sd 11037) * $signed(input_fmap_79[15:0]) +
	( 16'sd 17084) * $signed(input_fmap_80[15:0]) +
	( 10'sd 259) * $signed(input_fmap_81[15:0]) +
	( 15'sd 15296) * $signed(input_fmap_82[15:0]) +
	( 15'sd 8326) * $signed(input_fmap_83[15:0]) +
	( 15'sd 9270) * $signed(input_fmap_84[15:0]) +
	( 16'sd 22736) * $signed(input_fmap_85[15:0]) +
	( 15'sd 10856) * $signed(input_fmap_86[15:0]) +
	( 16'sd 30398) * $signed(input_fmap_87[15:0]) +
	( 16'sd 27975) * $signed(input_fmap_88[15:0]) +
	( 13'sd 3602) * $signed(input_fmap_89[15:0]) +
	( 16'sd 30596) * $signed(input_fmap_90[15:0]) +
	( 14'sd 5645) * $signed(input_fmap_91[15:0]) +
	( 14'sd 7431) * $signed(input_fmap_92[15:0]) +
	( 13'sd 2661) * $signed(input_fmap_93[15:0]) +
	( 16'sd 26501) * $signed(input_fmap_94[15:0]) +
	( 16'sd 19757) * $signed(input_fmap_95[15:0]) +
	( 14'sd 6667) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27196) * $signed(input_fmap_97[15:0]) +
	( 14'sd 5161) * $signed(input_fmap_98[15:0]) +
	( 16'sd 16873) * $signed(input_fmap_99[15:0]) +
	( 16'sd 18791) * $signed(input_fmap_100[15:0]) +
	( 16'sd 30087) * $signed(input_fmap_101[15:0]) +
	( 16'sd 25183) * $signed(input_fmap_102[15:0]) +
	( 14'sd 4595) * $signed(input_fmap_103[15:0]) +
	( 16'sd 17514) * $signed(input_fmap_104[15:0]) +
	( 16'sd 18097) * $signed(input_fmap_105[15:0]) +
	( 16'sd 32060) * $signed(input_fmap_106[15:0]) +
	( 15'sd 14139) * $signed(input_fmap_107[15:0]) +
	( 16'sd 29591) * $signed(input_fmap_108[15:0]) +
	( 15'sd 11112) * $signed(input_fmap_109[15:0]) +
	( 16'sd 25608) * $signed(input_fmap_110[15:0]) +
	( 16'sd 32230) * $signed(input_fmap_111[15:0]) +
	( 16'sd 32592) * $signed(input_fmap_112[15:0]) +
	( 14'sd 7665) * $signed(input_fmap_113[15:0]) +
	( 16'sd 30174) * $signed(input_fmap_114[15:0]) +
	( 16'sd 17567) * $signed(input_fmap_115[15:0]) +
	( 15'sd 13056) * $signed(input_fmap_116[15:0]) +
	( 15'sd 13128) * $signed(input_fmap_117[15:0]) +
	( 16'sd 27366) * $signed(input_fmap_118[15:0]) +
	( 16'sd 19017) * $signed(input_fmap_119[15:0]) +
	( 15'sd 11290) * $signed(input_fmap_120[15:0]) +
	( 16'sd 27667) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9917) * $signed(input_fmap_122[15:0]) +
	( 15'sd 9845) * $signed(input_fmap_123[15:0]) +
	( 16'sd 24048) * $signed(input_fmap_124[15:0]) +
	( 13'sd 2840) * $signed(input_fmap_125[15:0]) +
	( 16'sd 23344) * $signed(input_fmap_126[15:0]) +
	( 16'sd 24555) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 13'sd 3210) * $signed(input_fmap_0[15:0]) +
	( 15'sd 8981) * $signed(input_fmap_1[15:0]) +
	( 16'sd 28925) * $signed(input_fmap_2[15:0]) +
	( 16'sd 22502) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30345) * $signed(input_fmap_4[15:0]) +
	( 16'sd 31528) * $signed(input_fmap_5[15:0]) +
	( 15'sd 11827) * $signed(input_fmap_6[15:0]) +
	( 16'sd 28082) * $signed(input_fmap_7[15:0]) +
	( 15'sd 11823) * $signed(input_fmap_8[15:0]) +
	( 16'sd 17273) * $signed(input_fmap_9[15:0]) +
	( 16'sd 32527) * $signed(input_fmap_10[15:0]) +
	( 16'sd 29514) * $signed(input_fmap_11[15:0]) +
	( 15'sd 13256) * $signed(input_fmap_12[15:0]) +
	( 14'sd 4812) * $signed(input_fmap_13[15:0]) +
	( 16'sd 24780) * $signed(input_fmap_14[15:0]) +
	( 16'sd 21343) * $signed(input_fmap_15[15:0]) +
	( 14'sd 6533) * $signed(input_fmap_16[15:0]) +
	( 12'sd 1294) * $signed(input_fmap_17[15:0]) +
	( 15'sd 12400) * $signed(input_fmap_18[15:0]) +
	( 16'sd 20205) * $signed(input_fmap_19[15:0]) +
	( 16'sd 20190) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17410) * $signed(input_fmap_21[15:0]) +
	( 16'sd 29551) * $signed(input_fmap_22[15:0]) +
	( 16'sd 16518) * $signed(input_fmap_23[15:0]) +
	( 14'sd 4318) * $signed(input_fmap_24[15:0]) +
	( 9'sd 197) * $signed(input_fmap_25[15:0]) +
	( 16'sd 25512) * $signed(input_fmap_26[15:0]) +
	( 16'sd 25832) * $signed(input_fmap_27[15:0]) +
	( 16'sd 29229) * $signed(input_fmap_28[15:0]) +
	( 16'sd 22549) * $signed(input_fmap_29[15:0]) +
	( 16'sd 23228) * $signed(input_fmap_30[15:0]) +
	( 16'sd 19355) * $signed(input_fmap_31[15:0]) +
	( 15'sd 9047) * $signed(input_fmap_32[15:0]) +
	( 16'sd 26210) * $signed(input_fmap_33[15:0]) +
	( 14'sd 5602) * $signed(input_fmap_34[15:0]) +
	( 13'sd 2903) * $signed(input_fmap_35[15:0]) +
	( 16'sd 30647) * $signed(input_fmap_36[15:0]) +
	( 11'sd 820) * $signed(input_fmap_37[15:0]) +
	( 16'sd 28881) * $signed(input_fmap_38[15:0]) +
	( 14'sd 4545) * $signed(input_fmap_39[15:0]) +
	( 15'sd 13765) * $signed(input_fmap_40[15:0]) +
	( 15'sd 12385) * $signed(input_fmap_41[15:0]) +
	( 16'sd 30074) * $signed(input_fmap_42[15:0]) +
	( 16'sd 28559) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31789) * $signed(input_fmap_44[15:0]) +
	( 15'sd 14802) * $signed(input_fmap_45[15:0]) +
	( 16'sd 20133) * $signed(input_fmap_46[15:0]) +
	( 16'sd 22461) * $signed(input_fmap_47[15:0]) +
	( 16'sd 17451) * $signed(input_fmap_48[15:0]) +
	( 12'sd 1991) * $signed(input_fmap_49[15:0]) +
	( 15'sd 9961) * $signed(input_fmap_50[15:0]) +
	( 16'sd 22738) * $signed(input_fmap_51[15:0]) +
	( 14'sd 7812) * $signed(input_fmap_52[15:0]) +
	( 15'sd 13835) * $signed(input_fmap_53[15:0]) +
	( 16'sd 24131) * $signed(input_fmap_54[15:0]) +
	( 16'sd 18273) * $signed(input_fmap_55[15:0]) +
	( 15'sd 11150) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17980) * $signed(input_fmap_57[15:0]) +
	( 16'sd 22437) * $signed(input_fmap_58[15:0]) +
	( 16'sd 21402) * $signed(input_fmap_59[15:0]) +
	( 16'sd 25368) * $signed(input_fmap_60[15:0]) +
	( 13'sd 3932) * $signed(input_fmap_61[15:0]) +
	( 16'sd 22150) * $signed(input_fmap_62[15:0]) +
	( 15'sd 10807) * $signed(input_fmap_63[15:0]) +
	( 16'sd 18050) * $signed(input_fmap_64[15:0]) +
	( 16'sd 29541) * $signed(input_fmap_65[15:0]) +
	( 16'sd 17275) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28135) * $signed(input_fmap_67[15:0]) +
	( 11'sd 549) * $signed(input_fmap_68[15:0]) +
	( 15'sd 15302) * $signed(input_fmap_69[15:0]) +
	( 15'sd 14338) * $signed(input_fmap_70[15:0]) +
	( 15'sd 12692) * $signed(input_fmap_71[15:0]) +
	( 14'sd 5619) * $signed(input_fmap_72[15:0]) +
	( 16'sd 20623) * $signed(input_fmap_73[15:0]) +
	( 14'sd 7456) * $signed(input_fmap_74[15:0]) +
	( 15'sd 13302) * $signed(input_fmap_75[15:0]) +
	( 15'sd 13140) * $signed(input_fmap_76[15:0]) +
	( 14'sd 7641) * $signed(input_fmap_77[15:0]) +
	( 13'sd 2977) * $signed(input_fmap_78[15:0]) +
	( 16'sd 30713) * $signed(input_fmap_79[15:0]) +
	( 14'sd 8191) * $signed(input_fmap_80[15:0]) +
	( 15'sd 10668) * $signed(input_fmap_81[15:0]) +
	( 16'sd 29204) * $signed(input_fmap_82[15:0]) +
	( 14'sd 7167) * $signed(input_fmap_83[15:0]) +
	( 16'sd 26795) * $signed(input_fmap_84[15:0]) +
	( 16'sd 31937) * $signed(input_fmap_85[15:0]) +
	( 15'sd 8697) * $signed(input_fmap_86[15:0]) +
	( 16'sd 22732) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6193) * $signed(input_fmap_88[15:0]) +
	( 15'sd 9611) * $signed(input_fmap_89[15:0]) +
	( 12'sd 1448) * $signed(input_fmap_90[15:0]) +
	( 16'sd 17117) * $signed(input_fmap_91[15:0]) +
	( 15'sd 13642) * $signed(input_fmap_92[15:0]) +
	( 16'sd 25601) * $signed(input_fmap_93[15:0]) +
	( 15'sd 12819) * $signed(input_fmap_94[15:0]) +
	( 15'sd 8874) * $signed(input_fmap_95[15:0]) +
	( 15'sd 12309) * $signed(input_fmap_96[15:0]) +
	( 15'sd 15571) * $signed(input_fmap_97[15:0]) +
	( 13'sd 3571) * $signed(input_fmap_98[15:0]) +
	( 16'sd 27327) * $signed(input_fmap_99[15:0]) +
	( 15'sd 14976) * $signed(input_fmap_100[15:0]) +
	( 16'sd 28198) * $signed(input_fmap_101[15:0]) +
	( 16'sd 32224) * $signed(input_fmap_102[15:0]) +
	( 16'sd 32568) * $signed(input_fmap_103[15:0]) +
	( 13'sd 2260) * $signed(input_fmap_104[15:0]) +
	( 14'sd 7858) * $signed(input_fmap_105[15:0]) +
	( 15'sd 9702) * $signed(input_fmap_106[15:0]) +
	( 16'sd 30485) * $signed(input_fmap_107[15:0]) +
	( 16'sd 32401) * $signed(input_fmap_108[15:0]) +
	( 16'sd 31930) * $signed(input_fmap_109[15:0]) +
	( 16'sd 21768) * $signed(input_fmap_110[15:0]) +
	( 16'sd 25071) * $signed(input_fmap_111[15:0]) +
	( 15'sd 11523) * $signed(input_fmap_112[15:0]) +
	( 12'sd 1436) * $signed(input_fmap_113[15:0]) +
	( 16'sd 24220) * $signed(input_fmap_114[15:0]) +
	( 13'sd 2257) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15701) * $signed(input_fmap_116[15:0]) +
	( 13'sd 4053) * $signed(input_fmap_117[15:0]) +
	( 15'sd 13591) * $signed(input_fmap_118[15:0]) +
	( 14'sd 5501) * $signed(input_fmap_119[15:0]) +
	( 10'sd 260) * $signed(input_fmap_120[15:0]) +
	( 16'sd 30039) * $signed(input_fmap_121[15:0]) +
	( 16'sd 30742) * $signed(input_fmap_122[15:0]) +
	( 11'sd 742) * $signed(input_fmap_123[15:0]) +
	( 16'sd 23937) * $signed(input_fmap_124[15:0]) +
	( 15'sd 15640) * $signed(input_fmap_125[15:0]) +
	( 11'sd 726) * $signed(input_fmap_126[15:0]) +
	( 12'sd 2020) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 15'sd 10908) * $signed(input_fmap_0[15:0]) +
	( 13'sd 2575) * $signed(input_fmap_1[15:0]) +
	( 15'sd 10162) * $signed(input_fmap_2[15:0]) +
	( 16'sd 29501) * $signed(input_fmap_3[15:0]) +
	( 16'sd 29709) * $signed(input_fmap_4[15:0]) +
	( 12'sd 1773) * $signed(input_fmap_5[15:0]) +
	( 16'sd 19334) * $signed(input_fmap_6[15:0]) +
	( 13'sd 3841) * $signed(input_fmap_7[15:0]) +
	( 16'sd 32760) * $signed(input_fmap_8[15:0]) +
	( 16'sd 26025) * $signed(input_fmap_9[15:0]) +
	( 15'sd 9924) * $signed(input_fmap_10[15:0]) +
	( 15'sd 14694) * $signed(input_fmap_11[15:0]) +
	( 16'sd 30020) * $signed(input_fmap_12[15:0]) +
	( 15'sd 12625) * $signed(input_fmap_13[15:0]) +
	( 16'sd 19709) * $signed(input_fmap_14[15:0]) +
	( 15'sd 12640) * $signed(input_fmap_15[15:0]) +
	( 16'sd 28045) * $signed(input_fmap_16[15:0]) +
	( 15'sd 15547) * $signed(input_fmap_17[15:0]) +
	( 15'sd 13293) * $signed(input_fmap_18[15:0]) +
	( 16'sd 25655) * $signed(input_fmap_19[15:0]) +
	( 13'sd 3844) * $signed(input_fmap_20[15:0]) +
	( 16'sd 25415) * $signed(input_fmap_21[15:0]) +
	( 16'sd 19136) * $signed(input_fmap_22[15:0]) +
	( 16'sd 31404) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17680) * $signed(input_fmap_24[15:0]) +
	( 16'sd 31154) * $signed(input_fmap_25[15:0]) +
	( 15'sd 14067) * $signed(input_fmap_26[15:0]) +
	( 16'sd 25796) * $signed(input_fmap_27[15:0]) +
	( 12'sd 1561) * $signed(input_fmap_28[15:0]) +
	( 16'sd 18095) * $signed(input_fmap_29[15:0]) +
	( 15'sd 12025) * $signed(input_fmap_30[15:0]) +
	( 14'sd 6227) * $signed(input_fmap_31[15:0]) +
	( 14'sd 6313) * $signed(input_fmap_32[15:0]) +
	( 16'sd 25714) * $signed(input_fmap_33[15:0]) +
	( 15'sd 13955) * $signed(input_fmap_34[15:0]) +
	( 16'sd 28152) * $signed(input_fmap_35[15:0]) +
	( 16'sd 24836) * $signed(input_fmap_36[15:0]) +
	( 16'sd 27654) * $signed(input_fmap_37[15:0]) +
	( 16'sd 23984) * $signed(input_fmap_38[15:0]) +
	( 13'sd 3294) * $signed(input_fmap_39[15:0]) +
	( 13'sd 3348) * $signed(input_fmap_40[15:0]) +
	( 15'sd 12671) * $signed(input_fmap_41[15:0]) +
	( 16'sd 27622) * $signed(input_fmap_42[15:0]) +
	( 15'sd 15824) * $signed(input_fmap_43[15:0]) +
	( 15'sd 11603) * $signed(input_fmap_44[15:0]) +
	( 16'sd 20411) * $signed(input_fmap_45[15:0]) +
	( 16'sd 31707) * $signed(input_fmap_46[15:0]) +
	( 16'sd 16980) * $signed(input_fmap_47[15:0]) +
	( 16'sd 25115) * $signed(input_fmap_48[15:0]) +
	( 15'sd 15740) * $signed(input_fmap_49[15:0]) +
	( 16'sd 19608) * $signed(input_fmap_50[15:0]) +
	( 16'sd 30976) * $signed(input_fmap_51[15:0]) +
	( 16'sd 18127) * $signed(input_fmap_52[15:0]) +
	( 14'sd 7060) * $signed(input_fmap_53[15:0]) +
	( 15'sd 8750) * $signed(input_fmap_54[15:0]) +
	( 16'sd 27593) * $signed(input_fmap_55[15:0]) +
	( 16'sd 23238) * $signed(input_fmap_56[15:0]) +
	( 14'sd 6552) * $signed(input_fmap_57[15:0]) +
	( 16'sd 19999) * $signed(input_fmap_58[15:0]) +
	( 13'sd 2902) * $signed(input_fmap_59[15:0]) +
	( 16'sd 26292) * $signed(input_fmap_60[15:0]) +
	( 16'sd 24488) * $signed(input_fmap_61[15:0]) +
	( 15'sd 11101) * $signed(input_fmap_62[15:0]) +
	( 16'sd 16428) * $signed(input_fmap_63[15:0]) +
	( 14'sd 5223) * $signed(input_fmap_64[15:0]) +
	( 13'sd 2407) * $signed(input_fmap_65[15:0]) +
	( 15'sd 9169) * $signed(input_fmap_66[15:0]) +
	( 16'sd 30597) * $signed(input_fmap_67[15:0]) +
	( 16'sd 17294) * $signed(input_fmap_68[15:0]) +
	( 14'sd 5278) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31809) * $signed(input_fmap_70[15:0]) +
	( 15'sd 14970) * $signed(input_fmap_71[15:0]) +
	( 16'sd 32271) * $signed(input_fmap_72[15:0]) +
	( 13'sd 3518) * $signed(input_fmap_73[15:0]) +
	( 13'sd 2887) * $signed(input_fmap_74[15:0]) +
	( 15'sd 14735) * $signed(input_fmap_75[15:0]) +
	( 16'sd 29419) * $signed(input_fmap_76[15:0]) +
	( 16'sd 21021) * $signed(input_fmap_77[15:0]) +
	( 16'sd 16762) * $signed(input_fmap_78[15:0]) +
	( 13'sd 2625) * $signed(input_fmap_79[15:0]) +
	( 15'sd 14924) * $signed(input_fmap_80[15:0]) +
	( 16'sd 31152) * $signed(input_fmap_81[15:0]) +
	( 16'sd 16961) * $signed(input_fmap_82[15:0]) +
	( 15'sd 10402) * $signed(input_fmap_83[15:0]) +
	( 16'sd 30796) * $signed(input_fmap_84[15:0]) +
	( 16'sd 28127) * $signed(input_fmap_85[15:0]) +
	( 16'sd 19375) * $signed(input_fmap_86[15:0]) +
	( 16'sd 27297) * $signed(input_fmap_87[15:0]) +
	( 16'sd 22203) * $signed(input_fmap_88[15:0]) +
	( 16'sd 24552) * $signed(input_fmap_89[15:0]) +
	( 14'sd 6226) * $signed(input_fmap_90[15:0]) +
	( 15'sd 15674) * $signed(input_fmap_91[15:0]) +
	( 16'sd 18675) * $signed(input_fmap_92[15:0]) +
	( 16'sd 26196) * $signed(input_fmap_93[15:0]) +
	( 16'sd 28013) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25655) * $signed(input_fmap_95[15:0]) +
	( 16'sd 17382) * $signed(input_fmap_96[15:0]) +
	( 16'sd 25964) * $signed(input_fmap_97[15:0]) +
	( 16'sd 31872) * $signed(input_fmap_98[15:0]) +
	( 16'sd 29765) * $signed(input_fmap_99[15:0]) +
	( 15'sd 9692) * $signed(input_fmap_100[15:0]) +
	( 16'sd 22033) * $signed(input_fmap_101[15:0]) +
	( 11'sd 546) * $signed(input_fmap_102[15:0]) +
	( 16'sd 20820) * $signed(input_fmap_103[15:0]) +
	( 16'sd 30600) * $signed(input_fmap_104[15:0]) +
	( 12'sd 1427) * $signed(input_fmap_105[15:0]) +
	( 16'sd 27567) * $signed(input_fmap_106[15:0]) +
	( 16'sd 16818) * $signed(input_fmap_107[15:0]) +
	( 15'sd 13314) * $signed(input_fmap_108[15:0]) +
	( 15'sd 8921) * $signed(input_fmap_109[15:0]) +
	( 14'sd 4911) * $signed(input_fmap_110[15:0]) +
	( 14'sd 8066) * $signed(input_fmap_111[15:0]) +
	( 15'sd 11753) * $signed(input_fmap_112[15:0]) +
	( 15'sd 10954) * $signed(input_fmap_113[15:0]) +
	( 15'sd 11918) * $signed(input_fmap_114[15:0]) +
	( 16'sd 27355) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15319) * $signed(input_fmap_116[15:0]) +
	( 16'sd 20654) * $signed(input_fmap_117[15:0]) +
	( 16'sd 16497) * $signed(input_fmap_118[15:0]) +
	( 15'sd 12482) * $signed(input_fmap_119[15:0]) +
	( 14'sd 5958) * $signed(input_fmap_120[15:0]) +
	( 16'sd 18229) * $signed(input_fmap_121[15:0]) +
	( 13'sd 2790) * $signed(input_fmap_122[15:0]) +
	( 15'sd 14243) * $signed(input_fmap_123[15:0]) +
	( 13'sd 3464) * $signed(input_fmap_124[15:0]) +
	( 12'sd 1613) * $signed(input_fmap_125[15:0]) +
	( 16'sd 20069) * $signed(input_fmap_126[15:0]) +
	( 15'sd 10198) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 15'sd 11362) * $signed(input_fmap_0[15:0]) +
	( 15'sd 9979) * $signed(input_fmap_1[15:0]) +
	( 16'sd 20193) * $signed(input_fmap_2[15:0]) +
	( 15'sd 11556) * $signed(input_fmap_3[15:0]) +
	( 16'sd 22061) * $signed(input_fmap_4[15:0]) +
	( 15'sd 14381) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2133) * $signed(input_fmap_6[15:0]) +
	( 16'sd 31811) * $signed(input_fmap_7[15:0]) +
	( 14'sd 7914) * $signed(input_fmap_8[15:0]) +
	( 14'sd 5272) * $signed(input_fmap_9[15:0]) +
	( 16'sd 31541) * $signed(input_fmap_10[15:0]) +
	( 14'sd 7679) * $signed(input_fmap_11[15:0]) +
	( 16'sd 30215) * $signed(input_fmap_12[15:0]) +
	( 15'sd 13565) * $signed(input_fmap_13[15:0]) +
	( 16'sd 23988) * $signed(input_fmap_14[15:0]) +
	( 16'sd 31917) * $signed(input_fmap_15[15:0]) +
	( 16'sd 22386) * $signed(input_fmap_16[15:0]) +
	( 15'sd 12407) * $signed(input_fmap_17[15:0]) +
	( 12'sd 1050) * $signed(input_fmap_18[15:0]) +
	( 15'sd 8207) * $signed(input_fmap_19[15:0]) +
	( 12'sd 1586) * $signed(input_fmap_20[15:0]) +
	( 14'sd 4330) * $signed(input_fmap_21[15:0]) +
	( 16'sd 18287) * $signed(input_fmap_22[15:0]) +
	( 16'sd 17563) * $signed(input_fmap_23[15:0]) +
	( 14'sd 7099) * $signed(input_fmap_24[15:0]) +
	( 15'sd 8600) * $signed(input_fmap_25[15:0]) +
	( 16'sd 16589) * $signed(input_fmap_26[15:0]) +
	( 16'sd 24381) * $signed(input_fmap_27[15:0]) +
	( 15'sd 8929) * $signed(input_fmap_28[15:0]) +
	( 9'sd 214) * $signed(input_fmap_29[15:0]) +
	( 10'sd 393) * $signed(input_fmap_30[15:0]) +
	( 16'sd 18372) * $signed(input_fmap_31[15:0]) +
	( 16'sd 26682) * $signed(input_fmap_32[15:0]) +
	( 13'sd 3329) * $signed(input_fmap_33[15:0]) +
	( 16'sd 22456) * $signed(input_fmap_34[15:0]) +
	( 15'sd 10550) * $signed(input_fmap_35[15:0]) +
	( 16'sd 28870) * $signed(input_fmap_36[15:0]) +
	( 16'sd 31103) * $signed(input_fmap_37[15:0]) +
	( 16'sd 22297) * $signed(input_fmap_38[15:0]) +
	( 13'sd 3945) * $signed(input_fmap_39[15:0]) +
	( 9'sd 240) * $signed(input_fmap_40[15:0]) +
	( 16'sd 32628) * $signed(input_fmap_41[15:0]) +
	( 15'sd 13918) * $signed(input_fmap_42[15:0]) +
	( 16'sd 26374) * $signed(input_fmap_43[15:0]) +
	( 16'sd 22109) * $signed(input_fmap_44[15:0]) +
	( 16'sd 21627) * $signed(input_fmap_45[15:0]) +
	( 16'sd 22406) * $signed(input_fmap_46[15:0]) +
	( 14'sd 6513) * $signed(input_fmap_47[15:0]) +
	( 16'sd 26568) * $signed(input_fmap_48[15:0]) +
	( 16'sd 16587) * $signed(input_fmap_49[15:0]) +
	( 16'sd 32325) * $signed(input_fmap_50[15:0]) +
	( 15'sd 14508) * $signed(input_fmap_51[15:0]) +
	( 16'sd 16433) * $signed(input_fmap_52[15:0]) +
	( 15'sd 15618) * $signed(input_fmap_53[15:0]) +
	( 15'sd 16061) * $signed(input_fmap_54[15:0]) +
	( 14'sd 5328) * $signed(input_fmap_55[15:0]) +
	( 15'sd 12204) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17932) * $signed(input_fmap_57[15:0]) +
	( 15'sd 13529) * $signed(input_fmap_58[15:0]) +
	( 14'sd 5461) * $signed(input_fmap_59[15:0]) +
	( 15'sd 12442) * $signed(input_fmap_60[15:0]) +
	( 16'sd 18412) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3578) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20812) * $signed(input_fmap_63[15:0]) +
	( 16'sd 30471) * $signed(input_fmap_64[15:0]) +
	( 16'sd 18804) * $signed(input_fmap_65[15:0]) +
	( 15'sd 12594) * $signed(input_fmap_66[15:0]) +
	( 16'sd 17322) * $signed(input_fmap_67[15:0]) +
	( 15'sd 12523) * $signed(input_fmap_68[15:0]) +
	( 12'sd 1059) * $signed(input_fmap_69[15:0]) +
	( 16'sd 17676) * $signed(input_fmap_70[15:0]) +
	( 16'sd 26620) * $signed(input_fmap_71[15:0]) +
	( 15'sd 8473) * $signed(input_fmap_72[15:0]) +
	( 13'sd 2667) * $signed(input_fmap_73[15:0]) +
	( 12'sd 1628) * $signed(input_fmap_74[15:0]) +
	( 15'sd 9586) * $signed(input_fmap_75[15:0]) +
	( 16'sd 22696) * $signed(input_fmap_76[15:0]) +
	( 13'sd 3992) * $signed(input_fmap_77[15:0]) +
	( 16'sd 25332) * $signed(input_fmap_78[15:0]) +
	( 16'sd 23832) * $signed(input_fmap_79[15:0]) +
	( 16'sd 27047) * $signed(input_fmap_80[15:0]) +
	( 16'sd 17814) * $signed(input_fmap_81[15:0]) +
	( 16'sd 17036) * $signed(input_fmap_82[15:0]) +
	( 16'sd 27799) * $signed(input_fmap_83[15:0]) +
	( 14'sd 5663) * $signed(input_fmap_84[15:0]) +
	( 16'sd 17287) * $signed(input_fmap_85[15:0]) +
	( 14'sd 4752) * $signed(input_fmap_86[15:0]) +
	( 14'sd 5356) * $signed(input_fmap_87[15:0]) +
	( 13'sd 2479) * $signed(input_fmap_88[15:0]) +
	( 14'sd 4829) * $signed(input_fmap_89[15:0]) +
	( 16'sd 26127) * $signed(input_fmap_90[15:0]) +
	( 14'sd 5472) * $signed(input_fmap_91[15:0]) +
	( 10'sd 507) * $signed(input_fmap_92[15:0]) +
	( 16'sd 27122) * $signed(input_fmap_93[15:0]) +
	( 16'sd 16579) * $signed(input_fmap_94[15:0]) +
	( 13'sd 3551) * $signed(input_fmap_95[15:0]) +
	( 16'sd 32437) * $signed(input_fmap_96[15:0]) +
	( 16'sd 28687) * $signed(input_fmap_97[15:0]) +
	( 16'sd 16855) * $signed(input_fmap_98[15:0]) +
	( 13'sd 3230) * $signed(input_fmap_99[15:0]) +
	( 15'sd 13973) * $signed(input_fmap_100[15:0]) +
	( 15'sd 9763) * $signed(input_fmap_101[15:0]) +
	( 15'sd 16020) * $signed(input_fmap_102[15:0]) +
	( 16'sd 30083) * $signed(input_fmap_103[15:0]) +
	( 16'sd 27285) * $signed(input_fmap_104[15:0]) +
	( 15'sd 15677) * $signed(input_fmap_105[15:0]) +
	( 15'sd 10833) * $signed(input_fmap_106[15:0]) +
	( 16'sd 20627) * $signed(input_fmap_107[15:0]) +
	( 15'sd 13704) * $signed(input_fmap_108[15:0]) +
	( 16'sd 16947) * $signed(input_fmap_109[15:0]) +
	( 16'sd 24881) * $signed(input_fmap_110[15:0]) +
	( 16'sd 31770) * $signed(input_fmap_111[15:0]) +
	( 16'sd 27029) * $signed(input_fmap_112[15:0]) +
	( 15'sd 11000) * $signed(input_fmap_113[15:0]) +
	( 15'sd 10596) * $signed(input_fmap_114[15:0]) +
	( 16'sd 26881) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15681) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27397) * $signed(input_fmap_117[15:0]) +
	( 16'sd 30908) * $signed(input_fmap_118[15:0]) +
	( 14'sd 7962) * $signed(input_fmap_119[15:0]) +
	( 13'sd 2314) * $signed(input_fmap_120[15:0]) +
	( 16'sd 20103) * $signed(input_fmap_121[15:0]) +
	( 15'sd 8512) * $signed(input_fmap_122[15:0]) +
	( 16'sd 19224) * $signed(input_fmap_123[15:0]) +
	( 15'sd 13226) * $signed(input_fmap_124[15:0]) +
	( 15'sd 12588) * $signed(input_fmap_125[15:0]) +
	( 16'sd 27908) * $signed(input_fmap_126[15:0]) +
	( 15'sd 11645) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 16'sd 31471) * $signed(input_fmap_0[15:0]) +
	( 16'sd 31689) * $signed(input_fmap_1[15:0]) +
	( 13'sd 2164) * $signed(input_fmap_2[15:0]) +
	( 16'sd 23841) * $signed(input_fmap_3[15:0]) +
	( 16'sd 19317) * $signed(input_fmap_4[15:0]) +
	( 15'sd 10293) * $signed(input_fmap_5[15:0]) +
	( 15'sd 10679) * $signed(input_fmap_6[15:0]) +
	( 16'sd 23170) * $signed(input_fmap_7[15:0]) +
	( 14'sd 6892) * $signed(input_fmap_8[15:0]) +
	( 16'sd 23189) * $signed(input_fmap_9[15:0]) +
	( 13'sd 3882) * $signed(input_fmap_10[15:0]) +
	( 16'sd 18078) * $signed(input_fmap_11[15:0]) +
	( 16'sd 28564) * $signed(input_fmap_12[15:0]) +
	( 16'sd 28761) * $signed(input_fmap_13[15:0]) +
	( 16'sd 26656) * $signed(input_fmap_14[15:0]) +
	( 16'sd 24188) * $signed(input_fmap_15[15:0]) +
	( 16'sd 24072) * $signed(input_fmap_16[15:0]) +
	( 16'sd 16897) * $signed(input_fmap_17[15:0]) +
	( 15'sd 15039) * $signed(input_fmap_18[15:0]) +
	( 16'sd 19419) * $signed(input_fmap_19[15:0]) +
	( 15'sd 9546) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17117) * $signed(input_fmap_21[15:0]) +
	( 15'sd 10573) * $signed(input_fmap_22[15:0]) +
	( 15'sd 10992) * $signed(input_fmap_23[15:0]) +
	( 16'sd 31431) * $signed(input_fmap_24[15:0]) +
	( 16'sd 24481) * $signed(input_fmap_25[15:0]) +
	( 14'sd 5350) * $signed(input_fmap_26[15:0]) +
	( 14'sd 7028) * $signed(input_fmap_27[15:0]) +
	( 15'sd 10262) * $signed(input_fmap_28[15:0]) +
	( 15'sd 9704) * $signed(input_fmap_29[15:0]) +
	( 16'sd 18186) * $signed(input_fmap_30[15:0]) +
	( 16'sd 26462) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28944) * $signed(input_fmap_32[15:0]) +
	( 16'sd 20528) * $signed(input_fmap_33[15:0]) +
	( 16'sd 30865) * $signed(input_fmap_34[15:0]) +
	( 16'sd 22435) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11026) * $signed(input_fmap_36[15:0]) +
	( 16'sd 18454) * $signed(input_fmap_37[15:0]) +
	( 16'sd 21468) * $signed(input_fmap_38[15:0]) +
	( 14'sd 4283) * $signed(input_fmap_39[15:0]) +
	( 15'sd 8525) * $signed(input_fmap_40[15:0]) +
	( 16'sd 31184) * $signed(input_fmap_41[15:0]) +
	( 14'sd 8171) * $signed(input_fmap_42[15:0]) +
	( 14'sd 7925) * $signed(input_fmap_43[15:0]) +
	( 16'sd 21639) * $signed(input_fmap_44[15:0]) +
	( 15'sd 14145) * $signed(input_fmap_45[15:0]) +
	( 15'sd 10350) * $signed(input_fmap_46[15:0]) +
	( 16'sd 16906) * $signed(input_fmap_47[15:0]) +
	( 12'sd 1782) * $signed(input_fmap_48[15:0]) +
	( 15'sd 14731) * $signed(input_fmap_49[15:0]) +
	( 16'sd 17349) * $signed(input_fmap_50[15:0]) +
	( 16'sd 32650) * $signed(input_fmap_51[15:0]) +
	( 16'sd 28682) * $signed(input_fmap_52[15:0]) +
	( 15'sd 11257) * $signed(input_fmap_53[15:0]) +
	( 16'sd 28472) * $signed(input_fmap_54[15:0]) +
	( 16'sd 23736) * $signed(input_fmap_55[15:0]) +
	( 16'sd 26943) * $signed(input_fmap_56[15:0]) +
	( 16'sd 32192) * $signed(input_fmap_57[15:0]) +
	( 16'sd 19658) * $signed(input_fmap_58[15:0]) +
	( 16'sd 21854) * $signed(input_fmap_59[15:0]) +
	( 16'sd 16794) * $signed(input_fmap_60[15:0]) +
	( 16'sd 17968) * $signed(input_fmap_61[15:0]) +
	( 16'sd 24645) * $signed(input_fmap_62[15:0]) +
	( 13'sd 3491) * $signed(input_fmap_63[15:0]) +
	( 16'sd 28311) * $signed(input_fmap_64[15:0]) +
	( 16'sd 20711) * $signed(input_fmap_65[15:0]) +
	( 15'sd 9880) * $signed(input_fmap_66[15:0]) +
	( 16'sd 18598) * $signed(input_fmap_67[15:0]) +
	( 14'sd 6750) * $signed(input_fmap_68[15:0]) +
	( 12'sd 1471) * $signed(input_fmap_69[15:0]) +
	( 16'sd 25442) * $signed(input_fmap_70[15:0]) +
	( 16'sd 23235) * $signed(input_fmap_71[15:0]) +
	( 16'sd 27348) * $signed(input_fmap_72[15:0]) +
	( 16'sd 20293) * $signed(input_fmap_73[15:0]) +
	( 16'sd 30585) * $signed(input_fmap_74[15:0]) +
	( 15'sd 14894) * $signed(input_fmap_75[15:0]) +
	( 15'sd 10285) * $signed(input_fmap_76[15:0]) +
	( 16'sd 23346) * $signed(input_fmap_77[15:0]) +
	( 15'sd 10193) * $signed(input_fmap_78[15:0]) +
	( 16'sd 17771) * $signed(input_fmap_79[15:0]) +
	( 16'sd 19995) * $signed(input_fmap_80[15:0]) +
	( 14'sd 4689) * $signed(input_fmap_81[15:0]) +
	( 15'sd 12356) * $signed(input_fmap_82[15:0]) +
	( 16'sd 31775) * $signed(input_fmap_83[15:0]) +
	( 11'sd 909) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24652) * $signed(input_fmap_85[15:0]) +
	( 14'sd 4293) * $signed(input_fmap_86[15:0]) +
	( 15'sd 12346) * $signed(input_fmap_87[15:0]) +
	( 16'sd 19008) * $signed(input_fmap_88[15:0]) +
	( 16'sd 24606) * $signed(input_fmap_89[15:0]) +
	( 15'sd 11625) * $signed(input_fmap_90[15:0]) +
	( 16'sd 22136) * $signed(input_fmap_91[15:0]) +
	( 14'sd 6162) * $signed(input_fmap_92[15:0]) +
	( 14'sd 7080) * $signed(input_fmap_93[15:0]) +
	( 14'sd 7960) * $signed(input_fmap_94[15:0]) +
	( 16'sd 21852) * $signed(input_fmap_95[15:0]) +
	( 15'sd 10364) * $signed(input_fmap_96[15:0]) +
	( 16'sd 16962) * $signed(input_fmap_97[15:0]) +
	( 15'sd 11917) * $signed(input_fmap_98[15:0]) +
	( 16'sd 20413) * $signed(input_fmap_99[15:0]) +
	( 14'sd 4734) * $signed(input_fmap_100[15:0]) +
	( 13'sd 2482) * $signed(input_fmap_101[15:0]) +
	( 16'sd 21265) * $signed(input_fmap_102[15:0]) +
	( 16'sd 16985) * $signed(input_fmap_103[15:0]) +
	( 16'sd 28746) * $signed(input_fmap_104[15:0]) +
	( 14'sd 6566) * $signed(input_fmap_105[15:0]) +
	( 16'sd 17136) * $signed(input_fmap_106[15:0]) +
	( 12'sd 1721) * $signed(input_fmap_107[15:0]) +
	( 16'sd 29088) * $signed(input_fmap_108[15:0]) +
	( 16'sd 32351) * $signed(input_fmap_109[15:0]) +
	( 16'sd 29918) * $signed(input_fmap_110[15:0]) +
	( 16'sd 29333) * $signed(input_fmap_111[15:0]) +
	( 16'sd 28200) * $signed(input_fmap_112[15:0]) +
	( 13'sd 3926) * $signed(input_fmap_113[15:0]) +
	( 16'sd 18131) * $signed(input_fmap_114[15:0]) +
	( 16'sd 28578) * $signed(input_fmap_115[15:0]) +
	( 12'sd 1676) * $signed(input_fmap_116[15:0]) +
	( 14'sd 4818) * $signed(input_fmap_117[15:0]) +
	( 14'sd 5196) * $signed(input_fmap_118[15:0]) +
	( 15'sd 11539) * $signed(input_fmap_119[15:0]) +
	( 16'sd 19482) * $signed(input_fmap_120[15:0]) +
	( 16'sd 28650) * $signed(input_fmap_121[15:0]) +
	( 16'sd 23222) * $signed(input_fmap_122[15:0]) +
	( 16'sd 30827) * $signed(input_fmap_123[15:0]) +
	( 15'sd 15651) * $signed(input_fmap_124[15:0]) +
	( 15'sd 11046) * $signed(input_fmap_125[15:0]) +
	( 10'sd 411) * $signed(input_fmap_126[15:0]) +
	( 16'sd 25152) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 14'sd 6735) * $signed(input_fmap_0[15:0]) +
	( 14'sd 5486) * $signed(input_fmap_1[15:0]) +
	( 15'sd 8811) * $signed(input_fmap_2[15:0]) +
	( 16'sd 27421) * $signed(input_fmap_3[15:0]) +
	( 16'sd 18469) * $signed(input_fmap_4[15:0]) +
	( 16'sd 25326) * $signed(input_fmap_5[15:0]) +
	( 15'sd 10054) * $signed(input_fmap_6[15:0]) +
	( 14'sd 7727) * $signed(input_fmap_7[15:0]) +
	( 16'sd 17521) * $signed(input_fmap_8[15:0]) +
	( 13'sd 2640) * $signed(input_fmap_9[15:0]) +
	( 16'sd 31239) * $signed(input_fmap_10[15:0]) +
	( 15'sd 15708) * $signed(input_fmap_11[15:0]) +
	( 16'sd 28445) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24303) * $signed(input_fmap_13[15:0]) +
	( 14'sd 6890) * $signed(input_fmap_14[15:0]) +
	( 16'sd 21454) * $signed(input_fmap_15[15:0]) +
	( 15'sd 13149) * $signed(input_fmap_16[15:0]) +
	( 13'sd 3959) * $signed(input_fmap_17[15:0]) +
	( 14'sd 4505) * $signed(input_fmap_18[15:0]) +
	( 16'sd 20169) * $signed(input_fmap_19[15:0]) +
	( 13'sd 2668) * $signed(input_fmap_20[15:0]) +
	( 16'sd 26140) * $signed(input_fmap_21[15:0]) +
	( 16'sd 18505) * $signed(input_fmap_22[15:0]) +
	( 16'sd 21116) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17579) * $signed(input_fmap_24[15:0]) +
	( 15'sd 10465) * $signed(input_fmap_25[15:0]) +
	( 13'sd 3285) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9583) * $signed(input_fmap_27[15:0]) +
	( 16'sd 23755) * $signed(input_fmap_28[15:0]) +
	( 14'sd 7453) * $signed(input_fmap_29[15:0]) +
	( 12'sd 2025) * $signed(input_fmap_30[15:0]) +
	( 16'sd 29442) * $signed(input_fmap_31[15:0]) +
	( 16'sd 22941) * $signed(input_fmap_32[15:0]) +
	( 15'sd 16375) * $signed(input_fmap_33[15:0]) +
	( 14'sd 6918) * $signed(input_fmap_34[15:0]) +
	( 16'sd 25734) * $signed(input_fmap_35[15:0]) +
	( 16'sd 16654) * $signed(input_fmap_36[15:0]) +
	( 15'sd 8664) * $signed(input_fmap_37[15:0]) +
	( 16'sd 31855) * $signed(input_fmap_38[15:0]) +
	( 16'sd 17750) * $signed(input_fmap_39[15:0]) +
	( 15'sd 15702) * $signed(input_fmap_40[15:0]) +
	( 16'sd 18999) * $signed(input_fmap_41[15:0]) +
	( 14'sd 5910) * $signed(input_fmap_42[15:0]) +
	( 16'sd 26631) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31185) * $signed(input_fmap_44[15:0]) +
	( 14'sd 4804) * $signed(input_fmap_45[15:0]) +
	( 16'sd 21482) * $signed(input_fmap_46[15:0]) +
	( 12'sd 1701) * $signed(input_fmap_47[15:0]) +
	( 15'sd 10382) * $signed(input_fmap_48[15:0]) +
	( 15'sd 11276) * $signed(input_fmap_49[15:0]) +
	( 16'sd 29361) * $signed(input_fmap_50[15:0]) +
	( 10'sd 277) * $signed(input_fmap_51[15:0]) +
	( 16'sd 28448) * $signed(input_fmap_52[15:0]) +
	( 14'sd 5819) * $signed(input_fmap_53[15:0]) +
	( 15'sd 11749) * $signed(input_fmap_54[15:0]) +
	( 16'sd 24082) * $signed(input_fmap_55[15:0]) +
	( 16'sd 21739) * $signed(input_fmap_56[15:0]) +
	( 15'sd 12114) * $signed(input_fmap_57[15:0]) +
	( 13'sd 3905) * $signed(input_fmap_58[15:0]) +
	( 15'sd 13868) * $signed(input_fmap_59[15:0]) +
	( 16'sd 26546) * $signed(input_fmap_60[15:0]) +
	( 15'sd 15232) * $signed(input_fmap_61[15:0]) +
	( 15'sd 15775) * $signed(input_fmap_62[15:0]) +
	( 16'sd 19016) * $signed(input_fmap_63[15:0]) +
	( 15'sd 16206) * $signed(input_fmap_64[15:0]) +
	( 16'sd 28161) * $signed(input_fmap_65[15:0]) +
	( 13'sd 2425) * $signed(input_fmap_66[15:0]) +
	( 16'sd 19676) * $signed(input_fmap_67[15:0]) +
	( 13'sd 2540) * $signed(input_fmap_68[15:0]) +
	( 16'sd 18132) * $signed(input_fmap_69[15:0]) +
	( 16'sd 27199) * $signed(input_fmap_70[15:0]) +
	( 16'sd 30879) * $signed(input_fmap_71[15:0]) +
	( 14'sd 5368) * $signed(input_fmap_72[15:0]) +
	( 14'sd 5219) * $signed(input_fmap_73[15:0]) +
	( 16'sd 17641) * $signed(input_fmap_74[15:0]) +
	( 16'sd 28427) * $signed(input_fmap_75[15:0]) +
	( 14'sd 6337) * $signed(input_fmap_76[15:0]) +
	( 15'sd 8869) * $signed(input_fmap_77[15:0]) +
	( 14'sd 4865) * $signed(input_fmap_78[15:0]) +
	( 16'sd 19957) * $signed(input_fmap_79[15:0]) +
	( 15'sd 8760) * $signed(input_fmap_80[15:0]) +
	( 16'sd 19609) * $signed(input_fmap_81[15:0]) +
	( 16'sd 16802) * $signed(input_fmap_82[15:0]) +
	( 14'sd 7104) * $signed(input_fmap_83[15:0]) +
	( 16'sd 17241) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24915) * $signed(input_fmap_85[15:0]) +
	( 15'sd 15441) * $signed(input_fmap_86[15:0]) +
	( 16'sd 23042) * $signed(input_fmap_87[15:0]) +
	( 16'sd 21057) * $signed(input_fmap_88[15:0]) +
	( 16'sd 17218) * $signed(input_fmap_89[15:0]) +
	( 16'sd 24331) * $signed(input_fmap_90[15:0]) +
	( 15'sd 12284) * $signed(input_fmap_91[15:0]) +
	( 15'sd 15897) * $signed(input_fmap_92[15:0]) +
	( 13'sd 2763) * $signed(input_fmap_93[15:0]) +
	( 16'sd 31107) * $signed(input_fmap_94[15:0]) +
	( 15'sd 13712) * $signed(input_fmap_95[15:0]) +
	( 13'sd 3585) * $signed(input_fmap_96[15:0]) +
	( 15'sd 8488) * $signed(input_fmap_97[15:0]) +
	( 14'sd 4470) * $signed(input_fmap_98[15:0]) +
	( 15'sd 14555) * $signed(input_fmap_99[15:0]) +
	( 15'sd 11285) * $signed(input_fmap_100[15:0]) +
	( 16'sd 20953) * $signed(input_fmap_101[15:0]) +
	( 16'sd 30982) * $signed(input_fmap_102[15:0]) +
	( 14'sd 4182) * $signed(input_fmap_103[15:0]) +
	( 16'sd 22053) * $signed(input_fmap_104[15:0]) +
	( 14'sd 5442) * $signed(input_fmap_105[15:0]) +
	( 13'sd 2622) * $signed(input_fmap_106[15:0]) +
	( 15'sd 10972) * $signed(input_fmap_107[15:0]) +
	( 16'sd 32260) * $signed(input_fmap_108[15:0]) +
	( 15'sd 10548) * $signed(input_fmap_109[15:0]) +
	( 16'sd 17848) * $signed(input_fmap_110[15:0]) +
	( 16'sd 29515) * $signed(input_fmap_111[15:0]) +
	( 15'sd 8833) * $signed(input_fmap_112[15:0]) +
	( 10'sd 410) * $signed(input_fmap_113[15:0]) +
	( 15'sd 13129) * $signed(input_fmap_114[15:0]) +
	( 16'sd 31452) * $signed(input_fmap_115[15:0]) +
	( 16'sd 31419) * $signed(input_fmap_116[15:0]) +
	( 14'sd 6027) * $signed(input_fmap_117[15:0]) +
	( 16'sd 21389) * $signed(input_fmap_118[15:0]) +
	( 16'sd 21393) * $signed(input_fmap_119[15:0]) +
	( 15'sd 11815) * $signed(input_fmap_120[15:0]) +
	( 16'sd 26518) * $signed(input_fmap_121[15:0]) +
	( 16'sd 27829) * $signed(input_fmap_122[15:0]) +
	( 16'sd 29878) * $signed(input_fmap_123[15:0]) +
	( 10'sd 297) * $signed(input_fmap_124[15:0]) +
	( 16'sd 21845) * $signed(input_fmap_125[15:0]) +
	( 13'sd 3390) * $signed(input_fmap_126[15:0]) +
	( 8'sd 90) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 16'sd 17324) * $signed(input_fmap_0[15:0]) +
	( 15'sd 13788) * $signed(input_fmap_1[15:0]) +
	( 16'sd 23930) * $signed(input_fmap_2[15:0]) +
	( 16'sd 24780) * $signed(input_fmap_3[15:0]) +
	( 16'sd 17970) * $signed(input_fmap_4[15:0]) +
	( 16'sd 19233) * $signed(input_fmap_5[15:0]) +
	( 15'sd 12555) * $signed(input_fmap_6[15:0]) +
	( 16'sd 30636) * $signed(input_fmap_7[15:0]) +
	( 16'sd 25920) * $signed(input_fmap_8[15:0]) +
	( 15'sd 13018) * $signed(input_fmap_9[15:0]) +
	( 16'sd 17306) * $signed(input_fmap_10[15:0]) +
	( 16'sd 22013) * $signed(input_fmap_11[15:0]) +
	( 15'sd 11506) * $signed(input_fmap_12[15:0]) +
	( 14'sd 7154) * $signed(input_fmap_13[15:0]) +
	( 14'sd 7263) * $signed(input_fmap_14[15:0]) +
	( 15'sd 10102) * $signed(input_fmap_15[15:0]) +
	( 14'sd 4230) * $signed(input_fmap_16[15:0]) +
	( 16'sd 16720) * $signed(input_fmap_17[15:0]) +
	( 16'sd 28233) * $signed(input_fmap_18[15:0]) +
	( 16'sd 17931) * $signed(input_fmap_19[15:0]) +
	( 13'sd 4030) * $signed(input_fmap_20[15:0]) +
	( 16'sd 30456) * $signed(input_fmap_21[15:0]) +
	( 15'sd 13269) * $signed(input_fmap_22[15:0]) +
	( 15'sd 9665) * $signed(input_fmap_23[15:0]) +
	( 15'sd 15410) * $signed(input_fmap_24[15:0]) +
	( 15'sd 12272) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22221) * $signed(input_fmap_26[15:0]) +
	( 16'sd 18000) * $signed(input_fmap_27[15:0]) +
	( 16'sd 18056) * $signed(input_fmap_28[15:0]) +
	( 16'sd 16433) * $signed(input_fmap_29[15:0]) +
	( 16'sd 22709) * $signed(input_fmap_30[15:0]) +
	( 15'sd 14061) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28190) * $signed(input_fmap_32[15:0]) +
	( 15'sd 16222) * $signed(input_fmap_33[15:0]) +
	( 13'sd 2608) * $signed(input_fmap_34[15:0]) +
	( 16'sd 22839) * $signed(input_fmap_35[15:0]) +
	( 16'sd 17252) * $signed(input_fmap_36[15:0]) +
	( 16'sd 18047) * $signed(input_fmap_37[15:0]) +
	( 15'sd 11146) * $signed(input_fmap_38[15:0]) +
	( 16'sd 30015) * $signed(input_fmap_39[15:0]) +
	( 12'sd 1783) * $signed(input_fmap_40[15:0]) +
	( 16'sd 25881) * $signed(input_fmap_41[15:0]) +
	( 16'sd 25350) * $signed(input_fmap_42[15:0]) +
	( 16'sd 30969) * $signed(input_fmap_43[15:0]) +
	( 16'sd 19301) * $signed(input_fmap_44[15:0]) +
	( 14'sd 5854) * $signed(input_fmap_45[15:0]) +
	( 15'sd 13040) * $signed(input_fmap_46[15:0]) +
	( 13'sd 3363) * $signed(input_fmap_47[15:0]) +
	( 12'sd 1817) * $signed(input_fmap_48[15:0]) +
	( 16'sd 17335) * $signed(input_fmap_49[15:0]) +
	( 16'sd 18315) * $signed(input_fmap_50[15:0]) +
	( 14'sd 6125) * $signed(input_fmap_51[15:0]) +
	( 16'sd 31991) * $signed(input_fmap_52[15:0]) +
	( 15'sd 8905) * $signed(input_fmap_53[15:0]) +
	( 14'sd 5271) * $signed(input_fmap_54[15:0]) +
	( 16'sd 22902) * $signed(input_fmap_55[15:0]) +
	( 16'sd 32746) * $signed(input_fmap_56[15:0]) +
	( 16'sd 30658) * $signed(input_fmap_57[15:0]) +
	( 16'sd 31699) * $signed(input_fmap_58[15:0]) +
	( 16'sd 23264) * $signed(input_fmap_59[15:0]) +
	( 16'sd 16528) * $signed(input_fmap_60[15:0]) +
	( 16'sd 27894) * $signed(input_fmap_61[15:0]) +
	( 15'sd 15036) * $signed(input_fmap_62[15:0]) +
	( 16'sd 30262) * $signed(input_fmap_63[15:0]) +
	( 15'sd 15765) * $signed(input_fmap_64[15:0]) +
	( 14'sd 5147) * $signed(input_fmap_65[15:0]) +
	( 16'sd 31840) * $signed(input_fmap_66[15:0]) +
	( 14'sd 4243) * $signed(input_fmap_67[15:0]) +
	( 15'sd 14326) * $signed(input_fmap_68[15:0]) +
	( 15'sd 14877) * $signed(input_fmap_69[15:0]) +
	( 10'sd 256) * $signed(input_fmap_70[15:0]) +
	( 16'sd 27159) * $signed(input_fmap_71[15:0]) +
	( 16'sd 24913) * $signed(input_fmap_72[15:0]) +
	( 12'sd 1898) * $signed(input_fmap_73[15:0]) +
	( 16'sd 21973) * $signed(input_fmap_74[15:0]) +
	( 16'sd 22019) * $signed(input_fmap_75[15:0]) +
	( 14'sd 4361) * $signed(input_fmap_76[15:0]) +
	( 14'sd 5878) * $signed(input_fmap_77[15:0]) +
	( 14'sd 7676) * $signed(input_fmap_78[15:0]) +
	( 16'sd 24760) * $signed(input_fmap_79[15:0]) +
	( 16'sd 23749) * $signed(input_fmap_80[15:0]) +
	( 16'sd 21546) * $signed(input_fmap_81[15:0]) +
	( 16'sd 25643) * $signed(input_fmap_82[15:0]) +
	( 15'sd 15033) * $signed(input_fmap_83[15:0]) +
	( 16'sd 31933) * $signed(input_fmap_84[15:0]) +
	( 15'sd 12334) * $signed(input_fmap_85[15:0]) +
	( 16'sd 22068) * $signed(input_fmap_86[15:0]) +
	( 16'sd 24407) * $signed(input_fmap_87[15:0]) +
	( 14'sd 4285) * $signed(input_fmap_88[15:0]) +
	( 16'sd 23036) * $signed(input_fmap_89[15:0]) +
	( 16'sd 20211) * $signed(input_fmap_90[15:0]) +
	( 16'sd 17466) * $signed(input_fmap_91[15:0]) +
	( 16'sd 32737) * $signed(input_fmap_92[15:0]) +
	( 16'sd 23004) * $signed(input_fmap_93[15:0]) +
	( 16'sd 16944) * $signed(input_fmap_94[15:0]) +
	( 16'sd 30933) * $signed(input_fmap_95[15:0]) +
	( 16'sd 19686) * $signed(input_fmap_96[15:0]) +
	( 14'sd 5998) * $signed(input_fmap_97[15:0]) +
	( 16'sd 17732) * $signed(input_fmap_98[15:0]) +
	( 16'sd 19535) * $signed(input_fmap_99[15:0]) +
	( 15'sd 11140) * $signed(input_fmap_100[15:0]) +
	( 16'sd 17586) * $signed(input_fmap_101[15:0]) +
	( 16'sd 20662) * $signed(input_fmap_102[15:0]) +
	( 12'sd 2017) * $signed(input_fmap_103[15:0]) +
	( 16'sd 25254) * $signed(input_fmap_104[15:0]) +
	( 15'sd 10806) * $signed(input_fmap_105[15:0]) +
	( 16'sd 23321) * $signed(input_fmap_106[15:0]) +
	( 16'sd 29456) * $signed(input_fmap_107[15:0]) +
	( 16'sd 31856) * $signed(input_fmap_108[15:0]) +
	( 16'sd 18082) * $signed(input_fmap_109[15:0]) +
	( 16'sd 24532) * $signed(input_fmap_110[15:0]) +
	( 16'sd 31871) * $signed(input_fmap_111[15:0]) +
	( 15'sd 14007) * $signed(input_fmap_112[15:0]) +
	( 14'sd 8184) * $signed(input_fmap_113[15:0]) +
	( 15'sd 10349) * $signed(input_fmap_114[15:0]) +
	( 16'sd 27471) * $signed(input_fmap_115[15:0]) +
	( 16'sd 22457) * $signed(input_fmap_116[15:0]) +
	( 16'sd 28831) * $signed(input_fmap_117[15:0]) +
	( 16'sd 21185) * $signed(input_fmap_118[15:0]) +
	( 13'sd 2381) * $signed(input_fmap_119[15:0]) +
	( 14'sd 6173) * $signed(input_fmap_120[15:0]) +
	( 16'sd 21458) * $signed(input_fmap_121[15:0]) +
	( 16'sd 26614) * $signed(input_fmap_122[15:0]) +
	( 16'sd 22155) * $signed(input_fmap_123[15:0]) +
	( 16'sd 32608) * $signed(input_fmap_124[15:0]) +
	( 15'sd 9868) * $signed(input_fmap_125[15:0]) +
	( 15'sd 11009) * $signed(input_fmap_126[15:0]) +
	( 16'sd 21739) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 13'sd 2555) * $signed(input_fmap_0[15:0]) +
	( 16'sd 28169) * $signed(input_fmap_1[15:0]) +
	( 16'sd 21580) * $signed(input_fmap_2[15:0]) +
	( 16'sd 32220) * $signed(input_fmap_3[15:0]) +
	( 16'sd 29865) * $signed(input_fmap_4[15:0]) +
	( 16'sd 28584) * $signed(input_fmap_5[15:0]) +
	( 8'sd 78) * $signed(input_fmap_6[15:0]) +
	( 16'sd 32032) * $signed(input_fmap_7[15:0]) +
	( 16'sd 16816) * $signed(input_fmap_8[15:0]) +
	( 14'sd 4435) * $signed(input_fmap_9[15:0]) +
	( 15'sd 12445) * $signed(input_fmap_10[15:0]) +
	( 16'sd 16543) * $signed(input_fmap_11[15:0]) +
	( 13'sd 3011) * $signed(input_fmap_12[15:0]) +
	( 16'sd 29851) * $signed(input_fmap_13[15:0]) +
	( 15'sd 16334) * $signed(input_fmap_14[15:0]) +
	( 15'sd 13076) * $signed(input_fmap_15[15:0]) +
	( 13'sd 2868) * $signed(input_fmap_16[15:0]) +
	( 10'sd 428) * $signed(input_fmap_17[15:0]) +
	( 16'sd 20519) * $signed(input_fmap_18[15:0]) +
	( 15'sd 10401) * $signed(input_fmap_19[15:0]) +
	( 14'sd 6742) * $signed(input_fmap_20[15:0]) +
	( 15'sd 10144) * $signed(input_fmap_21[15:0]) +
	( 16'sd 25154) * $signed(input_fmap_22[15:0]) +
	( 15'sd 13001) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17458) * $signed(input_fmap_24[15:0]) +
	( 16'sd 30725) * $signed(input_fmap_25[15:0]) +
	( 16'sd 19034) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9445) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24537) * $signed(input_fmap_28[15:0]) +
	( 12'sd 1594) * $signed(input_fmap_29[15:0]) +
	( 14'sd 4848) * $signed(input_fmap_30[15:0]) +
	( 16'sd 22376) * $signed(input_fmap_31[15:0]) +
	( 16'sd 23860) * $signed(input_fmap_32[15:0]) +
	( 15'sd 16276) * $signed(input_fmap_33[15:0]) +
	( 15'sd 15360) * $signed(input_fmap_34[15:0]) +
	( 16'sd 31421) * $signed(input_fmap_35[15:0]) +
	( 14'sd 5589) * $signed(input_fmap_36[15:0]) +
	( 16'sd 32128) * $signed(input_fmap_37[15:0]) +
	( 11'sd 778) * $signed(input_fmap_38[15:0]) +
	( 16'sd 23521) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6830) * $signed(input_fmap_40[15:0]) +
	( 16'sd 28385) * $signed(input_fmap_41[15:0]) +
	( 16'sd 32581) * $signed(input_fmap_42[15:0]) +
	( 14'sd 6606) * $signed(input_fmap_43[15:0]) +
	( 16'sd 32386) * $signed(input_fmap_44[15:0]) +
	( 16'sd 24354) * $signed(input_fmap_45[15:0]) +
	( 16'sd 19433) * $signed(input_fmap_46[15:0]) +
	( 15'sd 11165) * $signed(input_fmap_47[15:0]) +
	( 14'sd 4417) * $signed(input_fmap_48[15:0]) +
	( 13'sd 2679) * $signed(input_fmap_49[15:0]) +
	( 16'sd 23982) * $signed(input_fmap_50[15:0]) +
	( 15'sd 8472) * $signed(input_fmap_51[15:0]) +
	( 16'sd 18861) * $signed(input_fmap_52[15:0]) +
	( 15'sd 11093) * $signed(input_fmap_53[15:0]) +
	( 15'sd 14971) * $signed(input_fmap_54[15:0]) +
	( 15'sd 8561) * $signed(input_fmap_55[15:0]) +
	( 16'sd 22880) * $signed(input_fmap_56[15:0]) +
	( 13'sd 3840) * $signed(input_fmap_57[15:0]) +
	( 14'sd 7352) * $signed(input_fmap_58[15:0]) +
	( 16'sd 30698) * $signed(input_fmap_59[15:0]) +
	( 16'sd 22854) * $signed(input_fmap_60[15:0]) +
	( 16'sd 32337) * $signed(input_fmap_61[15:0]) +
	( 16'sd 18076) * $signed(input_fmap_62[15:0]) +
	( 16'sd 17752) * $signed(input_fmap_63[15:0]) +
	( 15'sd 15819) * $signed(input_fmap_64[15:0]) +
	( 16'sd 28483) * $signed(input_fmap_65[15:0]) +
	( 13'sd 2796) * $signed(input_fmap_66[15:0]) +
	( 16'sd 27337) * $signed(input_fmap_67[15:0]) +
	( 16'sd 25143) * $signed(input_fmap_68[15:0]) +
	( 14'sd 5941) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31747) * $signed(input_fmap_70[15:0]) +
	( 15'sd 15763) * $signed(input_fmap_71[15:0]) +
	( 15'sd 8435) * $signed(input_fmap_72[15:0]) +
	( 16'sd 25269) * $signed(input_fmap_73[15:0]) +
	( 16'sd 28028) * $signed(input_fmap_74[15:0]) +
	( 16'sd 28833) * $signed(input_fmap_75[15:0]) +
	( 16'sd 28958) * $signed(input_fmap_76[15:0]) +
	( 15'sd 8819) * $signed(input_fmap_77[15:0]) +
	( 16'sd 17744) * $signed(input_fmap_78[15:0]) +
	( 15'sd 11035) * $signed(input_fmap_79[15:0]) +
	( 16'sd 19597) * $signed(input_fmap_80[15:0]) +
	( 16'sd 21500) * $signed(input_fmap_81[15:0]) +
	( 12'sd 1898) * $signed(input_fmap_82[15:0]) +
	( 15'sd 12126) * $signed(input_fmap_83[15:0]) +
	( 16'sd 23536) * $signed(input_fmap_84[15:0]) +
	( 14'sd 5969) * $signed(input_fmap_85[15:0]) +
	( 14'sd 5428) * $signed(input_fmap_86[15:0]) +
	( 16'sd 20720) * $signed(input_fmap_87[15:0]) +
	( 16'sd 27663) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5827) * $signed(input_fmap_89[15:0]) +
	( 15'sd 13540) * $signed(input_fmap_90[15:0]) +
	( 13'sd 3146) * $signed(input_fmap_91[15:0]) +
	( 15'sd 11499) * $signed(input_fmap_92[15:0]) +
	( 16'sd 27195) * $signed(input_fmap_93[15:0]) +
	( 16'sd 23000) * $signed(input_fmap_94[15:0]) +
	( 14'sd 4230) * $signed(input_fmap_95[15:0]) +
	( 16'sd 21863) * $signed(input_fmap_96[15:0]) +
	( 15'sd 8591) * $signed(input_fmap_97[15:0]) +
	( 14'sd 7764) * $signed(input_fmap_98[15:0]) +
	( 16'sd 19597) * $signed(input_fmap_99[15:0]) +
	( 16'sd 19837) * $signed(input_fmap_100[15:0]) +
	( 16'sd 26694) * $signed(input_fmap_101[15:0]) +
	( 15'sd 12490) * $signed(input_fmap_102[15:0]) +
	( 15'sd 14240) * $signed(input_fmap_103[15:0]) +
	( 15'sd 9903) * $signed(input_fmap_104[15:0]) +
	( 14'sd 5369) * $signed(input_fmap_105[15:0]) +
	( 16'sd 31211) * $signed(input_fmap_106[15:0]) +
	( 16'sd 18999) * $signed(input_fmap_107[15:0]) +
	( 16'sd 24023) * $signed(input_fmap_108[15:0]) +
	( 16'sd 28829) * $signed(input_fmap_109[15:0]) +
	( 14'sd 5724) * $signed(input_fmap_110[15:0]) +
	( 16'sd 26284) * $signed(input_fmap_111[15:0]) +
	( 13'sd 3078) * $signed(input_fmap_112[15:0]) +
	( 16'sd 22008) * $signed(input_fmap_113[15:0]) +
	( 7'sd 59) * $signed(input_fmap_114[15:0]) +
	( 14'sd 6937) * $signed(input_fmap_115[15:0]) +
	( 16'sd 20091) * $signed(input_fmap_116[15:0]) +
	( 14'sd 7503) * $signed(input_fmap_117[15:0]) +
	( 14'sd 7779) * $signed(input_fmap_118[15:0]) +
	( 16'sd 24806) * $signed(input_fmap_119[15:0]) +
	( 15'sd 15219) * $signed(input_fmap_120[15:0]) +
	( 13'sd 3481) * $signed(input_fmap_121[15:0]) +
	( 16'sd 29534) * $signed(input_fmap_122[15:0]) +
	( 14'sd 6297) * $signed(input_fmap_123[15:0]) +
	( 15'sd 13868) * $signed(input_fmap_124[15:0]) +
	( 16'sd 31941) * $signed(input_fmap_125[15:0]) +
	( 15'sd 9824) * $signed(input_fmap_126[15:0]) +
	( 16'sd 26962) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 16'sd 18873) * $signed(input_fmap_0[15:0]) +
	( 14'sd 7622) * $signed(input_fmap_1[15:0]) +
	( 13'sd 2288) * $signed(input_fmap_2[15:0]) +
	( 15'sd 13276) * $signed(input_fmap_3[15:0]) +
	( 16'sd 17341) * $signed(input_fmap_4[15:0]) +
	( 16'sd 20890) * $signed(input_fmap_5[15:0]) +
	( 15'sd 11337) * $signed(input_fmap_6[15:0]) +
	( 16'sd 20705) * $signed(input_fmap_7[15:0]) +
	( 16'sd 22888) * $signed(input_fmap_8[15:0]) +
	( 16'sd 29677) * $signed(input_fmap_9[15:0]) +
	( 15'sd 8517) * $signed(input_fmap_10[15:0]) +
	( 15'sd 9849) * $signed(input_fmap_11[15:0]) +
	( 14'sd 7000) * $signed(input_fmap_12[15:0]) +
	( 14'sd 6395) * $signed(input_fmap_13[15:0]) +
	( 10'sd 416) * $signed(input_fmap_14[15:0]) +
	( 13'sd 2120) * $signed(input_fmap_15[15:0]) +
	( 16'sd 21427) * $signed(input_fmap_16[15:0]) +
	( 16'sd 29996) * $signed(input_fmap_17[15:0]) +
	( 16'sd 31332) * $signed(input_fmap_18[15:0]) +
	( 16'sd 26980) * $signed(input_fmap_19[15:0]) +
	( 15'sd 11233) * $signed(input_fmap_20[15:0]) +
	( 16'sd 23490) * $signed(input_fmap_21[15:0]) +
	( 14'sd 5762) * $signed(input_fmap_22[15:0]) +
	( 16'sd 32019) * $signed(input_fmap_23[15:0]) +
	( 13'sd 2689) * $signed(input_fmap_24[15:0]) +
	( 16'sd 29918) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22042) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9674) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24112) * $signed(input_fmap_28[15:0]) +
	( 15'sd 10593) * $signed(input_fmap_29[15:0]) +
	( 16'sd 27583) * $signed(input_fmap_30[15:0]) +
	( 14'sd 5360) * $signed(input_fmap_31[15:0]) +
	( 14'sd 4394) * $signed(input_fmap_32[15:0]) +
	( 16'sd 26465) * $signed(input_fmap_33[15:0]) +
	( 13'sd 2265) * $signed(input_fmap_34[15:0]) +
	( 11'sd 719) * $signed(input_fmap_35[15:0]) +
	( 16'sd 21443) * $signed(input_fmap_36[15:0]) +
	( 16'sd 31704) * $signed(input_fmap_37[15:0]) +
	( 16'sd 16491) * $signed(input_fmap_38[15:0]) +
	( 16'sd 32052) * $signed(input_fmap_39[15:0]) +
	( 15'sd 11219) * $signed(input_fmap_40[15:0]) +
	( 15'sd 12250) * $signed(input_fmap_41[15:0]) +
	( 16'sd 23831) * $signed(input_fmap_42[15:0]) +
	( 16'sd 24041) * $signed(input_fmap_43[15:0]) +
	( 16'sd 22505) * $signed(input_fmap_44[15:0]) +
	( 16'sd 21306) * $signed(input_fmap_45[15:0]) +
	( 15'sd 14919) * $signed(input_fmap_46[15:0]) +
	( 16'sd 30840) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13470) * $signed(input_fmap_48[15:0]) +
	( 13'sd 3226) * $signed(input_fmap_49[15:0]) +
	( 15'sd 9376) * $signed(input_fmap_50[15:0]) +
	( 16'sd 20500) * $signed(input_fmap_51[15:0]) +
	( 16'sd 24838) * $signed(input_fmap_52[15:0]) +
	( 15'sd 15176) * $signed(input_fmap_53[15:0]) +
	( 16'sd 18231) * $signed(input_fmap_54[15:0]) +
	( 16'sd 21100) * $signed(input_fmap_55[15:0]) +
	( 13'sd 2342) * $signed(input_fmap_56[15:0]) +
	( 16'sd 28414) * $signed(input_fmap_57[15:0]) +
	( 16'sd 19680) * $signed(input_fmap_58[15:0]) +
	( 16'sd 18331) * $signed(input_fmap_59[15:0]) +
	( 16'sd 24960) * $signed(input_fmap_60[15:0]) +
	( 15'sd 8781) * $signed(input_fmap_61[15:0]) +
	( 16'sd 26017) * $signed(input_fmap_62[15:0]) +
	( 16'sd 24245) * $signed(input_fmap_63[15:0]) +
	( 15'sd 10877) * $signed(input_fmap_64[15:0]) +
	( 14'sd 6340) * $signed(input_fmap_65[15:0]) +
	( 16'sd 27763) * $signed(input_fmap_66[15:0]) +
	( 16'sd 19791) * $signed(input_fmap_67[15:0]) +
	( 16'sd 17138) * $signed(input_fmap_68[15:0]) +
	( 11'sd 894) * $signed(input_fmap_69[15:0]) +
	( 15'sd 9234) * $signed(input_fmap_70[15:0]) +
	( 14'sd 4921) * $signed(input_fmap_71[15:0]) +
	( 16'sd 29918) * $signed(input_fmap_72[15:0]) +
	( 16'sd 25155) * $signed(input_fmap_73[15:0]) +
	( 11'sd 860) * $signed(input_fmap_74[15:0]) +
	( 16'sd 17808) * $signed(input_fmap_75[15:0]) +
	( 16'sd 32282) * $signed(input_fmap_76[15:0]) +
	( 16'sd 24811) * $signed(input_fmap_77[15:0]) +
	( 13'sd 2237) * $signed(input_fmap_78[15:0]) +
	( 16'sd 17952) * $signed(input_fmap_79[15:0]) +
	( 14'sd 8098) * $signed(input_fmap_80[15:0]) +
	( 14'sd 5148) * $signed(input_fmap_81[15:0]) +
	( 16'sd 19404) * $signed(input_fmap_82[15:0]) +
	( 12'sd 1678) * $signed(input_fmap_83[15:0]) +
	( 15'sd 9107) * $signed(input_fmap_84[15:0]) +
	( 16'sd 22889) * $signed(input_fmap_85[15:0]) +
	( 16'sd 22296) * $signed(input_fmap_86[15:0]) +
	( 16'sd 32482) * $signed(input_fmap_87[15:0]) +
	( 16'sd 18051) * $signed(input_fmap_88[15:0]) +
	( 16'sd 29435) * $signed(input_fmap_89[15:0]) +
	( 15'sd 13402) * $signed(input_fmap_90[15:0]) +
	( 13'sd 2747) * $signed(input_fmap_91[15:0]) +
	( 14'sd 5284) * $signed(input_fmap_92[15:0]) +
	( 15'sd 9555) * $signed(input_fmap_93[15:0]) +
	( 16'sd 30810) * $signed(input_fmap_94[15:0]) +
	( 16'sd 22474) * $signed(input_fmap_95[15:0]) +
	( 13'sd 3649) * $signed(input_fmap_96[15:0]) +
	( 11'sd 981) * $signed(input_fmap_97[15:0]) +
	( 16'sd 22378) * $signed(input_fmap_98[15:0]) +
	( 11'sd 989) * $signed(input_fmap_99[15:0]) +
	( 16'sd 22588) * $signed(input_fmap_100[15:0]) +
	( 16'sd 25873) * $signed(input_fmap_101[15:0]) +
	( 16'sd 19741) * $signed(input_fmap_102[15:0]) +
	( 15'sd 9153) * $signed(input_fmap_103[15:0]) +
	( 14'sd 6750) * $signed(input_fmap_104[15:0]) +
	( 16'sd 27651) * $signed(input_fmap_105[15:0]) +
	( 15'sd 15003) * $signed(input_fmap_106[15:0]) +
	( 15'sd 9384) * $signed(input_fmap_107[15:0]) +
	( 14'sd 5694) * $signed(input_fmap_108[15:0]) +
	( 16'sd 30107) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22098) * $signed(input_fmap_110[15:0]) +
	( 15'sd 15760) * $signed(input_fmap_111[15:0]) +
	( 16'sd 32164) * $signed(input_fmap_112[15:0]) +
	( 16'sd 29520) * $signed(input_fmap_113[15:0]) +
	( 10'sd 364) * $signed(input_fmap_114[15:0]) +
	( 16'sd 18292) * $signed(input_fmap_115[15:0]) +
	( 15'sd 12742) * $signed(input_fmap_116[15:0]) +
	( 15'sd 14645) * $signed(input_fmap_117[15:0]) +
	( 16'sd 32389) * $signed(input_fmap_118[15:0]) +
	( 14'sd 7604) * $signed(input_fmap_119[15:0]) +
	( 16'sd 29506) * $signed(input_fmap_120[15:0]) +
	( 11'sd 673) * $signed(input_fmap_121[15:0]) +
	( 16'sd 24991) * $signed(input_fmap_122[15:0]) +
	( 15'sd 13780) * $signed(input_fmap_123[15:0]) +
	( 16'sd 16660) * $signed(input_fmap_124[15:0]) +
	( 15'sd 15905) * $signed(input_fmap_125[15:0]) +
	( 15'sd 16133) * $signed(input_fmap_126[15:0]) +
	( 15'sd 8525) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 16'sd 21782) * $signed(input_fmap_0[15:0]) +
	( 14'sd 5367) * $signed(input_fmap_1[15:0]) +
	( 15'sd 10549) * $signed(input_fmap_2[15:0]) +
	( 16'sd 18035) * $signed(input_fmap_3[15:0]) +
	( 12'sd 1761) * $signed(input_fmap_4[15:0]) +
	( 15'sd 8357) * $signed(input_fmap_5[15:0]) +
	( 15'sd 9450) * $signed(input_fmap_6[15:0]) +
	( 16'sd 21225) * $signed(input_fmap_7[15:0]) +
	( 16'sd 25063) * $signed(input_fmap_8[15:0]) +
	( 16'sd 16439) * $signed(input_fmap_9[15:0]) +
	( 16'sd 32270) * $signed(input_fmap_10[15:0]) +
	( 16'sd 16480) * $signed(input_fmap_11[15:0]) +
	( 16'sd 29953) * $signed(input_fmap_12[15:0]) +
	( 13'sd 2543) * $signed(input_fmap_13[15:0]) +
	( 16'sd 18014) * $signed(input_fmap_14[15:0]) +
	( 14'sd 6882) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10623) * $signed(input_fmap_16[15:0]) +
	( 16'sd 28061) * $signed(input_fmap_17[15:0]) +
	( 16'sd 25284) * $signed(input_fmap_18[15:0]) +
	( 16'sd 18041) * $signed(input_fmap_19[15:0]) +
	( 15'sd 8792) * $signed(input_fmap_20[15:0]) +
	( 11'sd 837) * $signed(input_fmap_21[15:0]) +
	( 15'sd 15933) * $signed(input_fmap_22[15:0]) +
	( 15'sd 9576) * $signed(input_fmap_23[15:0]) +
	( 15'sd 16345) * $signed(input_fmap_24[15:0]) +
	( 15'sd 8298) * $signed(input_fmap_25[15:0]) +
	( 14'sd 6912) * $signed(input_fmap_26[15:0]) +
	( 15'sd 11063) * $signed(input_fmap_27[15:0]) +
	( 16'sd 20173) * $signed(input_fmap_28[15:0]) +
	( 11'sd 566) * $signed(input_fmap_29[15:0]) +
	( 14'sd 7012) * $signed(input_fmap_30[15:0]) +
	( 16'sd 30161) * $signed(input_fmap_31[15:0]) +
	( 16'sd 18879) * $signed(input_fmap_32[15:0]) +
	( 14'sd 4486) * $signed(input_fmap_33[15:0]) +
	( 15'sd 8548) * $signed(input_fmap_34[15:0]) +
	( 16'sd 17412) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2291) * $signed(input_fmap_36[15:0]) +
	( 16'sd 27226) * $signed(input_fmap_37[15:0]) +
	( 16'sd 28285) * $signed(input_fmap_38[15:0]) +
	( 14'sd 6790) * $signed(input_fmap_39[15:0]) +
	( 16'sd 17683) * $signed(input_fmap_40[15:0]) +
	( 10'sd 339) * $signed(input_fmap_41[15:0]) +
	( 16'sd 18880) * $signed(input_fmap_42[15:0]) +
	( 11'sd 816) * $signed(input_fmap_43[15:0]) +
	( 16'sd 23457) * $signed(input_fmap_44[15:0]) +
	( 15'sd 15979) * $signed(input_fmap_45[15:0]) +
	( 13'sd 3747) * $signed(input_fmap_46[15:0]) +
	( 15'sd 12050) * $signed(input_fmap_47[15:0]) +
	( 15'sd 9447) * $signed(input_fmap_48[15:0]) +
	( 15'sd 13455) * $signed(input_fmap_49[15:0]) +
	( 16'sd 25527) * $signed(input_fmap_50[15:0]) +
	( 16'sd 19847) * $signed(input_fmap_51[15:0]) +
	( 15'sd 13840) * $signed(input_fmap_52[15:0]) +
	( 16'sd 28485) * $signed(input_fmap_53[15:0]) +
	( 16'sd 27536) * $signed(input_fmap_54[15:0]) +
	( 15'sd 13280) * $signed(input_fmap_55[15:0]) +
	( 16'sd 19992) * $signed(input_fmap_56[15:0]) +
	( 14'sd 5615) * $signed(input_fmap_57[15:0]) +
	( 16'sd 21695) * $signed(input_fmap_58[15:0]) +
	( 14'sd 7504) * $signed(input_fmap_59[15:0]) +
	( 16'sd 28644) * $signed(input_fmap_60[15:0]) +
	( 16'sd 24348) * $signed(input_fmap_61[15:0]) +
	( 13'sd 2509) * $signed(input_fmap_62[15:0]) +
	( 13'sd 3608) * $signed(input_fmap_63[15:0]) +
	( 16'sd 28930) * $signed(input_fmap_64[15:0]) +
	( 14'sd 4376) * $signed(input_fmap_65[15:0]) +
	( 15'sd 12961) * $signed(input_fmap_66[15:0]) +
	( 15'sd 9399) * $signed(input_fmap_67[15:0]) +
	( 16'sd 19207) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31568) * $signed(input_fmap_69[15:0]) +
	( 14'sd 5527) * $signed(input_fmap_70[15:0]) +
	( 15'sd 12369) * $signed(input_fmap_71[15:0]) +
	( 15'sd 12878) * $signed(input_fmap_72[15:0]) +
	( 16'sd 29098) * $signed(input_fmap_73[15:0]) +
	( 15'sd 10769) * $signed(input_fmap_74[15:0]) +
	( 16'sd 26997) * $signed(input_fmap_75[15:0]) +
	( 16'sd 27267) * $signed(input_fmap_76[15:0]) +
	( 15'sd 10140) * $signed(input_fmap_77[15:0]) +
	( 15'sd 11418) * $signed(input_fmap_78[15:0]) +
	( 16'sd 24518) * $signed(input_fmap_79[15:0]) +
	( 13'sd 3355) * $signed(input_fmap_80[15:0]) +
	( 16'sd 19918) * $signed(input_fmap_81[15:0]) +
	( 16'sd 28458) * $signed(input_fmap_82[15:0]) +
	( 12'sd 1094) * $signed(input_fmap_83[15:0]) +
	( 14'sd 7941) * $signed(input_fmap_84[15:0]) +
	( 14'sd 6084) * $signed(input_fmap_85[15:0]) +
	( 16'sd 22349) * $signed(input_fmap_86[15:0]) +
	( 16'sd 23440) * $signed(input_fmap_87[15:0]) +
	( 12'sd 1315) * $signed(input_fmap_88[15:0]) +
	( 16'sd 30674) * $signed(input_fmap_89[15:0]) +
	( 16'sd 22287) * $signed(input_fmap_90[15:0]) +
	( 16'sd 17884) * $signed(input_fmap_91[15:0]) +
	( 16'sd 20519) * $signed(input_fmap_92[15:0]) +
	( 14'sd 7566) * $signed(input_fmap_93[15:0]) +
	( 15'sd 12685) * $signed(input_fmap_94[15:0]) +
	( 12'sd 1833) * $signed(input_fmap_95[15:0]) +
	( 10'sd 256) * $signed(input_fmap_96[15:0]) +
	( 16'sd 31763) * $signed(input_fmap_97[15:0]) +
	( 16'sd 28601) * $signed(input_fmap_98[15:0]) +
	( 14'sd 4642) * $signed(input_fmap_99[15:0]) +
	( 15'sd 9415) * $signed(input_fmap_100[15:0]) +
	( 16'sd 25390) * $signed(input_fmap_101[15:0]) +
	( 15'sd 12999) * $signed(input_fmap_102[15:0]) +
	( 16'sd 22274) * $signed(input_fmap_103[15:0]) +
	( 14'sd 5273) * $signed(input_fmap_104[15:0]) +
	( 13'sd 3083) * $signed(input_fmap_105[15:0]) +
	( 15'sd 12247) * $signed(input_fmap_106[15:0]) +
	( 16'sd 22215) * $signed(input_fmap_107[15:0]) +
	( 16'sd 28005) * $signed(input_fmap_108[15:0]) +
	( 15'sd 13856) * $signed(input_fmap_109[15:0]) +
	( 12'sd 1213) * $signed(input_fmap_110[15:0]) +
	( 16'sd 20868) * $signed(input_fmap_111[15:0]) +
	( 16'sd 29136) * $signed(input_fmap_112[15:0]) +
	( 16'sd 29672) * $signed(input_fmap_113[15:0]) +
	( 16'sd 18782) * $signed(input_fmap_114[15:0]) +
	( 13'sd 2333) * $signed(input_fmap_115[15:0]) +
	( 16'sd 29067) * $signed(input_fmap_116[15:0]) +
	( 16'sd 18035) * $signed(input_fmap_117[15:0]) +
	( 16'sd 31590) * $signed(input_fmap_118[15:0]) +
	( 16'sd 21708) * $signed(input_fmap_119[15:0]) +
	( 16'sd 19169) * $signed(input_fmap_120[15:0]) +
	( 16'sd 17128) * $signed(input_fmap_121[15:0]) +
	( 13'sd 2253) * $signed(input_fmap_122[15:0]) +
	( 12'sd 1233) * $signed(input_fmap_123[15:0]) +
	( 16'sd 23497) * $signed(input_fmap_124[15:0]) +
	( 16'sd 29292) * $signed(input_fmap_125[15:0]) +
	( 16'sd 27807) * $signed(input_fmap_126[15:0]) +
	( 16'sd 19196) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 15'sd 13705) * $signed(input_fmap_0[15:0]) +
	( 15'sd 11737) * $signed(input_fmap_1[15:0]) +
	( 16'sd 27630) * $signed(input_fmap_2[15:0]) +
	( 16'sd 18764) * $signed(input_fmap_3[15:0]) +
	( 15'sd 11429) * $signed(input_fmap_4[15:0]) +
	( 15'sd 16185) * $signed(input_fmap_5[15:0]) +
	( 16'sd 21430) * $signed(input_fmap_6[15:0]) +
	( 16'sd 25323) * $signed(input_fmap_7[15:0]) +
	( 16'sd 23574) * $signed(input_fmap_8[15:0]) +
	( 16'sd 17563) * $signed(input_fmap_9[15:0]) +
	( 16'sd 30385) * $signed(input_fmap_10[15:0]) +
	( 14'sd 5873) * $signed(input_fmap_11[15:0]) +
	( 14'sd 6638) * $signed(input_fmap_12[15:0]) +
	( 15'sd 11451) * $signed(input_fmap_13[15:0]) +
	( 15'sd 9446) * $signed(input_fmap_14[15:0]) +
	( 16'sd 30952) * $signed(input_fmap_15[15:0]) +
	( 16'sd 31462) * $signed(input_fmap_16[15:0]) +
	( 16'sd 16760) * $signed(input_fmap_17[15:0]) +
	( 15'sd 10146) * $signed(input_fmap_18[15:0]) +
	( 15'sd 10110) * $signed(input_fmap_19[15:0]) +
	( 16'sd 16926) * $signed(input_fmap_20[15:0]) +
	( 15'sd 11526) * $signed(input_fmap_21[15:0]) +
	( 16'sd 24661) * $signed(input_fmap_22[15:0]) +
	( 15'sd 10802) * $signed(input_fmap_23[15:0]) +
	( 15'sd 10183) * $signed(input_fmap_24[15:0]) +
	( 16'sd 20688) * $signed(input_fmap_25[15:0]) +
	( 16'sd 19114) * $signed(input_fmap_26[15:0]) +
	( 14'sd 4787) * $signed(input_fmap_27[15:0]) +
	( 16'sd 26497) * $signed(input_fmap_28[15:0]) +
	( 10'sd 308) * $signed(input_fmap_29[15:0]) +
	( 16'sd 20454) * $signed(input_fmap_30[15:0]) +
	( 16'sd 24258) * $signed(input_fmap_31[15:0]) +
	( 16'sd 22863) * $signed(input_fmap_32[15:0]) +
	( 13'sd 3122) * $signed(input_fmap_33[15:0]) +
	( 16'sd 20853) * $signed(input_fmap_34[15:0]) +
	( 14'sd 4119) * $signed(input_fmap_35[15:0]) +
	( 15'sd 14714) * $signed(input_fmap_36[15:0]) +
	( 15'sd 14338) * $signed(input_fmap_37[15:0]) +
	( 16'sd 16482) * $signed(input_fmap_38[15:0]) +
	( 15'sd 12900) * $signed(input_fmap_39[15:0]) +
	( 16'sd 22960) * $signed(input_fmap_40[15:0]) +
	( 12'sd 1639) * $signed(input_fmap_41[15:0]) +
	( 16'sd 21005) * $signed(input_fmap_42[15:0]) +
	( 14'sd 7838) * $signed(input_fmap_43[15:0]) +
	( 14'sd 4834) * $signed(input_fmap_44[15:0]) +
	( 15'sd 15062) * $signed(input_fmap_45[15:0]) +
	( 10'sd 481) * $signed(input_fmap_46[15:0]) +
	( 13'sd 3556) * $signed(input_fmap_47[15:0]) +
	( 15'sd 10263) * $signed(input_fmap_48[15:0]) +
	( 16'sd 28354) * $signed(input_fmap_49[15:0]) +
	( 14'sd 7290) * $signed(input_fmap_50[15:0]) +
	( 14'sd 6867) * $signed(input_fmap_51[15:0]) +
	( 15'sd 12241) * $signed(input_fmap_52[15:0]) +
	( 12'sd 1828) * $signed(input_fmap_53[15:0]) +
	( 16'sd 24554) * $signed(input_fmap_54[15:0]) +
	( 16'sd 23582) * $signed(input_fmap_55[15:0]) +
	( 14'sd 6783) * $signed(input_fmap_56[15:0]) +
	( 14'sd 7957) * $signed(input_fmap_57[15:0]) +
	( 16'sd 21362) * $signed(input_fmap_58[15:0]) +
	( 16'sd 20144) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1279) * $signed(input_fmap_60[15:0]) +
	( 16'sd 18694) * $signed(input_fmap_61[15:0]) +
	( 16'sd 18761) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20158) * $signed(input_fmap_63[15:0]) +
	( 7'sd 52) * $signed(input_fmap_64[15:0]) +
	( 15'sd 15194) * $signed(input_fmap_65[15:0]) +
	( 16'sd 31736) * $signed(input_fmap_66[15:0]) +
	( 16'sd 30655) * $signed(input_fmap_67[15:0]) +
	( 16'sd 25443) * $signed(input_fmap_68[15:0]) +
	( 15'sd 9731) * $signed(input_fmap_69[15:0]) +
	( 16'sd 24675) * $signed(input_fmap_70[15:0]) +
	( 16'sd 25534) * $signed(input_fmap_71[15:0]) +
	( 16'sd 17801) * $signed(input_fmap_72[15:0]) +
	( 15'sd 14996) * $signed(input_fmap_73[15:0]) +
	( 16'sd 19416) * $signed(input_fmap_74[15:0]) +
	( 16'sd 18002) * $signed(input_fmap_75[15:0]) +
	( 16'sd 26119) * $signed(input_fmap_76[15:0]) +
	( 16'sd 25589) * $signed(input_fmap_77[15:0]) +
	( 15'sd 11923) * $signed(input_fmap_78[15:0]) +
	( 15'sd 11342) * $signed(input_fmap_79[15:0]) +
	( 15'sd 14228) * $signed(input_fmap_80[15:0]) +
	( 16'sd 17213) * $signed(input_fmap_81[15:0]) +
	( 16'sd 21840) * $signed(input_fmap_82[15:0]) +
	( 16'sd 30809) * $signed(input_fmap_83[15:0]) +
	( 13'sd 2941) * $signed(input_fmap_84[15:0]) +
	( 14'sd 7258) * $signed(input_fmap_85[15:0]) +
	( 15'sd 9214) * $signed(input_fmap_86[15:0]) +
	( 13'sd 3208) * $signed(input_fmap_87[15:0]) +
	( 16'sd 27207) * $signed(input_fmap_88[15:0]) +
	( 14'sd 6867) * $signed(input_fmap_89[15:0]) +
	( 14'sd 4760) * $signed(input_fmap_90[15:0]) +
	( 12'sd 1621) * $signed(input_fmap_91[15:0]) +
	( 13'sd 3458) * $signed(input_fmap_92[15:0]) +
	( 16'sd 22035) * $signed(input_fmap_93[15:0]) +
	( 16'sd 28012) * $signed(input_fmap_94[15:0]) +
	( 16'sd 20359) * $signed(input_fmap_95[15:0]) +
	( 16'sd 21439) * $signed(input_fmap_96[15:0]) +
	( 16'sd 23645) * $signed(input_fmap_97[15:0]) +
	( 16'sd 28218) * $signed(input_fmap_98[15:0]) +
	( 16'sd 19908) * $signed(input_fmap_99[15:0]) +
	( 14'sd 7293) * $signed(input_fmap_100[15:0]) +
	( 13'sd 3501) * $signed(input_fmap_101[15:0]) +
	( 16'sd 23165) * $signed(input_fmap_102[15:0]) +
	( 12'sd 1107) * $signed(input_fmap_103[15:0]) +
	( 15'sd 12405) * $signed(input_fmap_104[15:0]) +
	( 15'sd 13344) * $signed(input_fmap_105[15:0]) +
	( 16'sd 26108) * $signed(input_fmap_106[15:0]) +
	( 15'sd 10128) * $signed(input_fmap_107[15:0]) +
	( 15'sd 10262) * $signed(input_fmap_108[15:0]) +
	( 15'sd 9641) * $signed(input_fmap_109[15:0]) +
	( 16'sd 25772) * $signed(input_fmap_110[15:0]) +
	( 16'sd 21069) * $signed(input_fmap_111[15:0]) +
	( 14'sd 5979) * $signed(input_fmap_112[15:0]) +
	( 16'sd 21267) * $signed(input_fmap_113[15:0]) +
	( 16'sd 31245) * $signed(input_fmap_114[15:0]) +
	( 14'sd 7057) * $signed(input_fmap_115[15:0]) +
	( 16'sd 24562) * $signed(input_fmap_116[15:0]) +
	( 16'sd 24778) * $signed(input_fmap_117[15:0]) +
	( 15'sd 9398) * $signed(input_fmap_118[15:0]) +
	( 14'sd 6798) * $signed(input_fmap_119[15:0]) +
	( 15'sd 15788) * $signed(input_fmap_120[15:0]) +
	( 13'sd 2233) * $signed(input_fmap_121[15:0]) +
	( 14'sd 4921) * $signed(input_fmap_122[15:0]) +
	( 15'sd 10051) * $signed(input_fmap_123[15:0]) +
	( 16'sd 24976) * $signed(input_fmap_124[15:0]) +
	( 15'sd 11157) * $signed(input_fmap_125[15:0]) +
	( 14'sd 4247) * $signed(input_fmap_126[15:0]) +
	( 13'sd 2277) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 9'sd 155) * $signed(input_fmap_0[15:0]) +
	( 16'sd 25769) * $signed(input_fmap_1[15:0]) +
	( 16'sd 21971) * $signed(input_fmap_2[15:0]) +
	( 16'sd 28167) * $signed(input_fmap_3[15:0]) +
	( 15'sd 12291) * $signed(input_fmap_4[15:0]) +
	( 12'sd 1623) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2717) * $signed(input_fmap_6[15:0]) +
	( 16'sd 25052) * $signed(input_fmap_7[15:0]) +
	( 16'sd 18480) * $signed(input_fmap_8[15:0]) +
	( 15'sd 10227) * $signed(input_fmap_9[15:0]) +
	( 13'sd 3092) * $signed(input_fmap_10[15:0]) +
	( 14'sd 7001) * $signed(input_fmap_11[15:0]) +
	( 16'sd 27022) * $signed(input_fmap_12[15:0]) +
	( 15'sd 15621) * $signed(input_fmap_13[15:0]) +
	( 16'sd 20596) * $signed(input_fmap_14[15:0]) +
	( 16'sd 22750) * $signed(input_fmap_15[15:0]) +
	( 11'sd 856) * $signed(input_fmap_16[15:0]) +
	( 16'sd 30003) * $signed(input_fmap_17[15:0]) +
	( 16'sd 25792) * $signed(input_fmap_18[15:0]) +
	( 16'sd 28677) * $signed(input_fmap_19[15:0]) +
	( 15'sd 15458) * $signed(input_fmap_20[15:0]) +
	( 16'sd 20568) * $signed(input_fmap_21[15:0]) +
	( 15'sd 14698) * $signed(input_fmap_22[15:0]) +
	( 13'sd 3239) * $signed(input_fmap_23[15:0]) +
	( 16'sd 26514) * $signed(input_fmap_24[15:0]) +
	( 13'sd 3766) * $signed(input_fmap_25[15:0]) +
	( 14'sd 4543) * $signed(input_fmap_26[15:0]) +
	( 16'sd 21974) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24223) * $signed(input_fmap_28[15:0]) +
	( 14'sd 4322) * $signed(input_fmap_29[15:0]) +
	( 16'sd 17278) * $signed(input_fmap_30[15:0]) +
	( 16'sd 16821) * $signed(input_fmap_31[15:0]) +
	( 15'sd 11949) * $signed(input_fmap_32[15:0]) +
	( 11'sd 655) * $signed(input_fmap_33[15:0]) +
	( 14'sd 4873) * $signed(input_fmap_34[15:0]) +
	( 16'sd 32182) * $signed(input_fmap_35[15:0]) +
	( 16'sd 32650) * $signed(input_fmap_36[15:0]) +
	( 16'sd 24052) * $signed(input_fmap_37[15:0]) +
	( 15'sd 9008) * $signed(input_fmap_38[15:0]) +
	( 15'sd 13734) * $signed(input_fmap_39[15:0]) +
	( 16'sd 16706) * $signed(input_fmap_40[15:0]) +
	( 15'sd 14112) * $signed(input_fmap_41[15:0]) +
	( 16'sd 23791) * $signed(input_fmap_42[15:0]) +
	( 16'sd 23932) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31924) * $signed(input_fmap_44[15:0]) +
	( 16'sd 26142) * $signed(input_fmap_45[15:0]) +
	( 16'sd 21491) * $signed(input_fmap_46[15:0]) +
	( 16'sd 26243) * $signed(input_fmap_47[15:0]) +
	( 16'sd 25029) * $signed(input_fmap_48[15:0]) +
	( 16'sd 18592) * $signed(input_fmap_49[15:0]) +
	( 14'sd 6988) * $signed(input_fmap_50[15:0]) +
	( 14'sd 8119) * $signed(input_fmap_51[15:0]) +
	( 16'sd 28678) * $signed(input_fmap_52[15:0]) +
	( 16'sd 26402) * $signed(input_fmap_53[15:0]) +
	( 13'sd 2795) * $signed(input_fmap_54[15:0]) +
	( 16'sd 27072) * $signed(input_fmap_55[15:0]) +
	( 15'sd 16069) * $signed(input_fmap_56[15:0]) +
	( 15'sd 11715) * $signed(input_fmap_57[15:0]) +
	( 14'sd 4720) * $signed(input_fmap_58[15:0]) +
	( 16'sd 22091) * $signed(input_fmap_59[15:0]) +
	( 15'sd 15260) * $signed(input_fmap_60[15:0]) +
	( 16'sd 23729) * $signed(input_fmap_61[15:0]) +
	( 14'sd 4972) * $signed(input_fmap_62[15:0]) +
	( 15'sd 14183) * $signed(input_fmap_63[15:0]) +
	( 16'sd 32642) * $signed(input_fmap_64[15:0]) +
	( 16'sd 30186) * $signed(input_fmap_65[15:0]) +
	( 14'sd 8095) * $signed(input_fmap_66[15:0]) +
	( 16'sd 32257) * $signed(input_fmap_67[15:0]) +
	( 16'sd 19961) * $signed(input_fmap_68[15:0]) +
	( 16'sd 19888) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31492) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31283) * $signed(input_fmap_71[15:0]) +
	( 10'sd 360) * $signed(input_fmap_72[15:0]) +
	( 16'sd 16441) * $signed(input_fmap_73[15:0]) +
	( 15'sd 9936) * $signed(input_fmap_74[15:0]) +
	( 15'sd 16297) * $signed(input_fmap_75[15:0]) +
	( 15'sd 8600) * $signed(input_fmap_76[15:0]) +
	( 16'sd 25541) * $signed(input_fmap_77[15:0]) +
	( 16'sd 29138) * $signed(input_fmap_78[15:0]) +
	( 12'sd 1102) * $signed(input_fmap_79[15:0]) +
	( 16'sd 29242) * $signed(input_fmap_80[15:0]) +
	( 15'sd 15596) * $signed(input_fmap_81[15:0]) +
	( 15'sd 15601) * $signed(input_fmap_82[15:0]) +
	( 14'sd 8164) * $signed(input_fmap_83[15:0]) +
	( 16'sd 29951) * $signed(input_fmap_84[15:0]) +
	( 15'sd 11283) * $signed(input_fmap_85[15:0]) +
	( 11'sd 961) * $signed(input_fmap_86[15:0]) +
	( 15'sd 11124) * $signed(input_fmap_87[15:0]) +
	( 16'sd 20797) * $signed(input_fmap_88[15:0]) +
	( 15'sd 8804) * $signed(input_fmap_89[15:0]) +
	( 15'sd 13397) * $signed(input_fmap_90[15:0]) +
	( 16'sd 24559) * $signed(input_fmap_91[15:0]) +
	( 16'sd 28198) * $signed(input_fmap_92[15:0]) +
	( 16'sd 31523) * $signed(input_fmap_93[15:0]) +
	( 13'sd 4028) * $signed(input_fmap_94[15:0]) +
	( 15'sd 15490) * $signed(input_fmap_95[15:0]) +
	( 15'sd 11883) * $signed(input_fmap_96[15:0]) +
	( 16'sd 26461) * $signed(input_fmap_97[15:0]) +
	( 15'sd 9206) * $signed(input_fmap_98[15:0]) +
	( 14'sd 5872) * $signed(input_fmap_99[15:0]) +
	( 14'sd 4505) * $signed(input_fmap_100[15:0]) +
	( 15'sd 13667) * $signed(input_fmap_101[15:0]) +
	( 15'sd 15128) * $signed(input_fmap_102[15:0]) +
	( 13'sd 2673) * $signed(input_fmap_103[15:0]) +
	( 16'sd 19294) * $signed(input_fmap_104[15:0]) +
	( 16'sd 29785) * $signed(input_fmap_105[15:0]) +
	( 12'sd 1324) * $signed(input_fmap_106[15:0]) +
	( 15'sd 14179) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15698) * $signed(input_fmap_108[15:0]) +
	( 16'sd 29299) * $signed(input_fmap_109[15:0]) +
	( 15'sd 11504) * $signed(input_fmap_110[15:0]) +
	( 16'sd 26810) * $signed(input_fmap_111[15:0]) +
	( 15'sd 16009) * $signed(input_fmap_112[15:0]) +
	( 16'sd 31059) * $signed(input_fmap_113[15:0]) +
	( 15'sd 8715) * $signed(input_fmap_114[15:0]) +
	( 16'sd 30530) * $signed(input_fmap_115[15:0]) +
	( 16'sd 23068) * $signed(input_fmap_116[15:0]) +
	( 16'sd 18677) * $signed(input_fmap_117[15:0]) +
	( 16'sd 18591) * $signed(input_fmap_118[15:0]) +
	( 15'sd 10209) * $signed(input_fmap_119[15:0]) +
	( 16'sd 22957) * $signed(input_fmap_120[15:0]) +
	( 11'sd 535) * $signed(input_fmap_121[15:0]) +
	( 16'sd 25554) * $signed(input_fmap_122[15:0]) +
	( 14'sd 5076) * $signed(input_fmap_123[15:0]) +
	( 14'sd 5017) * $signed(input_fmap_124[15:0]) +
	( 16'sd 21014) * $signed(input_fmap_125[15:0]) +
	( 14'sd 7688) * $signed(input_fmap_126[15:0]) +
	( 15'sd 14261) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 14'sd 5889) * $signed(input_fmap_0[15:0]) +
	( 16'sd 30896) * $signed(input_fmap_1[15:0]) +
	( 14'sd 7078) * $signed(input_fmap_2[15:0]) +
	( 15'sd 12379) * $signed(input_fmap_3[15:0]) +
	( 16'sd 26557) * $signed(input_fmap_4[15:0]) +
	( 15'sd 14540) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2653) * $signed(input_fmap_6[15:0]) +
	( 10'sd 436) * $signed(input_fmap_7[15:0]) +
	( 16'sd 29765) * $signed(input_fmap_8[15:0]) +
	( 15'sd 9935) * $signed(input_fmap_9[15:0]) +
	( 16'sd 29144) * $signed(input_fmap_10[15:0]) +
	( 16'sd 24661) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20222) * $signed(input_fmap_12[15:0]) +
	( 12'sd 1707) * $signed(input_fmap_13[15:0]) +
	( 15'sd 10243) * $signed(input_fmap_14[15:0]) +
	( 15'sd 10206) * $signed(input_fmap_15[15:0]) +
	( 16'sd 27771) * $signed(input_fmap_16[15:0]) +
	( 16'sd 27823) * $signed(input_fmap_17[15:0]) +
	( 16'sd 22143) * $signed(input_fmap_18[15:0]) +
	( 16'sd 20402) * $signed(input_fmap_19[15:0]) +
	( 16'sd 23361) * $signed(input_fmap_20[15:0]) +
	( 15'sd 15091) * $signed(input_fmap_21[15:0]) +
	( 16'sd 18427) * $signed(input_fmap_22[15:0]) +
	( 16'sd 17661) * $signed(input_fmap_23[15:0]) +
	( 10'sd 405) * $signed(input_fmap_24[15:0]) +
	( 13'sd 2736) * $signed(input_fmap_25[15:0]) +
	( 16'sd 18965) * $signed(input_fmap_26[15:0]) +
	( 16'sd 22621) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24870) * $signed(input_fmap_28[15:0]) +
	( 16'sd 20890) * $signed(input_fmap_29[15:0]) +
	( 12'sd 1257) * $signed(input_fmap_30[15:0]) +
	( 16'sd 28835) * $signed(input_fmap_31[15:0]) +
	( 14'sd 7368) * $signed(input_fmap_32[15:0]) +
	( 16'sd 27058) * $signed(input_fmap_33[15:0]) +
	( 16'sd 32583) * $signed(input_fmap_34[15:0]) +
	( 16'sd 27617) * $signed(input_fmap_35[15:0]) +
	( 15'sd 9783) * $signed(input_fmap_36[15:0]) +
	( 13'sd 3187) * $signed(input_fmap_37[15:0]) +
	( 16'sd 20049) * $signed(input_fmap_38[15:0]) +
	( 14'sd 6397) * $signed(input_fmap_39[15:0]) +
	( 16'sd 17970) * $signed(input_fmap_40[15:0]) +
	( 14'sd 6920) * $signed(input_fmap_41[15:0]) +
	( 16'sd 28505) * $signed(input_fmap_42[15:0]) +
	( 14'sd 7759) * $signed(input_fmap_43[15:0]) +
	( 16'sd 22133) * $signed(input_fmap_44[15:0]) +
	( 16'sd 32245) * $signed(input_fmap_45[15:0]) +
	( 16'sd 30541) * $signed(input_fmap_46[15:0]) +
	( 16'sd 17601) * $signed(input_fmap_47[15:0]) +
	( 16'sd 17785) * $signed(input_fmap_48[15:0]) +
	( 16'sd 19261) * $signed(input_fmap_49[15:0]) +
	( 15'sd 15098) * $signed(input_fmap_50[15:0]) +
	( 16'sd 23711) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19439) * $signed(input_fmap_52[15:0]) +
	( 16'sd 17843) * $signed(input_fmap_53[15:0]) +
	( 16'sd 18679) * $signed(input_fmap_54[15:0]) +
	( 12'sd 1853) * $signed(input_fmap_55[15:0]) +
	( 16'sd 18496) * $signed(input_fmap_56[15:0]) +
	( 14'sd 6910) * $signed(input_fmap_57[15:0]) +
	( 13'sd 2091) * $signed(input_fmap_58[15:0]) +
	( 16'sd 24650) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1568) * $signed(input_fmap_60[15:0]) +
	( 16'sd 31513) * $signed(input_fmap_61[15:0]) +
	( 16'sd 22893) * $signed(input_fmap_62[15:0]) +
	( 16'sd 23235) * $signed(input_fmap_63[15:0]) +
	( 16'sd 27954) * $signed(input_fmap_64[15:0]) +
	( 16'sd 18813) * $signed(input_fmap_65[15:0]) +
	( 16'sd 23569) * $signed(input_fmap_66[15:0]) +
	( 16'sd 22263) * $signed(input_fmap_67[15:0]) +
	( 14'sd 5947) * $signed(input_fmap_68[15:0]) +
	( 14'sd 8152) * $signed(input_fmap_69[15:0]) +
	( 15'sd 14502) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11923) * $signed(input_fmap_71[15:0]) +
	( 16'sd 31875) * $signed(input_fmap_72[15:0]) +
	( 15'sd 14327) * $signed(input_fmap_73[15:0]) +
	( 16'sd 26524) * $signed(input_fmap_74[15:0]) +
	( 13'sd 2561) * $signed(input_fmap_75[15:0]) +
	( 9'sd 157) * $signed(input_fmap_76[15:0]) +
	( 15'sd 9233) * $signed(input_fmap_77[15:0]) +
	( 13'sd 3848) * $signed(input_fmap_78[15:0]) +
	( 16'sd 26976) * $signed(input_fmap_79[15:0]) +
	( 16'sd 19821) * $signed(input_fmap_80[15:0]) +
	( 13'sd 3876) * $signed(input_fmap_81[15:0]) +
	( 14'sd 4757) * $signed(input_fmap_82[15:0]) +
	( 16'sd 32104) * $signed(input_fmap_83[15:0]) +
	( 14'sd 5551) * $signed(input_fmap_84[15:0]) +
	( 16'sd 25821) * $signed(input_fmap_85[15:0]) +
	( 16'sd 20945) * $signed(input_fmap_86[15:0]) +
	( 15'sd 12740) * $signed(input_fmap_87[15:0]) +
	( 15'sd 16167) * $signed(input_fmap_88[15:0]) +
	( 16'sd 23042) * $signed(input_fmap_89[15:0]) +
	( 15'sd 13729) * $signed(input_fmap_90[15:0]) +
	( 16'sd 29155) * $signed(input_fmap_91[15:0]) +
	( 15'sd 15583) * $signed(input_fmap_92[15:0]) +
	( 14'sd 4711) * $signed(input_fmap_93[15:0]) +
	( 16'sd 21384) * $signed(input_fmap_94[15:0]) +
	( 15'sd 11239) * $signed(input_fmap_95[15:0]) +
	( 14'sd 6211) * $signed(input_fmap_96[15:0]) +
	( 13'sd 3554) * $signed(input_fmap_97[15:0]) +
	( 15'sd 12751) * $signed(input_fmap_98[15:0]) +
	( 11'sd 598) * $signed(input_fmap_99[15:0]) +
	( 16'sd 17052) * $signed(input_fmap_100[15:0]) +
	( 10'sd 343) * $signed(input_fmap_101[15:0]) +
	( 16'sd 16832) * $signed(input_fmap_102[15:0]) +
	( 16'sd 20692) * $signed(input_fmap_103[15:0]) +
	( 11'sd 876) * $signed(input_fmap_104[15:0]) +
	( 15'sd 13620) * $signed(input_fmap_105[15:0]) +
	( 16'sd 18546) * $signed(input_fmap_106[15:0]) +
	( 15'sd 16286) * $signed(input_fmap_107[15:0]) +
	( 16'sd 16869) * $signed(input_fmap_108[15:0]) +
	( 15'sd 11703) * $signed(input_fmap_109[15:0]) +
	( 14'sd 4824) * $signed(input_fmap_110[15:0]) +
	( 16'sd 23298) * $signed(input_fmap_111[15:0]) +
	( 16'sd 28314) * $signed(input_fmap_112[15:0]) +
	( 16'sd 27772) * $signed(input_fmap_113[15:0]) +
	( 14'sd 5814) * $signed(input_fmap_114[15:0]) +
	( 14'sd 4766) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15082) * $signed(input_fmap_116[15:0]) +
	( 16'sd 18658) * $signed(input_fmap_117[15:0]) +
	( 16'sd 30425) * $signed(input_fmap_118[15:0]) +
	( 16'sd 18652) * $signed(input_fmap_119[15:0]) +
	( 13'sd 2833) * $signed(input_fmap_120[15:0]) +
	( 16'sd 23678) * $signed(input_fmap_121[15:0]) +
	( 16'sd 18149) * $signed(input_fmap_122[15:0]) +
	( 15'sd 11961) * $signed(input_fmap_123[15:0]) +
	( 13'sd 2655) * $signed(input_fmap_124[15:0]) +
	( 12'sd 1538) * $signed(input_fmap_125[15:0]) +
	( 16'sd 18024) * $signed(input_fmap_126[15:0]) +
	( 14'sd 6856) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 16'sd 21840) * $signed(input_fmap_0[15:0]) +
	( 13'sd 3511) * $signed(input_fmap_1[15:0]) +
	( 15'sd 12375) * $signed(input_fmap_2[15:0]) +
	( 16'sd 29088) * $signed(input_fmap_3[15:0]) +
	( 14'sd 5500) * $signed(input_fmap_4[15:0]) +
	( 16'sd 21337) * $signed(input_fmap_5[15:0]) +
	( 16'sd 22563) * $signed(input_fmap_6[15:0]) +
	( 16'sd 18598) * $signed(input_fmap_7[15:0]) +
	( 16'sd 28235) * $signed(input_fmap_8[15:0]) +
	( 16'sd 22236) * $signed(input_fmap_9[15:0]) +
	( 16'sd 22337) * $signed(input_fmap_10[15:0]) +
	( 16'sd 29048) * $signed(input_fmap_11[15:0]) +
	( 16'sd 31867) * $signed(input_fmap_12[15:0]) +
	( 16'sd 23195) * $signed(input_fmap_13[15:0]) +
	( 16'sd 20970) * $signed(input_fmap_14[15:0]) +
	( 10'sd 367) * $signed(input_fmap_15[15:0]) +
	( 14'sd 6090) * $signed(input_fmap_16[15:0]) +
	( 15'sd 8754) * $signed(input_fmap_17[15:0]) +
	( 15'sd 8318) * $signed(input_fmap_18[15:0]) +
	( 16'sd 20226) * $signed(input_fmap_19[15:0]) +
	( 16'sd 29751) * $signed(input_fmap_20[15:0]) +
	( 16'sd 32551) * $signed(input_fmap_21[15:0]) +
	( 16'sd 21008) * $signed(input_fmap_22[15:0]) +
	( 15'sd 16013) * $signed(input_fmap_23[15:0]) +
	( 15'sd 11557) * $signed(input_fmap_24[15:0]) +
	( 16'sd 24698) * $signed(input_fmap_25[15:0]) +
	( 15'sd 9734) * $signed(input_fmap_26[15:0]) +
	( 16'sd 22200) * $signed(input_fmap_27[15:0]) +
	( 15'sd 12491) * $signed(input_fmap_28[15:0]) +
	( 16'sd 16735) * $signed(input_fmap_29[15:0]) +
	( 15'sd 13020) * $signed(input_fmap_30[15:0]) +
	( 16'sd 23082) * $signed(input_fmap_31[15:0]) +
	( 14'sd 7178) * $signed(input_fmap_32[15:0]) +
	( 15'sd 15740) * $signed(input_fmap_33[15:0]) +
	( 15'sd 14567) * $signed(input_fmap_34[15:0]) +
	( 14'sd 5203) * $signed(input_fmap_35[15:0]) +
	( 16'sd 17917) * $signed(input_fmap_36[15:0]) +
	( 15'sd 9531) * $signed(input_fmap_37[15:0]) +
	( 16'sd 16895) * $signed(input_fmap_38[15:0]) +
	( 14'sd 8107) * $signed(input_fmap_39[15:0]) +
	( 14'sd 7232) * $signed(input_fmap_40[15:0]) +
	( 14'sd 7449) * $signed(input_fmap_41[15:0]) +
	( 14'sd 4114) * $signed(input_fmap_42[15:0]) +
	( 14'sd 6620) * $signed(input_fmap_43[15:0]) +
	( 15'sd 13317) * $signed(input_fmap_44[15:0]) +
	( 16'sd 24769) * $signed(input_fmap_45[15:0]) +
	( 16'sd 21234) * $signed(input_fmap_46[15:0]) +
	( 15'sd 13066) * $signed(input_fmap_47[15:0]) +
	( 16'sd 16619) * $signed(input_fmap_48[15:0]) +
	( 9'sd 238) * $signed(input_fmap_49[15:0]) +
	( 16'sd 21417) * $signed(input_fmap_50[15:0]) +
	( 16'sd 31576) * $signed(input_fmap_51[15:0]) +
	( 15'sd 12645) * $signed(input_fmap_52[15:0]) +
	( 16'sd 26986) * $signed(input_fmap_53[15:0]) +
	( 16'sd 21334) * $signed(input_fmap_54[15:0]) +
	( 14'sd 5664) * $signed(input_fmap_55[15:0]) +
	( 16'sd 23690) * $signed(input_fmap_56[15:0]) +
	( 16'sd 23296) * $signed(input_fmap_57[15:0]) +
	( 15'sd 10120) * $signed(input_fmap_58[15:0]) +
	( 15'sd 8789) * $signed(input_fmap_59[15:0]) +
	( 11'sd 909) * $signed(input_fmap_60[15:0]) +
	( 14'sd 4878) * $signed(input_fmap_61[15:0]) +
	( 16'sd 18569) * $signed(input_fmap_62[15:0]) +
	( 14'sd 4479) * $signed(input_fmap_63[15:0]) +
	( 13'sd 3789) * $signed(input_fmap_64[15:0]) +
	( 15'sd 9906) * $signed(input_fmap_65[15:0]) +
	( 16'sd 16979) * $signed(input_fmap_66[15:0]) +
	( 16'sd 23245) * $signed(input_fmap_67[15:0]) +
	( 16'sd 22306) * $signed(input_fmap_68[15:0]) +
	( 16'sd 29732) * $signed(input_fmap_69[15:0]) +
	( 16'sd 19877) * $signed(input_fmap_70[15:0]) +
	( 15'sd 12948) * $signed(input_fmap_71[15:0]) +
	( 14'sd 7066) * $signed(input_fmap_72[15:0]) +
	( 16'sd 26457) * $signed(input_fmap_73[15:0]) +
	( 16'sd 31882) * $signed(input_fmap_74[15:0]) +
	( 15'sd 15771) * $signed(input_fmap_75[15:0]) +
	( 16'sd 18029) * $signed(input_fmap_76[15:0]) +
	( 16'sd 20236) * $signed(input_fmap_77[15:0]) +
	( 16'sd 32300) * $signed(input_fmap_78[15:0]) +
	( 16'sd 29303) * $signed(input_fmap_79[15:0]) +
	( 15'sd 9817) * $signed(input_fmap_80[15:0]) +
	( 16'sd 20996) * $signed(input_fmap_81[15:0]) +
	( 14'sd 5924) * $signed(input_fmap_82[15:0]) +
	( 13'sd 3998) * $signed(input_fmap_83[15:0]) +
	( 16'sd 27607) * $signed(input_fmap_84[15:0]) +
	( 16'sd 23817) * $signed(input_fmap_85[15:0]) +
	( 16'sd 24677) * $signed(input_fmap_86[15:0]) +
	( 16'sd 17461) * $signed(input_fmap_87[15:0]) +
	( 16'sd 20912) * $signed(input_fmap_88[15:0]) +
	( 14'sd 4106) * $signed(input_fmap_89[15:0]) +
	( 16'sd 21280) * $signed(input_fmap_90[15:0]) +
	( 16'sd 31798) * $signed(input_fmap_91[15:0]) +
	( 15'sd 14449) * $signed(input_fmap_92[15:0]) +
	( 16'sd 26177) * $signed(input_fmap_93[15:0]) +
	( 15'sd 9003) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25217) * $signed(input_fmap_95[15:0]) +
	( 13'sd 3341) * $signed(input_fmap_96[15:0]) +
	( 15'sd 10964) * $signed(input_fmap_97[15:0]) +
	( 15'sd 8357) * $signed(input_fmap_98[15:0]) +
	( 16'sd 24908) * $signed(input_fmap_99[15:0]) +
	( 16'sd 28956) * $signed(input_fmap_100[15:0]) +
	( 13'sd 2159) * $signed(input_fmap_101[15:0]) +
	( 14'sd 4984) * $signed(input_fmap_102[15:0]) +
	( 14'sd 7860) * $signed(input_fmap_103[15:0]) +
	( 16'sd 20086) * $signed(input_fmap_104[15:0]) +
	( 15'sd 9878) * $signed(input_fmap_105[15:0]) +
	( 15'sd 13558) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27025) * $signed(input_fmap_107[15:0]) +
	( 16'sd 28663) * $signed(input_fmap_108[15:0]) +
	( 15'sd 11015) * $signed(input_fmap_109[15:0]) +
	( 15'sd 11611) * $signed(input_fmap_110[15:0]) +
	( 15'sd 12407) * $signed(input_fmap_111[15:0]) +
	( 14'sd 6116) * $signed(input_fmap_112[15:0]) +
	( 14'sd 7116) * $signed(input_fmap_113[15:0]) +
	( 15'sd 13684) * $signed(input_fmap_114[15:0]) +
	( 16'sd 23032) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15247) * $signed(input_fmap_116[15:0]) +
	( 14'sd 8098) * $signed(input_fmap_117[15:0]) +
	( 16'sd 17807) * $signed(input_fmap_118[15:0]) +
	( 15'sd 10075) * $signed(input_fmap_119[15:0]) +
	( 16'sd 31257) * $signed(input_fmap_120[15:0]) +
	( 13'sd 2889) * $signed(input_fmap_121[15:0]) +
	( 14'sd 5817) * $signed(input_fmap_122[15:0]) +
	( 16'sd 23529) * $signed(input_fmap_123[15:0]) +
	( 14'sd 5338) * $signed(input_fmap_124[15:0]) +
	( 16'sd 27263) * $signed(input_fmap_125[15:0]) +
	( 15'sd 12760) * $signed(input_fmap_126[15:0]) +
	( 16'sd 21014) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 15'sd 14000) * $signed(input_fmap_0[15:0]) +
	( 16'sd 25315) * $signed(input_fmap_1[15:0]) +
	( 16'sd 21505) * $signed(input_fmap_2[15:0]) +
	( 16'sd 32682) * $signed(input_fmap_3[15:0]) +
	( 16'sd 27193) * $signed(input_fmap_4[15:0]) +
	( 16'sd 24302) * $signed(input_fmap_5[15:0]) +
	( 16'sd 23109) * $signed(input_fmap_6[15:0]) +
	( 12'sd 1571) * $signed(input_fmap_7[15:0]) +
	( 16'sd 19620) * $signed(input_fmap_8[15:0]) +
	( 14'sd 7107) * $signed(input_fmap_9[15:0]) +
	( 16'sd 25890) * $signed(input_fmap_10[15:0]) +
	( 16'sd 25455) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20458) * $signed(input_fmap_12[15:0]) +
	( 16'sd 18763) * $signed(input_fmap_13[15:0]) +
	( 13'sd 2617) * $signed(input_fmap_14[15:0]) +
	( 15'sd 12475) * $signed(input_fmap_15[15:0]) +
	( 16'sd 18714) * $signed(input_fmap_16[15:0]) +
	( 16'sd 23990) * $signed(input_fmap_17[15:0]) +
	( 14'sd 6564) * $signed(input_fmap_18[15:0]) +
	( 13'sd 3141) * $signed(input_fmap_19[15:0]) +
	( 16'sd 25824) * $signed(input_fmap_20[15:0]) +
	( 16'sd 24516) * $signed(input_fmap_21[15:0]) +
	( 14'sd 4429) * $signed(input_fmap_22[15:0]) +
	( 15'sd 10324) * $signed(input_fmap_23[15:0]) +
	( 13'sd 2631) * $signed(input_fmap_24[15:0]) +
	( 16'sd 19420) * $signed(input_fmap_25[15:0]) +
	( 16'sd 23901) * $signed(input_fmap_26[15:0]) +
	( 16'sd 30330) * $signed(input_fmap_27[15:0]) +
	( 15'sd 12654) * $signed(input_fmap_28[15:0]) +
	( 16'sd 18171) * $signed(input_fmap_29[15:0]) +
	( 15'sd 15309) * $signed(input_fmap_30[15:0]) +
	( 15'sd 8260) * $signed(input_fmap_31[15:0]) +
	( 16'sd 25247) * $signed(input_fmap_32[15:0]) +
	( 16'sd 27506) * $signed(input_fmap_33[15:0]) +
	( 16'sd 25879) * $signed(input_fmap_34[15:0]) +
	( 16'sd 17536) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2254) * $signed(input_fmap_36[15:0]) +
	( 16'sd 19655) * $signed(input_fmap_37[15:0]) +
	( 16'sd 30823) * $signed(input_fmap_38[15:0]) +
	( 14'sd 7336) * $signed(input_fmap_39[15:0]) +
	( 14'sd 7509) * $signed(input_fmap_40[15:0]) +
	( 15'sd 9013) * $signed(input_fmap_41[15:0]) +
	( 15'sd 9673) * $signed(input_fmap_42[15:0]) +
	( 12'sd 1716) * $signed(input_fmap_43[15:0]) +
	( 16'sd 24078) * $signed(input_fmap_44[15:0]) +
	( 16'sd 22118) * $signed(input_fmap_45[15:0]) +
	( 15'sd 11302) * $signed(input_fmap_46[15:0]) +
	( 15'sd 8427) * $signed(input_fmap_47[15:0]) +
	( 14'sd 7982) * $signed(input_fmap_48[15:0]) +
	( 11'sd 1011) * $signed(input_fmap_49[15:0]) +
	( 16'sd 20334) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15997) * $signed(input_fmap_51[15:0]) +
	( 16'sd 17644) * $signed(input_fmap_52[15:0]) +
	( 16'sd 29502) * $signed(input_fmap_53[15:0]) +
	( 15'sd 16288) * $signed(input_fmap_54[15:0]) +
	( 16'sd 23260) * $signed(input_fmap_55[15:0]) +
	( 16'sd 30629) * $signed(input_fmap_56[15:0]) +
	( 13'sd 3097) * $signed(input_fmap_57[15:0]) +
	( 16'sd 26784) * $signed(input_fmap_58[15:0]) +
	( 16'sd 26499) * $signed(input_fmap_59[15:0]) +
	( 15'sd 8522) * $signed(input_fmap_60[15:0]) +
	( 16'sd 28123) * $signed(input_fmap_61[15:0]) +
	( 16'sd 25853) * $signed(input_fmap_62[15:0]) +
	( 16'sd 17970) * $signed(input_fmap_63[15:0]) +
	( 16'sd 31133) * $signed(input_fmap_64[15:0]) +
	( 16'sd 26439) * $signed(input_fmap_65[15:0]) +
	( 16'sd 17537) * $signed(input_fmap_66[15:0]) +
	( 15'sd 12361) * $signed(input_fmap_67[15:0]) +
	( 15'sd 14463) * $signed(input_fmap_68[15:0]) +
	( 16'sd 24819) * $signed(input_fmap_69[15:0]) +
	( 14'sd 5279) * $signed(input_fmap_70[15:0]) +
	( 16'sd 25129) * $signed(input_fmap_71[15:0]) +
	( 14'sd 7630) * $signed(input_fmap_72[15:0]) +
	( 15'sd 14353) * $signed(input_fmap_73[15:0]) +
	( 16'sd 23463) * $signed(input_fmap_74[15:0]) +
	( 16'sd 24688) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19363) * $signed(input_fmap_76[15:0]) +
	( 13'sd 2181) * $signed(input_fmap_77[15:0]) +
	( 16'sd 31998) * $signed(input_fmap_78[15:0]) +
	( 16'sd 21061) * $signed(input_fmap_79[15:0]) +
	( 16'sd 27371) * $signed(input_fmap_80[15:0]) +
	( 16'sd 31061) * $signed(input_fmap_81[15:0]) +
	( 11'sd 671) * $signed(input_fmap_82[15:0]) +
	( 15'sd 16309) * $signed(input_fmap_83[15:0]) +
	( 16'sd 21070) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24038) * $signed(input_fmap_85[15:0]) +
	( 12'sd 1725) * $signed(input_fmap_86[15:0]) +
	( 13'sd 2954) * $signed(input_fmap_87[15:0]) +
	( 15'sd 15940) * $signed(input_fmap_88[15:0]) +
	( 16'sd 26483) * $signed(input_fmap_89[15:0]) +
	( 15'sd 9848) * $signed(input_fmap_90[15:0]) +
	( 16'sd 25452) * $signed(input_fmap_91[15:0]) +
	( 15'sd 8734) * $signed(input_fmap_92[15:0]) +
	( 16'sd 25347) * $signed(input_fmap_93[15:0]) +
	( 16'sd 18471) * $signed(input_fmap_94[15:0]) +
	( 16'sd 23968) * $signed(input_fmap_95[15:0]) +
	( 15'sd 13863) * $signed(input_fmap_96[15:0]) +
	( 11'sd 696) * $signed(input_fmap_97[15:0]) +
	( 16'sd 19443) * $signed(input_fmap_98[15:0]) +
	( 14'sd 7555) * $signed(input_fmap_99[15:0]) +
	( 16'sd 20673) * $signed(input_fmap_100[15:0]) +
	( 15'sd 12982) * $signed(input_fmap_101[15:0]) +
	( 16'sd 31142) * $signed(input_fmap_102[15:0]) +
	( 16'sd 18023) * $signed(input_fmap_103[15:0]) +
	( 15'sd 12588) * $signed(input_fmap_104[15:0]) +
	( 14'sd 5218) * $signed(input_fmap_105[15:0]) +
	( 16'sd 26647) * $signed(input_fmap_106[15:0]) +
	( 16'sd 17151) * $signed(input_fmap_107[15:0]) +
	( 16'sd 18816) * $signed(input_fmap_108[15:0]) +
	( 13'sd 2445) * $signed(input_fmap_109[15:0]) +
	( 14'sd 7698) * $signed(input_fmap_110[15:0]) +
	( 14'sd 7241) * $signed(input_fmap_111[15:0]) +
	( 15'sd 13720) * $signed(input_fmap_112[15:0]) +
	( 16'sd 22616) * $signed(input_fmap_113[15:0]) +
	( 15'sd 8716) * $signed(input_fmap_114[15:0]) +
	( 16'sd 17386) * $signed(input_fmap_115[15:0]) +
	( 16'sd 16933) * $signed(input_fmap_116[15:0]) +
	( 13'sd 3597) * $signed(input_fmap_117[15:0]) +
	( 14'sd 4594) * $signed(input_fmap_118[15:0]) +
	( 16'sd 25875) * $signed(input_fmap_119[15:0]) +
	( 15'sd 9692) * $signed(input_fmap_120[15:0]) +
	( 16'sd 26231) * $signed(input_fmap_121[15:0]) +
	( 16'sd 22347) * $signed(input_fmap_122[15:0]) +
	( 14'sd 8164) * $signed(input_fmap_123[15:0]) +
	( 16'sd 17432) * $signed(input_fmap_124[15:0]) +
	( 15'sd 8833) * $signed(input_fmap_125[15:0]) +
	( 16'sd 22133) * $signed(input_fmap_126[15:0]) +
	( 14'sd 6104) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 16'sd 23495) * $signed(input_fmap_0[15:0]) +
	( 15'sd 11853) * $signed(input_fmap_1[15:0]) +
	( 16'sd 28333) * $signed(input_fmap_2[15:0]) +
	( 16'sd 22943) * $signed(input_fmap_3[15:0]) +
	( 15'sd 11043) * $signed(input_fmap_4[15:0]) +
	( 16'sd 18930) * $signed(input_fmap_5[15:0]) +
	( 13'sd 3295) * $signed(input_fmap_6[15:0]) +
	( 16'sd 23878) * $signed(input_fmap_7[15:0]) +
	( 15'sd 10757) * $signed(input_fmap_8[15:0]) +
	( 15'sd 11679) * $signed(input_fmap_9[15:0]) +
	( 11'sd 970) * $signed(input_fmap_10[15:0]) +
	( 16'sd 31211) * $signed(input_fmap_11[15:0]) +
	( 14'sd 6893) * $signed(input_fmap_12[15:0]) +
	( 16'sd 21731) * $signed(input_fmap_13[15:0]) +
	( 15'sd 12485) * $signed(input_fmap_14[15:0]) +
	( 16'sd 24227) * $signed(input_fmap_15[15:0]) +
	( 13'sd 3033) * $signed(input_fmap_16[15:0]) +
	( 15'sd 14717) * $signed(input_fmap_17[15:0]) +
	( 16'sd 18302) * $signed(input_fmap_18[15:0]) +
	( 14'sd 5177) * $signed(input_fmap_19[15:0]) +
	( 15'sd 12923) * $signed(input_fmap_20[15:0]) +
	( 16'sd 21881) * $signed(input_fmap_21[15:0]) +
	( 15'sd 9600) * $signed(input_fmap_22[15:0]) +
	( 16'sd 22607) * $signed(input_fmap_23[15:0]) +
	( 16'sd 21863) * $signed(input_fmap_24[15:0]) +
	( 14'sd 4407) * $signed(input_fmap_25[15:0]) +
	( 16'sd 19370) * $signed(input_fmap_26[15:0]) +
	( 16'sd 16420) * $signed(input_fmap_27[15:0]) +
	( 14'sd 7026) * $signed(input_fmap_28[15:0]) +
	( 15'sd 11541) * $signed(input_fmap_29[15:0]) +
	( 13'sd 2269) * $signed(input_fmap_30[15:0]) +
	( 16'sd 30235) * $signed(input_fmap_31[15:0]) +
	( 12'sd 1907) * $signed(input_fmap_32[15:0]) +
	( 16'sd 32665) * $signed(input_fmap_33[15:0]) +
	( 15'sd 9636) * $signed(input_fmap_34[15:0]) +
	( 14'sd 7150) * $signed(input_fmap_35[15:0]) +
	( 16'sd 30496) * $signed(input_fmap_36[15:0]) +
	( 16'sd 28294) * $signed(input_fmap_37[15:0]) +
	( 16'sd 24952) * $signed(input_fmap_38[15:0]) +
	( 16'sd 19640) * $signed(input_fmap_39[15:0]) +
	( 16'sd 32027) * $signed(input_fmap_40[15:0]) +
	( 16'sd 21108) * $signed(input_fmap_41[15:0]) +
	( 14'sd 4910) * $signed(input_fmap_42[15:0]) +
	( 15'sd 13040) * $signed(input_fmap_43[15:0]) +
	( 16'sd 19684) * $signed(input_fmap_44[15:0]) +
	( 15'sd 15181) * $signed(input_fmap_45[15:0]) +
	( 16'sd 30213) * $signed(input_fmap_46[15:0]) +
	( 15'sd 15777) * $signed(input_fmap_47[15:0]) +
	( 15'sd 11086) * $signed(input_fmap_48[15:0]) +
	( 15'sd 11030) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22731) * $signed(input_fmap_50[15:0]) +
	( 16'sd 18025) * $signed(input_fmap_51[15:0]) +
	( 16'sd 26705) * $signed(input_fmap_52[15:0]) +
	( 15'sd 15437) * $signed(input_fmap_53[15:0]) +
	( 16'sd 24655) * $signed(input_fmap_54[15:0]) +
	( 16'sd 19165) * $signed(input_fmap_55[15:0]) +
	( 16'sd 24690) * $signed(input_fmap_56[15:0]) +
	( 16'sd 24926) * $signed(input_fmap_57[15:0]) +
	( 16'sd 23138) * $signed(input_fmap_58[15:0]) +
	( 13'sd 3612) * $signed(input_fmap_59[15:0]) +
	( 15'sd 11200) * $signed(input_fmap_60[15:0]) +
	( 16'sd 16486) * $signed(input_fmap_61[15:0]) +
	( 16'sd 28586) * $signed(input_fmap_62[15:0]) +
	( 16'sd 32761) * $signed(input_fmap_63[15:0]) +
	( 16'sd 30720) * $signed(input_fmap_64[15:0]) +
	( 16'sd 16920) * $signed(input_fmap_65[15:0]) +
	( 14'sd 5837) * $signed(input_fmap_66[15:0]) +
	( 16'sd 25475) * $signed(input_fmap_67[15:0]) +
	( 16'sd 25051) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31489) * $signed(input_fmap_69[15:0]) +
	( 14'sd 5801) * $signed(input_fmap_70[15:0]) +
	( 14'sd 7152) * $signed(input_fmap_71[15:0]) +
	( 15'sd 11185) * $signed(input_fmap_72[15:0]) +
	( 16'sd 30211) * $signed(input_fmap_73[15:0]) +
	( 16'sd 29501) * $signed(input_fmap_74[15:0]) +
	( 16'sd 26391) * $signed(input_fmap_75[15:0]) +
	( 15'sd 13255) * $signed(input_fmap_76[15:0]) +
	( 15'sd 16033) * $signed(input_fmap_77[15:0]) +
	( 14'sd 5413) * $signed(input_fmap_78[15:0]) +
	( 14'sd 8014) * $signed(input_fmap_79[15:0]) +
	( 16'sd 27896) * $signed(input_fmap_80[15:0]) +
	( 15'sd 12615) * $signed(input_fmap_81[15:0]) +
	( 16'sd 22507) * $signed(input_fmap_82[15:0]) +
	( 16'sd 28237) * $signed(input_fmap_83[15:0]) +
	( 13'sd 3857) * $signed(input_fmap_84[15:0]) +
	( 16'sd 29153) * $signed(input_fmap_85[15:0]) +
	( 15'sd 12973) * $signed(input_fmap_86[15:0]) +
	( 15'sd 9762) * $signed(input_fmap_87[15:0]) +
	( 16'sd 28045) * $signed(input_fmap_88[15:0]) +
	( 11'sd 596) * $signed(input_fmap_89[15:0]) +
	( 12'sd 1770) * $signed(input_fmap_90[15:0]) +
	( 15'sd 13179) * $signed(input_fmap_91[15:0]) +
	( 15'sd 15666) * $signed(input_fmap_92[15:0]) +
	( 13'sd 3536) * $signed(input_fmap_93[15:0]) +
	( 16'sd 19342) * $signed(input_fmap_94[15:0]) +
	( 15'sd 8986) * $signed(input_fmap_95[15:0]) +
	( 15'sd 16199) * $signed(input_fmap_96[15:0]) +
	( 16'sd 24928) * $signed(input_fmap_97[15:0]) +
	( 16'sd 30598) * $signed(input_fmap_98[15:0]) +
	( 16'sd 30540) * $signed(input_fmap_99[15:0]) +
	( 16'sd 22981) * $signed(input_fmap_100[15:0]) +
	( 16'sd 18071) * $signed(input_fmap_101[15:0]) +
	( 15'sd 8906) * $signed(input_fmap_102[15:0]) +
	( 15'sd 12274) * $signed(input_fmap_103[15:0]) +
	( 16'sd 29470) * $signed(input_fmap_104[15:0]) +
	( 16'sd 23812) * $signed(input_fmap_105[15:0]) +
	( 16'sd 17830) * $signed(input_fmap_106[15:0]) +
	( 16'sd 32174) * $signed(input_fmap_107[15:0]) +
	( 13'sd 2554) * $signed(input_fmap_108[15:0]) +
	( 16'sd 23534) * $signed(input_fmap_109[15:0]) +
	( 16'sd 29622) * $signed(input_fmap_110[15:0]) +
	( 16'sd 31259) * $signed(input_fmap_111[15:0]) +
	( 16'sd 28897) * $signed(input_fmap_112[15:0]) +
	( 16'sd 18659) * $signed(input_fmap_113[15:0]) +
	( 16'sd 26307) * $signed(input_fmap_114[15:0]) +
	( 14'sd 5436) * $signed(input_fmap_115[15:0]) +
	( 16'sd 18361) * $signed(input_fmap_116[15:0]) +
	( 16'sd 31731) * $signed(input_fmap_117[15:0]) +
	( 15'sd 9920) * $signed(input_fmap_118[15:0]) +
	( 15'sd 9026) * $signed(input_fmap_119[15:0]) +
	( 14'sd 4976) * $signed(input_fmap_120[15:0]) +
	( 14'sd 5848) * $signed(input_fmap_121[15:0]) +
	( 16'sd 22655) * $signed(input_fmap_122[15:0]) +
	( 16'sd 30868) * $signed(input_fmap_123[15:0]) +
	( 16'sd 24427) * $signed(input_fmap_124[15:0]) +
	( 15'sd 12763) * $signed(input_fmap_125[15:0]) +
	( 15'sd 13324) * $signed(input_fmap_126[15:0]) +
	( 16'sd 16900) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 15'sd 10096) * $signed(input_fmap_0[15:0]) +
	( 16'sd 28109) * $signed(input_fmap_1[15:0]) +
	( 16'sd 19661) * $signed(input_fmap_2[15:0]) +
	( 11'sd 829) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30427) * $signed(input_fmap_4[15:0]) +
	( 16'sd 27944) * $signed(input_fmap_5[15:0]) +
	( 14'sd 6505) * $signed(input_fmap_6[15:0]) +
	( 16'sd 20682) * $signed(input_fmap_7[15:0]) +
	( 15'sd 16163) * $signed(input_fmap_8[15:0]) +
	( 16'sd 29656) * $signed(input_fmap_9[15:0]) +
	( 16'sd 16448) * $signed(input_fmap_10[15:0]) +
	( 16'sd 26554) * $signed(input_fmap_11[15:0]) +
	( 14'sd 5272) * $signed(input_fmap_12[15:0]) +
	( 16'sd 29096) * $signed(input_fmap_13[15:0]) +
	( 16'sd 32151) * $signed(input_fmap_14[15:0]) +
	( 13'sd 3396) * $signed(input_fmap_15[15:0]) +
	( 16'sd 16747) * $signed(input_fmap_16[15:0]) +
	( 15'sd 11760) * $signed(input_fmap_17[15:0]) +
	( 15'sd 10978) * $signed(input_fmap_18[15:0]) +
	( 16'sd 25052) * $signed(input_fmap_19[15:0]) +
	( 16'sd 16534) * $signed(input_fmap_20[15:0]) +
	( 13'sd 3556) * $signed(input_fmap_21[15:0]) +
	( 15'sd 8484) * $signed(input_fmap_22[15:0]) +
	( 16'sd 29714) * $signed(input_fmap_23[15:0]) +
	( 16'sd 25254) * $signed(input_fmap_24[15:0]) +
	( 16'sd 30631) * $signed(input_fmap_25[15:0]) +
	( 16'sd 28459) * $signed(input_fmap_26[15:0]) +
	( 15'sd 12359) * $signed(input_fmap_27[15:0]) +
	( 13'sd 4031) * $signed(input_fmap_28[15:0]) +
	( 15'sd 12215) * $signed(input_fmap_29[15:0]) +
	( 15'sd 11316) * $signed(input_fmap_30[15:0]) +
	( 16'sd 18900) * $signed(input_fmap_31[15:0]) +
	( 16'sd 20662) * $signed(input_fmap_32[15:0]) +
	( 15'sd 9535) * $signed(input_fmap_33[15:0]) +
	( 16'sd 30076) * $signed(input_fmap_34[15:0]) +
	( 16'sd 23621) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11688) * $signed(input_fmap_36[15:0]) +
	( 16'sd 27089) * $signed(input_fmap_37[15:0]) +
	( 14'sd 5499) * $signed(input_fmap_38[15:0]) +
	( 16'sd 31045) * $signed(input_fmap_39[15:0]) +
	( 16'sd 17011) * $signed(input_fmap_40[15:0]) +
	( 15'sd 16010) * $signed(input_fmap_41[15:0]) +
	( 12'sd 1174) * $signed(input_fmap_42[15:0]) +
	( 14'sd 6240) * $signed(input_fmap_43[15:0]) +
	( 15'sd 12189) * $signed(input_fmap_44[15:0]) +
	( 15'sd 8901) * $signed(input_fmap_45[15:0]) +
	( 16'sd 24470) * $signed(input_fmap_46[15:0]) +
	( 16'sd 16649) * $signed(input_fmap_47[15:0]) +
	( 11'sd 578) * $signed(input_fmap_48[15:0]) +
	( 16'sd 18763) * $signed(input_fmap_49[15:0]) +
	( 13'sd 2582) * $signed(input_fmap_50[15:0]) +
	( 16'sd 28661) * $signed(input_fmap_51[15:0]) +
	( 15'sd 9120) * $signed(input_fmap_52[15:0]) +
	( 16'sd 32688) * $signed(input_fmap_53[15:0]) +
	( 15'sd 13684) * $signed(input_fmap_54[15:0]) +
	( 14'sd 6101) * $signed(input_fmap_55[15:0]) +
	( 16'sd 21675) * $signed(input_fmap_56[15:0]) +
	( 16'sd 24723) * $signed(input_fmap_57[15:0]) +
	( 16'sd 23646) * $signed(input_fmap_58[15:0]) +
	( 14'sd 5927) * $signed(input_fmap_59[15:0]) +
	( 16'sd 22768) * $signed(input_fmap_60[15:0]) +
	( 14'sd 7192) * $signed(input_fmap_61[15:0]) +
	( 16'sd 19538) * $signed(input_fmap_62[15:0]) +
	( 16'sd 31480) * $signed(input_fmap_63[15:0]) +
	( 14'sd 4179) * $signed(input_fmap_64[15:0]) +
	( 16'sd 29179) * $signed(input_fmap_65[15:0]) +
	( 14'sd 5834) * $signed(input_fmap_66[15:0]) +
	( 16'sd 25264) * $signed(input_fmap_67[15:0]) +
	( 16'sd 21230) * $signed(input_fmap_68[15:0]) +
	( 16'sd 16512) * $signed(input_fmap_69[15:0]) +
	( 16'sd 16841) * $signed(input_fmap_70[15:0]) +
	( 16'sd 24839) * $signed(input_fmap_71[15:0]) +
	( 8'sd 116) * $signed(input_fmap_72[15:0]) +
	( 15'sd 10778) * $signed(input_fmap_73[15:0]) +
	( 14'sd 6306) * $signed(input_fmap_74[15:0]) +
	( 13'sd 3783) * $signed(input_fmap_75[15:0]) +
	( 16'sd 16587) * $signed(input_fmap_76[15:0]) +
	( 16'sd 27222) * $signed(input_fmap_77[15:0]) +
	( 15'sd 15612) * $signed(input_fmap_78[15:0]) +
	( 15'sd 12165) * $signed(input_fmap_79[15:0]) +
	( 15'sd 12709) * $signed(input_fmap_80[15:0]) +
	( 15'sd 10567) * $signed(input_fmap_81[15:0]) +
	( 15'sd 11103) * $signed(input_fmap_82[15:0]) +
	( 15'sd 14993) * $signed(input_fmap_83[15:0]) +
	( 16'sd 18447) * $signed(input_fmap_84[15:0]) +
	( 16'sd 26486) * $signed(input_fmap_85[15:0]) +
	( 14'sd 6614) * $signed(input_fmap_86[15:0]) +
	( 15'sd 12400) * $signed(input_fmap_87[15:0]) +
	( 13'sd 3893) * $signed(input_fmap_88[15:0]) +
	( 14'sd 6100) * $signed(input_fmap_89[15:0]) +
	( 15'sd 12730) * $signed(input_fmap_90[15:0]) +
	( 15'sd 16374) * $signed(input_fmap_91[15:0]) +
	( 15'sd 14653) * $signed(input_fmap_92[15:0]) +
	( 16'sd 32701) * $signed(input_fmap_93[15:0]) +
	( 13'sd 3071) * $signed(input_fmap_94[15:0]) +
	( 9'sd 220) * $signed(input_fmap_95[15:0]) +
	( 15'sd 10848) * $signed(input_fmap_96[15:0]) +
	( 16'sd 26658) * $signed(input_fmap_97[15:0]) +
	( 14'sd 4506) * $signed(input_fmap_98[15:0]) +
	( 16'sd 30305) * $signed(input_fmap_99[15:0]) +
	( 16'sd 27372) * $signed(input_fmap_100[15:0]) +
	( 10'sd 321) * $signed(input_fmap_101[15:0]) +
	( 16'sd 18132) * $signed(input_fmap_102[15:0]) +
	( 14'sd 6158) * $signed(input_fmap_103[15:0]) +
	( 15'sd 10278) * $signed(input_fmap_104[15:0]) +
	( 14'sd 6631) * $signed(input_fmap_105[15:0]) +
	( 16'sd 29830) * $signed(input_fmap_106[15:0]) +
	( 16'sd 29188) * $signed(input_fmap_107[15:0]) +
	( 16'sd 26227) * $signed(input_fmap_108[15:0]) +
	( 16'sd 31823) * $signed(input_fmap_109[15:0]) +
	( 13'sd 3267) * $signed(input_fmap_110[15:0]) +
	( 16'sd 26955) * $signed(input_fmap_111[15:0]) +
	( 16'sd 22636) * $signed(input_fmap_112[15:0]) +
	( 13'sd 3648) * $signed(input_fmap_113[15:0]) +
	( 16'sd 20564) * $signed(input_fmap_114[15:0]) +
	( 14'sd 6011) * $signed(input_fmap_115[15:0]) +
	( 14'sd 4274) * $signed(input_fmap_116[15:0]) +
	( 7'sd 49) * $signed(input_fmap_117[15:0]) +
	( 16'sd 29747) * $signed(input_fmap_118[15:0]) +
	( 16'sd 30516) * $signed(input_fmap_119[15:0]) +
	( 16'sd 25865) * $signed(input_fmap_120[15:0]) +
	( 16'sd 28042) * $signed(input_fmap_121[15:0]) +
	( 15'sd 10506) * $signed(input_fmap_122[15:0]) +
	( 16'sd 23789) * $signed(input_fmap_123[15:0]) +
	( 16'sd 17088) * $signed(input_fmap_124[15:0]) +
	( 16'sd 19057) * $signed(input_fmap_125[15:0]) +
	( 11'sd 979) * $signed(input_fmap_126[15:0]) +
	( 14'sd 6992) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 16'sd 27964) * $signed(input_fmap_0[15:0]) +
	( 16'sd 28107) * $signed(input_fmap_1[15:0]) +
	( 16'sd 18419) * $signed(input_fmap_2[15:0]) +
	( 16'sd 16384) * $signed(input_fmap_3[15:0]) +
	( 13'sd 2927) * $signed(input_fmap_4[15:0]) +
	( 14'sd 5316) * $signed(input_fmap_5[15:0]) +
	( 16'sd 30460) * $signed(input_fmap_6[15:0]) +
	( 16'sd 28910) * $signed(input_fmap_7[15:0]) +
	( 15'sd 11557) * $signed(input_fmap_8[15:0]) +
	( 15'sd 13419) * $signed(input_fmap_9[15:0]) +
	( 14'sd 5784) * $signed(input_fmap_10[15:0]) +
	( 14'sd 6893) * $signed(input_fmap_11[15:0]) +
	( 16'sd 22827) * $signed(input_fmap_12[15:0]) +
	( 16'sd 17169) * $signed(input_fmap_13[15:0]) +
	( 15'sd 10852) * $signed(input_fmap_14[15:0]) +
	( 15'sd 11148) * $signed(input_fmap_15[15:0]) +
	( 16'sd 21292) * $signed(input_fmap_16[15:0]) +
	( 16'sd 24911) * $signed(input_fmap_17[15:0]) +
	( 16'sd 30933) * $signed(input_fmap_18[15:0]) +
	( 13'sd 3410) * $signed(input_fmap_19[15:0]) +
	( 15'sd 13186) * $signed(input_fmap_20[15:0]) +
	( 16'sd 24753) * $signed(input_fmap_21[15:0]) +
	( 16'sd 25990) * $signed(input_fmap_22[15:0]) +
	( 16'sd 27127) * $signed(input_fmap_23[15:0]) +
	( 15'sd 13000) * $signed(input_fmap_24[15:0]) +
	( 16'sd 22839) * $signed(input_fmap_25[15:0]) +
	( 15'sd 12057) * $signed(input_fmap_26[15:0]) +
	( 15'sd 10638) * $signed(input_fmap_27[15:0]) +
	( 6'sd 29) * $signed(input_fmap_28[15:0]) +
	( 10'sd 393) * $signed(input_fmap_29[15:0]) +
	( 15'sd 16035) * $signed(input_fmap_30[15:0]) +
	( 14'sd 6300) * $signed(input_fmap_31[15:0]) +
	( 15'sd 9134) * $signed(input_fmap_32[15:0]) +
	( 11'sd 756) * $signed(input_fmap_33[15:0]) +
	( 15'sd 15543) * $signed(input_fmap_34[15:0]) +
	( 16'sd 19138) * $signed(input_fmap_35[15:0]) +
	( 15'sd 12957) * $signed(input_fmap_36[15:0]) +
	( 16'sd 28404) * $signed(input_fmap_37[15:0]) +
	( 16'sd 28990) * $signed(input_fmap_38[15:0]) +
	( 16'sd 25357) * $signed(input_fmap_39[15:0]) +
	( 15'sd 14959) * $signed(input_fmap_40[15:0]) +
	( 12'sd 2024) * $signed(input_fmap_41[15:0]) +
	( 16'sd 24608) * $signed(input_fmap_42[15:0]) +
	( 16'sd 31982) * $signed(input_fmap_43[15:0]) +
	( 15'sd 12007) * $signed(input_fmap_44[15:0]) +
	( 15'sd 10737) * $signed(input_fmap_45[15:0]) +
	( 16'sd 17971) * $signed(input_fmap_46[15:0]) +
	( 16'sd 24212) * $signed(input_fmap_47[15:0]) +
	( 14'sd 7517) * $signed(input_fmap_48[15:0]) +
	( 15'sd 15253) * $signed(input_fmap_49[15:0]) +
	( 16'sd 24939) * $signed(input_fmap_50[15:0]) +
	( 13'sd 3963) * $signed(input_fmap_51[15:0]) +
	( 15'sd 10675) * $signed(input_fmap_52[15:0]) +
	( 12'sd 1256) * $signed(input_fmap_53[15:0]) +
	( 16'sd 20516) * $signed(input_fmap_54[15:0]) +
	( 14'sd 6957) * $signed(input_fmap_55[15:0]) +
	( 15'sd 9387) * $signed(input_fmap_56[15:0]) +
	( 16'sd 29464) * $signed(input_fmap_57[15:0]) +
	( 16'sd 27692) * $signed(input_fmap_58[15:0]) +
	( 16'sd 23904) * $signed(input_fmap_59[15:0]) +
	( 15'sd 13502) * $signed(input_fmap_60[15:0]) +
	( 14'sd 7509) * $signed(input_fmap_61[15:0]) +
	( 15'sd 16232) * $signed(input_fmap_62[15:0]) +
	( 14'sd 4697) * $signed(input_fmap_63[15:0]) +
	( 14'sd 6810) * $signed(input_fmap_64[15:0]) +
	( 15'sd 9462) * $signed(input_fmap_65[15:0]) +
	( 16'sd 23373) * $signed(input_fmap_66[15:0]) +
	( 14'sd 6203) * $signed(input_fmap_67[15:0]) +
	( 16'sd 31762) * $signed(input_fmap_68[15:0]) +
	( 16'sd 26184) * $signed(input_fmap_69[15:0]) +
	( 15'sd 13538) * $signed(input_fmap_70[15:0]) +
	( 15'sd 14549) * $signed(input_fmap_71[15:0]) +
	( 15'sd 9192) * $signed(input_fmap_72[15:0]) +
	( 13'sd 3371) * $signed(input_fmap_73[15:0]) +
	( 15'sd 15747) * $signed(input_fmap_74[15:0]) +
	( 15'sd 12804) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19096) * $signed(input_fmap_76[15:0]) +
	( 16'sd 22712) * $signed(input_fmap_77[15:0]) +
	( 15'sd 10079) * $signed(input_fmap_78[15:0]) +
	( 16'sd 28564) * $signed(input_fmap_79[15:0]) +
	( 14'sd 7343) * $signed(input_fmap_80[15:0]) +
	( 15'sd 11226) * $signed(input_fmap_81[15:0]) +
	( 13'sd 4016) * $signed(input_fmap_82[15:0]) +
	( 15'sd 8999) * $signed(input_fmap_83[15:0]) +
	( 14'sd 5132) * $signed(input_fmap_84[15:0]) +
	( 14'sd 5197) * $signed(input_fmap_85[15:0]) +
	( 14'sd 5501) * $signed(input_fmap_86[15:0]) +
	( 15'sd 9275) * $signed(input_fmap_87[15:0]) +
	( 16'sd 25650) * $signed(input_fmap_88[15:0]) +
	( 15'sd 15027) * $signed(input_fmap_89[15:0]) +
	( 10'sd 489) * $signed(input_fmap_90[15:0]) +
	( 16'sd 17694) * $signed(input_fmap_91[15:0]) +
	( 12'sd 2010) * $signed(input_fmap_92[15:0]) +
	( 16'sd 25252) * $signed(input_fmap_93[15:0]) +
	( 15'sd 8993) * $signed(input_fmap_94[15:0]) +
	( 15'sd 16155) * $signed(input_fmap_95[15:0]) +
	( 16'sd 28466) * $signed(input_fmap_96[15:0]) +
	( 16'sd 32252) * $signed(input_fmap_97[15:0]) +
	( 16'sd 19291) * $signed(input_fmap_98[15:0]) +
	( 16'sd 16593) * $signed(input_fmap_99[15:0]) +
	( 15'sd 10539) * $signed(input_fmap_100[15:0]) +
	( 16'sd 31241) * $signed(input_fmap_101[15:0]) +
	( 16'sd 23496) * $signed(input_fmap_102[15:0]) +
	( 14'sd 5391) * $signed(input_fmap_103[15:0]) +
	( 16'sd 16776) * $signed(input_fmap_104[15:0]) +
	( 16'sd 25208) * $signed(input_fmap_105[15:0]) +
	( 14'sd 6792) * $signed(input_fmap_106[15:0]) +
	( 16'sd 30913) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15472) * $signed(input_fmap_108[15:0]) +
	( 16'sd 25709) * $signed(input_fmap_109[15:0]) +
	( 16'sd 21932) * $signed(input_fmap_110[15:0]) +
	( 14'sd 5982) * $signed(input_fmap_111[15:0]) +
	( 15'sd 12455) * $signed(input_fmap_112[15:0]) +
	( 15'sd 12332) * $signed(input_fmap_113[15:0]) +
	( 15'sd 13700) * $signed(input_fmap_114[15:0]) +
	( 16'sd 23283) * $signed(input_fmap_115[15:0]) +
	( 13'sd 3292) * $signed(input_fmap_116[15:0]) +
	( 14'sd 7625) * $signed(input_fmap_117[15:0]) +
	( 16'sd 28321) * $signed(input_fmap_118[15:0]) +
	( 16'sd 24308) * $signed(input_fmap_119[15:0]) +
	( 13'sd 3870) * $signed(input_fmap_120[15:0]) +
	( 16'sd 32310) * $signed(input_fmap_121[15:0]) +
	( 12'sd 1571) * $signed(input_fmap_122[15:0]) +
	( 15'sd 10227) * $signed(input_fmap_123[15:0]) +
	( 16'sd 29576) * $signed(input_fmap_124[15:0]) +
	( 16'sd 23550) * $signed(input_fmap_125[15:0]) +
	( 15'sd 9753) * $signed(input_fmap_126[15:0]) +
	( 13'sd 3235) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 15'sd 15876) * $signed(input_fmap_0[15:0]) +
	( 14'sd 7475) * $signed(input_fmap_1[15:0]) +
	( 16'sd 17972) * $signed(input_fmap_2[15:0]) +
	( 15'sd 12607) * $signed(input_fmap_3[15:0]) +
	( 15'sd 13192) * $signed(input_fmap_4[15:0]) +
	( 16'sd 22451) * $signed(input_fmap_5[15:0]) +
	( 15'sd 13701) * $signed(input_fmap_6[15:0]) +
	( 13'sd 3544) * $signed(input_fmap_7[15:0]) +
	( 16'sd 26091) * $signed(input_fmap_8[15:0]) +
	( 14'sd 5732) * $signed(input_fmap_9[15:0]) +
	( 16'sd 19088) * $signed(input_fmap_10[15:0]) +
	( 15'sd 8632) * $signed(input_fmap_11[15:0]) +
	( 15'sd 9309) * $signed(input_fmap_12[15:0]) +
	( 13'sd 3378) * $signed(input_fmap_13[15:0]) +
	( 16'sd 23955) * $signed(input_fmap_14[15:0]) +
	( 16'sd 30645) * $signed(input_fmap_15[15:0]) +
	( 16'sd 26390) * $signed(input_fmap_16[15:0]) +
	( 15'sd 16113) * $signed(input_fmap_17[15:0]) +
	( 16'sd 20575) * $signed(input_fmap_18[15:0]) +
	( 16'sd 17241) * $signed(input_fmap_19[15:0]) +
	( 15'sd 11350) * $signed(input_fmap_20[15:0]) +
	( 16'sd 28895) * $signed(input_fmap_21[15:0]) +
	( 15'sd 15681) * $signed(input_fmap_22[15:0]) +
	( 15'sd 12721) * $signed(input_fmap_23[15:0]) +
	( 16'sd 26300) * $signed(input_fmap_24[15:0]) +
	( 12'sd 1973) * $signed(input_fmap_25[15:0]) +
	( 16'sd 29227) * $signed(input_fmap_26[15:0]) +
	( 16'sd 31897) * $signed(input_fmap_27[15:0]) +
	( 16'sd 32251) * $signed(input_fmap_28[15:0]) +
	( 16'sd 21960) * $signed(input_fmap_29[15:0]) +
	( 16'sd 32598) * $signed(input_fmap_30[15:0]) +
	( 16'sd 30961) * $signed(input_fmap_31[15:0]) +
	( 16'sd 30311) * $signed(input_fmap_32[15:0]) +
	( 14'sd 5125) * $signed(input_fmap_33[15:0]) +
	( 15'sd 13077) * $signed(input_fmap_34[15:0]) +
	( 16'sd 30294) * $signed(input_fmap_35[15:0]) +
	( 16'sd 24971) * $signed(input_fmap_36[15:0]) +
	( 15'sd 11666) * $signed(input_fmap_37[15:0]) +
	( 16'sd 18616) * $signed(input_fmap_38[15:0]) +
	( 16'sd 31673) * $signed(input_fmap_39[15:0]) +
	( 14'sd 5541) * $signed(input_fmap_40[15:0]) +
	( 16'sd 27877) * $signed(input_fmap_41[15:0]) +
	( 15'sd 12520) * $signed(input_fmap_42[15:0]) +
	( 15'sd 15944) * $signed(input_fmap_43[15:0]) +
	( 15'sd 9304) * $signed(input_fmap_44[15:0]) +
	( 15'sd 16121) * $signed(input_fmap_45[15:0]) +
	( 15'sd 8725) * $signed(input_fmap_46[15:0]) +
	( 16'sd 25679) * $signed(input_fmap_47[15:0]) +
	( 16'sd 19896) * $signed(input_fmap_48[15:0]) +
	( 14'sd 4228) * $signed(input_fmap_49[15:0]) +
	( 16'sd 28441) * $signed(input_fmap_50[15:0]) +
	( 16'sd 18296) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3515) * $signed(input_fmap_52[15:0]) +
	( 16'sd 32234) * $signed(input_fmap_53[15:0]) +
	( 16'sd 17471) * $signed(input_fmap_54[15:0]) +
	( 16'sd 21092) * $signed(input_fmap_55[15:0]) +
	( 13'sd 2946) * $signed(input_fmap_56[15:0]) +
	( 16'sd 32572) * $signed(input_fmap_57[15:0]) +
	( 14'sd 6166) * $signed(input_fmap_58[15:0]) +
	( 16'sd 30592) * $signed(input_fmap_59[15:0]) +
	( 13'sd 2614) * $signed(input_fmap_60[15:0]) +
	( 16'sd 30039) * $signed(input_fmap_61[15:0]) +
	( 12'sd 1768) * $signed(input_fmap_62[15:0]) +
	( 16'sd 30818) * $signed(input_fmap_63[15:0]) +
	( 15'sd 11349) * $signed(input_fmap_64[15:0]) +
	( 15'sd 14757) * $signed(input_fmap_65[15:0]) +
	( 15'sd 11370) * $signed(input_fmap_66[15:0]) +
	( 15'sd 15376) * $signed(input_fmap_67[15:0]) +
	( 15'sd 9738) * $signed(input_fmap_68[15:0]) +
	( 15'sd 11627) * $signed(input_fmap_69[15:0]) +
	( 14'sd 6836) * $signed(input_fmap_70[15:0]) +
	( 16'sd 21117) * $signed(input_fmap_71[15:0]) +
	( 12'sd 1260) * $signed(input_fmap_72[15:0]) +
	( 16'sd 18439) * $signed(input_fmap_73[15:0]) +
	( 16'sd 23302) * $signed(input_fmap_74[15:0]) +
	( 16'sd 29056) * $signed(input_fmap_75[15:0]) +
	( 15'sd 13242) * $signed(input_fmap_76[15:0]) +
	( 15'sd 12537) * $signed(input_fmap_77[15:0]) +
	( 16'sd 20223) * $signed(input_fmap_78[15:0]) +
	( 16'sd 31349) * $signed(input_fmap_79[15:0]) +
	( 16'sd 29541) * $signed(input_fmap_80[15:0]) +
	( 16'sd 16837) * $signed(input_fmap_81[15:0]) +
	( 16'sd 18197) * $signed(input_fmap_82[15:0]) +
	( 16'sd 20113) * $signed(input_fmap_83[15:0]) +
	( 16'sd 17676) * $signed(input_fmap_84[15:0]) +
	( 15'sd 13382) * $signed(input_fmap_85[15:0]) +
	( 14'sd 7155) * $signed(input_fmap_86[15:0]) +
	( 15'sd 13147) * $signed(input_fmap_87[15:0]) +
	( 14'sd 4128) * $signed(input_fmap_88[15:0]) +
	( 14'sd 6001) * $signed(input_fmap_89[15:0]) +
	( 15'sd 8873) * $signed(input_fmap_90[15:0]) +
	( 8'sd 101) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25253) * $signed(input_fmap_92[15:0]) +
	( 16'sd 24215) * $signed(input_fmap_93[15:0]) +
	( 15'sd 15955) * $signed(input_fmap_94[15:0]) +
	( 16'sd 26178) * $signed(input_fmap_95[15:0]) +
	( 16'sd 31105) * $signed(input_fmap_96[15:0]) +
	( 16'sd 16594) * $signed(input_fmap_97[15:0]) +
	( 16'sd 27797) * $signed(input_fmap_98[15:0]) +
	( 12'sd 1232) * $signed(input_fmap_99[15:0]) +
	( 7'sd 51) * $signed(input_fmap_100[15:0]) +
	( 16'sd 17204) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5629) * $signed(input_fmap_102[15:0]) +
	( 16'sd 18334) * $signed(input_fmap_103[15:0]) +
	( 16'sd 30806) * $signed(input_fmap_104[15:0]) +
	( 16'sd 23662) * $signed(input_fmap_105[15:0]) +
	( 16'sd 19990) * $signed(input_fmap_106[15:0]) +
	( 16'sd 23811) * $signed(input_fmap_107[15:0]) +
	( 12'sd 1892) * $signed(input_fmap_108[15:0]) +
	( 14'sd 7248) * $signed(input_fmap_109[15:0]) +
	( 15'sd 12051) * $signed(input_fmap_110[15:0]) +
	( 15'sd 13323) * $signed(input_fmap_111[15:0]) +
	( 11'sd 582) * $signed(input_fmap_112[15:0]) +
	( 13'sd 3844) * $signed(input_fmap_113[15:0]) +
	( 16'sd 20965) * $signed(input_fmap_114[15:0]) +
	( 16'sd 30312) * $signed(input_fmap_115[15:0]) +
	( 10'sd 285) * $signed(input_fmap_116[15:0]) +
	( 16'sd 19249) * $signed(input_fmap_117[15:0]) +
	( 16'sd 26165) * $signed(input_fmap_118[15:0]) +
	( 14'sd 7450) * $signed(input_fmap_119[15:0]) +
	( 16'sd 22315) * $signed(input_fmap_120[15:0]) +
	( 15'sd 12491) * $signed(input_fmap_121[15:0]) +
	( 10'sd 406) * $signed(input_fmap_122[15:0]) +
	( 15'sd 11743) * $signed(input_fmap_123[15:0]) +
	( 16'sd 22020) * $signed(input_fmap_124[15:0]) +
	( 16'sd 28421) * $signed(input_fmap_125[15:0]) +
	( 16'sd 28066) * $signed(input_fmap_126[15:0]) +
	( 16'sd 20783) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 15'sd 13832) * $signed(input_fmap_0[15:0]) +
	( 16'sd 23235) * $signed(input_fmap_1[15:0]) +
	( 16'sd 27052) * $signed(input_fmap_2[15:0]) +
	( 13'sd 3122) * $signed(input_fmap_3[15:0]) +
	( 13'sd 3336) * $signed(input_fmap_4[15:0]) +
	( 16'sd 27182) * $signed(input_fmap_5[15:0]) +
	( 13'sd 3321) * $signed(input_fmap_6[15:0]) +
	( 15'sd 12521) * $signed(input_fmap_7[15:0]) +
	( 15'sd 10146) * $signed(input_fmap_8[15:0]) +
	( 14'sd 7028) * $signed(input_fmap_9[15:0]) +
	( 15'sd 15186) * $signed(input_fmap_10[15:0]) +
	( 16'sd 20672) * $signed(input_fmap_11[15:0]) +
	( 15'sd 15856) * $signed(input_fmap_12[15:0]) +
	( 16'sd 23890) * $signed(input_fmap_13[15:0]) +
	( 16'sd 19426) * $signed(input_fmap_14[15:0]) +
	( 15'sd 9337) * $signed(input_fmap_15[15:0]) +
	( 15'sd 12573) * $signed(input_fmap_16[15:0]) +
	( 16'sd 23682) * $signed(input_fmap_17[15:0]) +
	( 16'sd 31710) * $signed(input_fmap_18[15:0]) +
	( 16'sd 32057) * $signed(input_fmap_19[15:0]) +
	( 14'sd 4363) * $signed(input_fmap_20[15:0]) +
	( 13'sd 3096) * $signed(input_fmap_21[15:0]) +
	( 11'sd 980) * $signed(input_fmap_22[15:0]) +
	( 15'sd 11775) * $signed(input_fmap_23[15:0]) +
	( 15'sd 15549) * $signed(input_fmap_24[15:0]) +
	( 14'sd 7088) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22254) * $signed(input_fmap_26[15:0]) +
	( 15'sd 15071) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24080) * $signed(input_fmap_28[15:0]) +
	( 16'sd 31010) * $signed(input_fmap_29[15:0]) +
	( 15'sd 14163) * $signed(input_fmap_30[15:0]) +
	( 12'sd 1539) * $signed(input_fmap_31[15:0]) +
	( 16'sd 19508) * $signed(input_fmap_32[15:0]) +
	( 16'sd 17825) * $signed(input_fmap_33[15:0]) +
	( 15'sd 10093) * $signed(input_fmap_34[15:0]) +
	( 16'sd 18991) * $signed(input_fmap_35[15:0]) +
	( 15'sd 12996) * $signed(input_fmap_36[15:0]) +
	( 16'sd 30859) * $signed(input_fmap_37[15:0]) +
	( 11'sd 895) * $signed(input_fmap_38[15:0]) +
	( 16'sd 28656) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6950) * $signed(input_fmap_40[15:0]) +
	( 16'sd 31817) * $signed(input_fmap_41[15:0]) +
	( 13'sd 3736) * $signed(input_fmap_42[15:0]) +
	( 16'sd 19777) * $signed(input_fmap_43[15:0]) +
	( 16'sd 32379) * $signed(input_fmap_44[15:0]) +
	( 12'sd 1931) * $signed(input_fmap_45[15:0]) +
	( 16'sd 17096) * $signed(input_fmap_46[15:0]) +
	( 16'sd 29033) * $signed(input_fmap_47[15:0]) +
	( 16'sd 21930) * $signed(input_fmap_48[15:0]) +
	( 13'sd 3491) * $signed(input_fmap_49[15:0]) +
	( 15'sd 13835) * $signed(input_fmap_50[15:0]) +
	( 16'sd 28603) * $signed(input_fmap_51[15:0]) +
	( 16'sd 22225) * $signed(input_fmap_52[15:0]) +
	( 12'sd 1426) * $signed(input_fmap_53[15:0]) +
	( 15'sd 13125) * $signed(input_fmap_54[15:0]) +
	( 16'sd 25743) * $signed(input_fmap_55[15:0]) +
	( 16'sd 18400) * $signed(input_fmap_56[15:0]) +
	( 16'sd 21648) * $signed(input_fmap_57[15:0]) +
	( 15'sd 9274) * $signed(input_fmap_58[15:0]) +
	( 16'sd 23485) * $signed(input_fmap_59[15:0]) +
	( 16'sd 19040) * $signed(input_fmap_60[15:0]) +
	( 16'sd 28390) * $signed(input_fmap_61[15:0]) +
	( 16'sd 21301) * $signed(input_fmap_62[15:0]) +
	( 15'sd 14568) * $signed(input_fmap_63[15:0]) +
	( 16'sd 21215) * $signed(input_fmap_64[15:0]) +
	( 16'sd 24943) * $signed(input_fmap_65[15:0]) +
	( 16'sd 21535) * $signed(input_fmap_66[15:0]) +
	( 14'sd 6224) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26903) * $signed(input_fmap_68[15:0]) +
	( 16'sd 22969) * $signed(input_fmap_69[15:0]) +
	( 16'sd 32655) * $signed(input_fmap_70[15:0]) +
	( 15'sd 15546) * $signed(input_fmap_71[15:0]) +
	( 16'sd 30497) * $signed(input_fmap_72[15:0]) +
	( 16'sd 24997) * $signed(input_fmap_73[15:0]) +
	( 14'sd 6526) * $signed(input_fmap_74[15:0]) +
	( 15'sd 11660) * $signed(input_fmap_75[15:0]) +
	( 14'sd 8026) * $signed(input_fmap_76[15:0]) +
	( 15'sd 12016) * $signed(input_fmap_77[15:0]) +
	( 15'sd 14062) * $signed(input_fmap_78[15:0]) +
	( 16'sd 30345) * $signed(input_fmap_79[15:0]) +
	( 16'sd 30126) * $signed(input_fmap_80[15:0]) +
	( 14'sd 7918) * $signed(input_fmap_81[15:0]) +
	( 16'sd 27139) * $signed(input_fmap_82[15:0]) +
	( 15'sd 10760) * $signed(input_fmap_83[15:0]) +
	( 15'sd 11268) * $signed(input_fmap_84[15:0]) +
	( 16'sd 27339) * $signed(input_fmap_85[15:0]) +
	( 15'sd 10114) * $signed(input_fmap_86[15:0]) +
	( 8'sd 125) * $signed(input_fmap_87[15:0]) +
	( 14'sd 7352) * $signed(input_fmap_88[15:0]) +
	( 16'sd 31181) * $signed(input_fmap_89[15:0]) +
	( 15'sd 9974) * $signed(input_fmap_90[15:0]) +
	( 16'sd 27355) * $signed(input_fmap_91[15:0]) +
	( 16'sd 19685) * $signed(input_fmap_92[15:0]) +
	( 15'sd 12045) * $signed(input_fmap_93[15:0]) +
	( 16'sd 22734) * $signed(input_fmap_94[15:0]) +
	( 16'sd 21865) * $signed(input_fmap_95[15:0]) +
	( 14'sd 7876) * $signed(input_fmap_96[15:0]) +
	( 16'sd 30305) * $signed(input_fmap_97[15:0]) +
	( 16'sd 26834) * $signed(input_fmap_98[15:0]) +
	( 15'sd 8546) * $signed(input_fmap_99[15:0]) +
	( 14'sd 7924) * $signed(input_fmap_100[15:0]) +
	( 16'sd 18618) * $signed(input_fmap_101[15:0]) +
	( 15'sd 15869) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28300) * $signed(input_fmap_103[15:0]) +
	( 16'sd 19609) * $signed(input_fmap_104[15:0]) +
	( 16'sd 25137) * $signed(input_fmap_105[15:0]) +
	( 16'sd 24511) * $signed(input_fmap_106[15:0]) +
	( 16'sd 22244) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15590) * $signed(input_fmap_108[15:0]) +
	( 15'sd 13863) * $signed(input_fmap_109[15:0]) +
	( 16'sd 25730) * $signed(input_fmap_110[15:0]) +
	( 15'sd 12155) * $signed(input_fmap_111[15:0]) +
	( 16'sd 24957) * $signed(input_fmap_112[15:0]) +
	( 16'sd 22101) * $signed(input_fmap_113[15:0]) +
	( 14'sd 5717) * $signed(input_fmap_114[15:0]) +
	( 14'sd 5715) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26896) * $signed(input_fmap_116[15:0]) +
	( 15'sd 12679) * $signed(input_fmap_117[15:0]) +
	( 13'sd 2961) * $signed(input_fmap_118[15:0]) +
	( 14'sd 4371) * $signed(input_fmap_119[15:0]) +
	( 16'sd 25903) * $signed(input_fmap_120[15:0]) +
	( 16'sd 31359) * $signed(input_fmap_121[15:0]) +
	( 16'sd 27278) * $signed(input_fmap_122[15:0]) +
	( 16'sd 24293) * $signed(input_fmap_123[15:0]) +
	( 13'sd 3217) * $signed(input_fmap_124[15:0]) +
	( 16'sd 16417) * $signed(input_fmap_125[15:0]) +
	( 16'sd 30956) * $signed(input_fmap_126[15:0]) +
	( 16'sd 18131) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 15'sd 13583) * $signed(input_fmap_0[15:0]) +
	( 15'sd 12707) * $signed(input_fmap_1[15:0]) +
	( 15'sd 12209) * $signed(input_fmap_2[15:0]) +
	( 16'sd 26167) * $signed(input_fmap_3[15:0]) +
	( 15'sd 10546) * $signed(input_fmap_4[15:0]) +
	( 16'sd 20411) * $signed(input_fmap_5[15:0]) +
	( 16'sd 31672) * $signed(input_fmap_6[15:0]) +
	( 12'sd 1167) * $signed(input_fmap_7[15:0]) +
	( 16'sd 23563) * $signed(input_fmap_8[15:0]) +
	( 13'sd 2628) * $signed(input_fmap_9[15:0]) +
	( 16'sd 26066) * $signed(input_fmap_10[15:0]) +
	( 16'sd 24289) * $signed(input_fmap_11[15:0]) +
	( 14'sd 4314) * $signed(input_fmap_12[15:0]) +
	( 15'sd 10147) * $signed(input_fmap_13[15:0]) +
	( 16'sd 25235) * $signed(input_fmap_14[15:0]) +
	( 13'sd 3638) * $signed(input_fmap_15[15:0]) +
	( 15'sd 13902) * $signed(input_fmap_16[15:0]) +
	( 15'sd 15847) * $signed(input_fmap_17[15:0]) +
	( 14'sd 4773) * $signed(input_fmap_18[15:0]) +
	( 15'sd 16204) * $signed(input_fmap_19[15:0]) +
	( 10'sd 262) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17564) * $signed(input_fmap_21[15:0]) +
	( 16'sd 19096) * $signed(input_fmap_22[15:0]) +
	( 11'sd 920) * $signed(input_fmap_23[15:0]) +
	( 16'sd 27753) * $signed(input_fmap_24[15:0]) +
	( 16'sd 31523) * $signed(input_fmap_25[15:0]) +
	( 16'sd 32676) * $signed(input_fmap_26[15:0]) +
	( 16'sd 23491) * $signed(input_fmap_27[15:0]) +
	( 13'sd 4045) * $signed(input_fmap_28[15:0]) +
	( 15'sd 11221) * $signed(input_fmap_29[15:0]) +
	( 15'sd 10213) * $signed(input_fmap_30[15:0]) +
	( 16'sd 17981) * $signed(input_fmap_31[15:0]) +
	( 15'sd 14165) * $signed(input_fmap_32[15:0]) +
	( 16'sd 25549) * $signed(input_fmap_33[15:0]) +
	( 16'sd 24897) * $signed(input_fmap_34[15:0]) +
	( 15'sd 14566) * $signed(input_fmap_35[15:0]) +
	( 16'sd 24759) * $signed(input_fmap_36[15:0]) +
	( 16'sd 20750) * $signed(input_fmap_37[15:0]) +
	( 14'sd 6213) * $signed(input_fmap_38[15:0]) +
	( 16'sd 26170) * $signed(input_fmap_39[15:0]) +
	( 16'sd 22686) * $signed(input_fmap_40[15:0]) +
	( 16'sd 23738) * $signed(input_fmap_41[15:0]) +
	( 16'sd 25063) * $signed(input_fmap_42[15:0]) +
	( 16'sd 22065) * $signed(input_fmap_43[15:0]) +
	( 16'sd 23611) * $signed(input_fmap_44[15:0]) +
	( 16'sd 23296) * $signed(input_fmap_45[15:0]) +
	( 16'sd 22008) * $signed(input_fmap_46[15:0]) +
	( 16'sd 31423) * $signed(input_fmap_47[15:0]) +
	( 16'sd 30011) * $signed(input_fmap_48[15:0]) +
	( 14'sd 5498) * $signed(input_fmap_49[15:0]) +
	( 16'sd 28620) * $signed(input_fmap_50[15:0]) +
	( 16'sd 26386) * $signed(input_fmap_51[15:0]) +
	( 16'sd 26070) * $signed(input_fmap_52[15:0]) +
	( 15'sd 10775) * $signed(input_fmap_53[15:0]) +
	( 16'sd 23527) * $signed(input_fmap_54[15:0]) +
	( 12'sd 1866) * $signed(input_fmap_55[15:0]) +
	( 16'sd 25901) * $signed(input_fmap_56[15:0]) +
	( 14'sd 4616) * $signed(input_fmap_57[15:0]) +
	( 16'sd 17814) * $signed(input_fmap_58[15:0]) +
	( 16'sd 31465) * $signed(input_fmap_59[15:0]) +
	( 16'sd 28757) * $signed(input_fmap_60[15:0]) +
	( 16'sd 26139) * $signed(input_fmap_61[15:0]) +
	( 15'sd 14521) * $signed(input_fmap_62[15:0]) +
	( 12'sd 1349) * $signed(input_fmap_63[15:0]) +
	( 16'sd 28519) * $signed(input_fmap_64[15:0]) +
	( 15'sd 13249) * $signed(input_fmap_65[15:0]) +
	( 16'sd 22227) * $signed(input_fmap_66[15:0]) +
	( 15'sd 9430) * $signed(input_fmap_67[15:0]) +
	( 15'sd 10161) * $signed(input_fmap_68[15:0]) +
	( 16'sd 19437) * $signed(input_fmap_69[15:0]) +
	( 13'sd 3843) * $signed(input_fmap_70[15:0]) +
	( 16'sd 27498) * $signed(input_fmap_71[15:0]) +
	( 16'sd 18276) * $signed(input_fmap_72[15:0]) +
	( 16'sd 19764) * $signed(input_fmap_73[15:0]) +
	( 13'sd 3479) * $signed(input_fmap_74[15:0]) +
	( 13'sd 2267) * $signed(input_fmap_75[15:0]) +
	( 16'sd 23575) * $signed(input_fmap_76[15:0]) +
	( 16'sd 18900) * $signed(input_fmap_77[15:0]) +
	( 16'sd 18843) * $signed(input_fmap_78[15:0]) +
	( 16'sd 16664) * $signed(input_fmap_79[15:0]) +
	( 15'sd 15130) * $signed(input_fmap_80[15:0]) +
	( 12'sd 1647) * $signed(input_fmap_81[15:0]) +
	( 15'sd 15638) * $signed(input_fmap_82[15:0]) +
	( 15'sd 16050) * $signed(input_fmap_83[15:0]) +
	( 12'sd 1353) * $signed(input_fmap_84[15:0]) +
	( 16'sd 21130) * $signed(input_fmap_85[15:0]) +
	( 16'sd 16843) * $signed(input_fmap_86[15:0]) +
	( 13'sd 3530) * $signed(input_fmap_87[15:0]) +
	( 16'sd 24736) * $signed(input_fmap_88[15:0]) +
	( 16'sd 27137) * $signed(input_fmap_89[15:0]) +
	( 16'sd 21348) * $signed(input_fmap_90[15:0]) +
	( 16'sd 25423) * $signed(input_fmap_91[15:0]) +
	( 16'sd 31933) * $signed(input_fmap_92[15:0]) +
	( 16'sd 21793) * $signed(input_fmap_93[15:0]) +
	( 15'sd 15464) * $signed(input_fmap_94[15:0]) +
	( 14'sd 6850) * $signed(input_fmap_95[15:0]) +
	( 16'sd 32696) * $signed(input_fmap_96[15:0]) +
	( 13'sd 3514) * $signed(input_fmap_97[15:0]) +
	( 16'sd 25639) * $signed(input_fmap_98[15:0]) +
	( 14'sd 4771) * $signed(input_fmap_99[15:0]) +
	( 12'sd 1104) * $signed(input_fmap_100[15:0]) +
	( 14'sd 7174) * $signed(input_fmap_101[15:0]) +
	( 15'sd 8471) * $signed(input_fmap_102[15:0]) +
	( 14'sd 7002) * $signed(input_fmap_103[15:0]) +
	( 14'sd 6279) * $signed(input_fmap_104[15:0]) +
	( 16'sd 31828) * $signed(input_fmap_105[15:0]) +
	( 16'sd 18480) * $signed(input_fmap_106[15:0]) +
	( 15'sd 14152) * $signed(input_fmap_107[15:0]) +
	( 16'sd 18566) * $signed(input_fmap_108[15:0]) +
	( 16'sd 29151) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22143) * $signed(input_fmap_110[15:0]) +
	( 16'sd 29530) * $signed(input_fmap_111[15:0]) +
	( 15'sd 13081) * $signed(input_fmap_112[15:0]) +
	( 16'sd 18552) * $signed(input_fmap_113[15:0]) +
	( 16'sd 18968) * $signed(input_fmap_114[15:0]) +
	( 14'sd 7388) * $signed(input_fmap_115[15:0]) +
	( 14'sd 5719) * $signed(input_fmap_116[15:0]) +
	( 16'sd 20163) * $signed(input_fmap_117[15:0]) +
	( 16'sd 28713) * $signed(input_fmap_118[15:0]) +
	( 16'sd 16613) * $signed(input_fmap_119[15:0]) +
	( 15'sd 9779) * $signed(input_fmap_120[15:0]) +
	( 16'sd 30248) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9726) * $signed(input_fmap_122[15:0]) +
	( 16'sd 17282) * $signed(input_fmap_123[15:0]) +
	( 16'sd 19920) * $signed(input_fmap_124[15:0]) +
	( 14'sd 4520) * $signed(input_fmap_125[15:0]) +
	( 15'sd 12722) * $signed(input_fmap_126[15:0]) +
	( 11'sd 761) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 16'sd 18553) * $signed(input_fmap_0[15:0]) +
	( 15'sd 11335) * $signed(input_fmap_1[15:0]) +
	( 15'sd 15745) * $signed(input_fmap_2[15:0]) +
	( 16'sd 18047) * $signed(input_fmap_3[15:0]) +
	( 13'sd 2759) * $signed(input_fmap_4[15:0]) +
	( 14'sd 6833) * $signed(input_fmap_5[15:0]) +
	( 15'sd 14433) * $signed(input_fmap_6[15:0]) +
	( 16'sd 16631) * $signed(input_fmap_7[15:0]) +
	( 16'sd 20751) * $signed(input_fmap_8[15:0]) +
	( 16'sd 26182) * $signed(input_fmap_9[15:0]) +
	( 13'sd 3359) * $signed(input_fmap_10[15:0]) +
	( 16'sd 18614) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20263) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24319) * $signed(input_fmap_13[15:0]) +
	( 16'sd 32455) * $signed(input_fmap_14[15:0]) +
	( 16'sd 17937) * $signed(input_fmap_15[15:0]) +
	( 15'sd 12488) * $signed(input_fmap_16[15:0]) +
	( 16'sd 16885) * $signed(input_fmap_17[15:0]) +
	( 16'sd 23478) * $signed(input_fmap_18[15:0]) +
	( 16'sd 28802) * $signed(input_fmap_19[15:0]) +
	( 16'sd 21033) * $signed(input_fmap_20[15:0]) +
	( 16'sd 20855) * $signed(input_fmap_21[15:0]) +
	( 16'sd 29079) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28895) * $signed(input_fmap_23[15:0]) +
	( 16'sd 16490) * $signed(input_fmap_24[15:0]) +
	( 15'sd 15278) * $signed(input_fmap_25[15:0]) +
	( 15'sd 14724) * $signed(input_fmap_26[15:0]) +
	( 14'sd 4778) * $signed(input_fmap_27[15:0]) +
	( 15'sd 15821) * $signed(input_fmap_28[15:0]) +
	( 15'sd 13149) * $signed(input_fmap_29[15:0]) +
	( 15'sd 12940) * $signed(input_fmap_30[15:0]) +
	( 15'sd 8521) * $signed(input_fmap_31[15:0]) +
	( 16'sd 17464) * $signed(input_fmap_32[15:0]) +
	( 12'sd 1666) * $signed(input_fmap_33[15:0]) +
	( 16'sd 16501) * $signed(input_fmap_34[15:0]) +
	( 15'sd 12771) * $signed(input_fmap_35[15:0]) +
	( 16'sd 16681) * $signed(input_fmap_36[15:0]) +
	( 16'sd 28897) * $signed(input_fmap_37[15:0]) +
	( 15'sd 10933) * $signed(input_fmap_38[15:0]) +
	( 16'sd 29173) * $signed(input_fmap_39[15:0]) +
	( 16'sd 22238) * $signed(input_fmap_40[15:0]) +
	( 16'sd 19836) * $signed(input_fmap_41[15:0]) +
	( 16'sd 16823) * $signed(input_fmap_42[15:0]) +
	( 16'sd 26113) * $signed(input_fmap_43[15:0]) +
	( 16'sd 27267) * $signed(input_fmap_44[15:0]) +
	( 15'sd 13686) * $signed(input_fmap_45[15:0]) +
	( 13'sd 3149) * $signed(input_fmap_46[15:0]) +
	( 14'sd 4342) * $signed(input_fmap_47[15:0]) +
	( 14'sd 7754) * $signed(input_fmap_48[15:0]) +
	( 16'sd 23370) * $signed(input_fmap_49[15:0]) +
	( 13'sd 2178) * $signed(input_fmap_50[15:0]) +
	( 16'sd 24696) * $signed(input_fmap_51[15:0]) +
	( 16'sd 26457) * $signed(input_fmap_52[15:0]) +
	( 16'sd 30843) * $signed(input_fmap_53[15:0]) +
	( 15'sd 13490) * $signed(input_fmap_54[15:0]) +
	( 16'sd 17121) * $signed(input_fmap_55[15:0]) +
	( 13'sd 2925) * $signed(input_fmap_56[15:0]) +
	( 14'sd 8008) * $signed(input_fmap_57[15:0]) +
	( 16'sd 22911) * $signed(input_fmap_58[15:0]) +
	( 16'sd 25480) * $signed(input_fmap_59[15:0]) +
	( 16'sd 26578) * $signed(input_fmap_60[15:0]) +
	( 16'sd 28368) * $signed(input_fmap_61[15:0]) +
	( 16'sd 21129) * $signed(input_fmap_62[15:0]) +
	( 15'sd 15300) * $signed(input_fmap_63[15:0]) +
	( 14'sd 4343) * $signed(input_fmap_64[15:0]) +
	( 16'sd 32522) * $signed(input_fmap_65[15:0]) +
	( 16'sd 26729) * $signed(input_fmap_66[15:0]) +
	( 14'sd 7642) * $signed(input_fmap_67[15:0]) +
	( 16'sd 22808) * $signed(input_fmap_68[15:0]) +
	( 16'sd 27918) * $signed(input_fmap_69[15:0]) +
	( 15'sd 9639) * $signed(input_fmap_70[15:0]) +
	( 16'sd 19817) * $signed(input_fmap_71[15:0]) +
	( 13'sd 3274) * $signed(input_fmap_72[15:0]) +
	( 15'sd 11018) * $signed(input_fmap_73[15:0]) +
	( 16'sd 31227) * $signed(input_fmap_74[15:0]) +
	( 15'sd 14944) * $signed(input_fmap_75[15:0]) +
	( 16'sd 25257) * $signed(input_fmap_76[15:0]) +
	( 15'sd 13618) * $signed(input_fmap_77[15:0]) +
	( 16'sd 23700) * $signed(input_fmap_78[15:0]) +
	( 12'sd 1608) * $signed(input_fmap_79[15:0]) +
	( 15'sd 15984) * $signed(input_fmap_80[15:0]) +
	( 16'sd 21527) * $signed(input_fmap_81[15:0]) +
	( 16'sd 32198) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25627) * $signed(input_fmap_83[15:0]) +
	( 15'sd 12395) * $signed(input_fmap_84[15:0]) +
	( 9'sd 232) * $signed(input_fmap_85[15:0]) +
	( 16'sd 27430) * $signed(input_fmap_86[15:0]) +
	( 13'sd 3422) * $signed(input_fmap_87[15:0]) +
	( 13'sd 3644) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5870) * $signed(input_fmap_89[15:0]) +
	( 16'sd 21209) * $signed(input_fmap_90[15:0]) +
	( 16'sd 20467) * $signed(input_fmap_91[15:0]) +
	( 14'sd 6157) * $signed(input_fmap_92[15:0]) +
	( 15'sd 9798) * $signed(input_fmap_93[15:0]) +
	( 15'sd 13913) * $signed(input_fmap_94[15:0]) +
	( 16'sd 21921) * $signed(input_fmap_95[15:0]) +
	( 16'sd 17832) * $signed(input_fmap_96[15:0]) +
	( 16'sd 18664) * $signed(input_fmap_97[15:0]) +
	( 16'sd 17734) * $signed(input_fmap_98[15:0]) +
	( 15'sd 14523) * $signed(input_fmap_99[15:0]) +
	( 16'sd 21608) * $signed(input_fmap_100[15:0]) +
	( 15'sd 10270) * $signed(input_fmap_101[15:0]) +
	( 16'sd 25678) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28430) * $signed(input_fmap_103[15:0]) +
	( 16'sd 32516) * $signed(input_fmap_104[15:0]) +
	( 14'sd 7485) * $signed(input_fmap_105[15:0]) +
	( 16'sd 20955) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27636) * $signed(input_fmap_107[15:0]) +
	( 15'sd 9199) * $signed(input_fmap_108[15:0]) +
	( 16'sd 17759) * $signed(input_fmap_109[15:0]) +
	( 16'sd 23722) * $signed(input_fmap_110[15:0]) +
	( 16'sd 21338) * $signed(input_fmap_111[15:0]) +
	( 16'sd 24710) * $signed(input_fmap_112[15:0]) +
	( 14'sd 5316) * $signed(input_fmap_113[15:0]) +
	( 15'sd 14026) * $signed(input_fmap_114[15:0]) +
	( 14'sd 7202) * $signed(input_fmap_115[15:0]) +
	( 16'sd 27659) * $signed(input_fmap_116[15:0]) +
	( 16'sd 28410) * $signed(input_fmap_117[15:0]) +
	( 12'sd 1328) * $signed(input_fmap_118[15:0]) +
	( 16'sd 28287) * $signed(input_fmap_119[15:0]) +
	( 15'sd 11313) * $signed(input_fmap_120[15:0]) +
	( 16'sd 23812) * $signed(input_fmap_121[15:0]) +
	( 16'sd 25029) * $signed(input_fmap_122[15:0]) +
	( 15'sd 10608) * $signed(input_fmap_123[15:0]) +
	( 12'sd 1460) * $signed(input_fmap_124[15:0]) +
	( 15'sd 11400) * $signed(input_fmap_125[15:0]) +
	( 12'sd 1795) * $signed(input_fmap_126[15:0]) +
	( 15'sd 9115) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 16'sd 21669) * $signed(input_fmap_0[15:0]) +
	( 15'sd 13425) * $signed(input_fmap_1[15:0]) +
	( 15'sd 10424) * $signed(input_fmap_2[15:0]) +
	( 16'sd 20493) * $signed(input_fmap_3[15:0]) +
	( 15'sd 13901) * $signed(input_fmap_4[15:0]) +
	( 15'sd 9935) * $signed(input_fmap_5[15:0]) +
	( 16'sd 22242) * $signed(input_fmap_6[15:0]) +
	( 16'sd 21866) * $signed(input_fmap_7[15:0]) +
	( 15'sd 9016) * $signed(input_fmap_8[15:0]) +
	( 16'sd 16623) * $signed(input_fmap_9[15:0]) +
	( 16'sd 27241) * $signed(input_fmap_10[15:0]) +
	( 14'sd 5309) * $signed(input_fmap_11[15:0]) +
	( 15'sd 15425) * $signed(input_fmap_12[15:0]) +
	( 15'sd 14077) * $signed(input_fmap_13[15:0]) +
	( 16'sd 31816) * $signed(input_fmap_14[15:0]) +
	( 16'sd 22414) * $signed(input_fmap_15[15:0]) +
	( 13'sd 3481) * $signed(input_fmap_16[15:0]) +
	( 15'sd 14209) * $signed(input_fmap_17[15:0]) +
	( 12'sd 1306) * $signed(input_fmap_18[15:0]) +
	( 14'sd 7433) * $signed(input_fmap_19[15:0]) +
	( 16'sd 20782) * $signed(input_fmap_20[15:0]) +
	( 16'sd 29746) * $signed(input_fmap_21[15:0]) +
	( 16'sd 27393) * $signed(input_fmap_22[15:0]) +
	( 16'sd 29708) * $signed(input_fmap_23[15:0]) +
	( 16'sd 21632) * $signed(input_fmap_24[15:0]) +
	( 16'sd 24760) * $signed(input_fmap_25[15:0]) +
	( 14'sd 4727) * $signed(input_fmap_26[15:0]) +
	( 16'sd 18464) * $signed(input_fmap_27[15:0]) +
	( 13'sd 2636) * $signed(input_fmap_28[15:0]) +
	( 16'sd 27042) * $signed(input_fmap_29[15:0]) +
	( 16'sd 16965) * $signed(input_fmap_30[15:0]) +
	( 16'sd 24930) * $signed(input_fmap_31[15:0]) +
	( 14'sd 4110) * $signed(input_fmap_32[15:0]) +
	( 16'sd 28516) * $signed(input_fmap_33[15:0]) +
	( 16'sd 24949) * $signed(input_fmap_34[15:0]) +
	( 16'sd 22158) * $signed(input_fmap_35[15:0]) +
	( 16'sd 25574) * $signed(input_fmap_36[15:0]) +
	( 16'sd 31867) * $signed(input_fmap_37[15:0]) +
	( 15'sd 9407) * $signed(input_fmap_38[15:0]) +
	( 15'sd 9709) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6271) * $signed(input_fmap_40[15:0]) +
	( 16'sd 29004) * $signed(input_fmap_41[15:0]) +
	( 16'sd 27801) * $signed(input_fmap_42[15:0]) +
	( 16'sd 31807) * $signed(input_fmap_43[15:0]) +
	( 16'sd 21823) * $signed(input_fmap_44[15:0]) +
	( 16'sd 28418) * $signed(input_fmap_45[15:0]) +
	( 16'sd 17065) * $signed(input_fmap_46[15:0]) +
	( 11'sd 869) * $signed(input_fmap_47[15:0]) +
	( 10'sd 338) * $signed(input_fmap_48[15:0]) +
	( 16'sd 29119) * $signed(input_fmap_49[15:0]) +
	( 14'sd 4684) * $signed(input_fmap_50[15:0]) +
	( 15'sd 13323) * $signed(input_fmap_51[15:0]) +
	( 16'sd 24134) * $signed(input_fmap_52[15:0]) +
	( 15'sd 12849) * $signed(input_fmap_53[15:0]) +
	( 15'sd 12415) * $signed(input_fmap_54[15:0]) +
	( 16'sd 31333) * $signed(input_fmap_55[15:0]) +
	( 14'sd 6976) * $signed(input_fmap_56[15:0]) +
	( 15'sd 9202) * $signed(input_fmap_57[15:0]) +
	( 16'sd 28302) * $signed(input_fmap_58[15:0]) +
	( 15'sd 12406) * $signed(input_fmap_59[15:0]) +
	( 15'sd 11225) * $signed(input_fmap_60[15:0]) +
	( 14'sd 4899) * $signed(input_fmap_61[15:0]) +
	( 15'sd 13178) * $signed(input_fmap_62[15:0]) +
	( 15'sd 9262) * $signed(input_fmap_63[15:0]) +
	( 15'sd 15675) * $signed(input_fmap_64[15:0]) +
	( 16'sd 25082) * $signed(input_fmap_65[15:0]) +
	( 16'sd 22723) * $signed(input_fmap_66[15:0]) +
	( 16'sd 20744) * $signed(input_fmap_67[15:0]) +
	( 16'sd 31543) * $signed(input_fmap_68[15:0]) +
	( 16'sd 19388) * $signed(input_fmap_69[15:0]) +
	( 13'sd 2466) * $signed(input_fmap_70[15:0]) +
	( 14'sd 7370) * $signed(input_fmap_71[15:0]) +
	( 15'sd 12977) * $signed(input_fmap_72[15:0]) +
	( 16'sd 29734) * $signed(input_fmap_73[15:0]) +
	( 15'sd 12505) * $signed(input_fmap_74[15:0]) +
	( 11'sd 759) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19385) * $signed(input_fmap_76[15:0]) +
	( 16'sd 31448) * $signed(input_fmap_77[15:0]) +
	( 14'sd 7078) * $signed(input_fmap_78[15:0]) +
	( 16'sd 27460) * $signed(input_fmap_79[15:0]) +
	( 16'sd 20670) * $signed(input_fmap_80[15:0]) +
	( 15'sd 15719) * $signed(input_fmap_81[15:0]) +
	( 13'sd 2502) * $signed(input_fmap_82[15:0]) +
	( 11'sd 974) * $signed(input_fmap_83[15:0]) +
	( 14'sd 8105) * $signed(input_fmap_84[15:0]) +
	( 16'sd 19219) * $signed(input_fmap_85[15:0]) +
	( 16'sd 17326) * $signed(input_fmap_86[15:0]) +
	( 16'sd 22336) * $signed(input_fmap_87[15:0]) +
	( 12'sd 1514) * $signed(input_fmap_88[15:0]) +
	( 16'sd 29043) * $signed(input_fmap_89[15:0]) +
	( 15'sd 10095) * $signed(input_fmap_90[15:0]) +
	( 14'sd 4114) * $signed(input_fmap_91[15:0]) +
	( 12'sd 1555) * $signed(input_fmap_92[15:0]) +
	( 15'sd 15561) * $signed(input_fmap_93[15:0]) +
	( 11'sd 984) * $signed(input_fmap_94[15:0]) +
	( 15'sd 10927) * $signed(input_fmap_95[15:0]) +
	( 14'sd 6355) * $signed(input_fmap_96[15:0]) +
	( 16'sd 17933) * $signed(input_fmap_97[15:0]) +
	( 16'sd 27057) * $signed(input_fmap_98[15:0]) +
	( 13'sd 3623) * $signed(input_fmap_99[15:0]) +
	( 15'sd 16187) * $signed(input_fmap_100[15:0]) +
	( 16'sd 23934) * $signed(input_fmap_101[15:0]) +
	( 16'sd 17309) * $signed(input_fmap_102[15:0]) +
	( 16'sd 30544) * $signed(input_fmap_103[15:0]) +
	( 15'sd 10677) * $signed(input_fmap_104[15:0]) +
	( 16'sd 17206) * $signed(input_fmap_105[15:0]) +
	( 15'sd 14716) * $signed(input_fmap_106[15:0]) +
	( 15'sd 12843) * $signed(input_fmap_107[15:0]) +
	( 14'sd 6292) * $signed(input_fmap_108[15:0]) +
	( 16'sd 25219) * $signed(input_fmap_109[15:0]) +
	( 14'sd 6101) * $signed(input_fmap_110[15:0]) +
	( 16'sd 26630) * $signed(input_fmap_111[15:0]) +
	( 13'sd 3258) * $signed(input_fmap_112[15:0]) +
	( 15'sd 10583) * $signed(input_fmap_113[15:0]) +
	( 15'sd 15234) * $signed(input_fmap_114[15:0]) +
	( 15'sd 9371) * $signed(input_fmap_115[15:0]) +
	( 13'sd 2502) * $signed(input_fmap_116[15:0]) +
	( 13'sd 2327) * $signed(input_fmap_117[15:0]) +
	( 14'sd 6522) * $signed(input_fmap_118[15:0]) +
	( 15'sd 12753) * $signed(input_fmap_119[15:0]) +
	( 16'sd 16627) * $signed(input_fmap_120[15:0]) +
	( 16'sd 23520) * $signed(input_fmap_121[15:0]) +
	( 16'sd 18289) * $signed(input_fmap_122[15:0]) +
	( 16'sd 32607) * $signed(input_fmap_123[15:0]) +
	( 15'sd 15449) * $signed(input_fmap_124[15:0]) +
	( 16'sd 25222) * $signed(input_fmap_125[15:0]) +
	( 15'sd 10380) * $signed(input_fmap_126[15:0]) +
	( 16'sd 28978) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 15'sd 15405) * $signed(input_fmap_0[15:0]) +
	( 16'sd 25372) * $signed(input_fmap_1[15:0]) +
	( 16'sd 30284) * $signed(input_fmap_2[15:0]) +
	( 16'sd 17972) * $signed(input_fmap_3[15:0]) +
	( 16'sd 22691) * $signed(input_fmap_4[15:0]) +
	( 16'sd 28080) * $signed(input_fmap_5[15:0]) +
	( 15'sd 9899) * $signed(input_fmap_6[15:0]) +
	( 16'sd 23278) * $signed(input_fmap_7[15:0]) +
	( 14'sd 6499) * $signed(input_fmap_8[15:0]) +
	( 15'sd 9314) * $signed(input_fmap_9[15:0]) +
	( 16'sd 17330) * $signed(input_fmap_10[15:0]) +
	( 16'sd 28368) * $signed(input_fmap_11[15:0]) +
	( 16'sd 19633) * $signed(input_fmap_12[15:0]) +
	( 16'sd 23431) * $signed(input_fmap_13[15:0]) +
	( 14'sd 7802) * $signed(input_fmap_14[15:0]) +
	( 16'sd 25538) * $signed(input_fmap_15[15:0]) +
	( 16'sd 30979) * $signed(input_fmap_16[15:0]) +
	( 16'sd 30363) * $signed(input_fmap_17[15:0]) +
	( 16'sd 31409) * $signed(input_fmap_18[15:0]) +
	( 15'sd 12789) * $signed(input_fmap_19[15:0]) +
	( 13'sd 2385) * $signed(input_fmap_20[15:0]) +
	( 16'sd 21558) * $signed(input_fmap_21[15:0]) +
	( 15'sd 11503) * $signed(input_fmap_22[15:0]) +
	( 14'sd 5373) * $signed(input_fmap_23[15:0]) +
	( 10'sd 422) * $signed(input_fmap_24[15:0]) +
	( 16'sd 23337) * $signed(input_fmap_25[15:0]) +
	( 16'sd 21611) * $signed(input_fmap_26[15:0]) +
	( 14'sd 6003) * $signed(input_fmap_27[15:0]) +
	( 16'sd 22372) * $signed(input_fmap_28[15:0]) +
	( 14'sd 6931) * $signed(input_fmap_29[15:0]) +
	( 15'sd 9741) * $signed(input_fmap_30[15:0]) +
	( 16'sd 32412) * $signed(input_fmap_31[15:0]) +
	( 16'sd 24977) * $signed(input_fmap_32[15:0]) +
	( 14'sd 6172) * $signed(input_fmap_33[15:0]) +
	( 15'sd 15364) * $signed(input_fmap_34[15:0]) +
	( 16'sd 23289) * $signed(input_fmap_35[15:0]) +
	( 16'sd 22213) * $signed(input_fmap_36[15:0]) +
	( 15'sd 10886) * $signed(input_fmap_37[15:0]) +
	( 11'sd 741) * $signed(input_fmap_38[15:0]) +
	( 14'sd 7636) * $signed(input_fmap_39[15:0]) +
	( 14'sd 4383) * $signed(input_fmap_40[15:0]) +
	( 16'sd 31365) * $signed(input_fmap_41[15:0]) +
	( 16'sd 16753) * $signed(input_fmap_42[15:0]) +
	( 14'sd 6453) * $signed(input_fmap_43[15:0]) +
	( 15'sd 14693) * $signed(input_fmap_44[15:0]) +
	( 15'sd 10388) * $signed(input_fmap_45[15:0]) +
	( 16'sd 31005) * $signed(input_fmap_46[15:0]) +
	( 14'sd 4298) * $signed(input_fmap_47[15:0]) +
	( 16'sd 28410) * $signed(input_fmap_48[15:0]) +
	( 16'sd 22936) * $signed(input_fmap_49[15:0]) +
	( 15'sd 11469) * $signed(input_fmap_50[15:0]) +
	( 16'sd 25986) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19004) * $signed(input_fmap_52[15:0]) +
	( 11'sd 834) * $signed(input_fmap_53[15:0]) +
	( 16'sd 30445) * $signed(input_fmap_54[15:0]) +
	( 15'sd 11234) * $signed(input_fmap_55[15:0]) +
	( 16'sd 22040) * $signed(input_fmap_56[15:0]) +
	( 13'sd 2740) * $signed(input_fmap_57[15:0]) +
	( 16'sd 28914) * $signed(input_fmap_58[15:0]) +
	( 16'sd 19895) * $signed(input_fmap_59[15:0]) +
	( 15'sd 11137) * $signed(input_fmap_60[15:0]) +
	( 16'sd 20949) * $signed(input_fmap_61[15:0]) +
	( 16'sd 31581) * $signed(input_fmap_62[15:0]) +
	( 16'sd 29536) * $signed(input_fmap_63[15:0]) +
	( 12'sd 1318) * $signed(input_fmap_64[15:0]) +
	( 15'sd 16168) * $signed(input_fmap_65[15:0]) +
	( 15'sd 10373) * $signed(input_fmap_66[15:0]) +
	( 16'sd 17462) * $signed(input_fmap_67[15:0]) +
	( 16'sd 22973) * $signed(input_fmap_68[15:0]) +
	( 16'sd 21650) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31688) * $signed(input_fmap_70[15:0]) +
	( 16'sd 29562) * $signed(input_fmap_71[15:0]) +
	( 15'sd 14299) * $signed(input_fmap_72[15:0]) +
	( 16'sd 21313) * $signed(input_fmap_73[15:0]) +
	( 13'sd 3861) * $signed(input_fmap_74[15:0]) +
	( 14'sd 6694) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19153) * $signed(input_fmap_76[15:0]) +
	( 16'sd 30238) * $signed(input_fmap_77[15:0]) +
	( 16'sd 29726) * $signed(input_fmap_78[15:0]) +
	( 16'sd 18233) * $signed(input_fmap_79[15:0]) +
	( 14'sd 7087) * $signed(input_fmap_80[15:0]) +
	( 14'sd 7454) * $signed(input_fmap_81[15:0]) +
	( 14'sd 6689) * $signed(input_fmap_82[15:0]) +
	( 15'sd 8398) * $signed(input_fmap_83[15:0]) +
	( 16'sd 17880) * $signed(input_fmap_84[15:0]) +
	( 16'sd 26481) * $signed(input_fmap_85[15:0]) +
	( 16'sd 16612) * $signed(input_fmap_86[15:0]) +
	( 16'sd 18691) * $signed(input_fmap_87[15:0]) +
	( 16'sd 24443) * $signed(input_fmap_88[15:0]) +
	( 16'sd 31358) * $signed(input_fmap_89[15:0]) +
	( 16'sd 17003) * $signed(input_fmap_90[15:0]) +
	( 15'sd 10512) * $signed(input_fmap_91[15:0]) +
	( 15'sd 8502) * $signed(input_fmap_92[15:0]) +
	( 16'sd 16702) * $signed(input_fmap_93[15:0]) +
	( 15'sd 11857) * $signed(input_fmap_94[15:0]) +
	( 16'sd 28292) * $signed(input_fmap_95[15:0]) +
	( 16'sd 28060) * $signed(input_fmap_96[15:0]) +
	( 16'sd 17736) * $signed(input_fmap_97[15:0]) +
	( 16'sd 24269) * $signed(input_fmap_98[15:0]) +
	( 16'sd 29923) * $signed(input_fmap_99[15:0]) +
	( 14'sd 5681) * $signed(input_fmap_100[15:0]) +
	( 16'sd 24170) * $signed(input_fmap_101[15:0]) +
	( 16'sd 19600) * $signed(input_fmap_102[15:0]) +
	( 15'sd 11305) * $signed(input_fmap_103[15:0]) +
	( 16'sd 24847) * $signed(input_fmap_104[15:0]) +
	( 16'sd 22832) * $signed(input_fmap_105[15:0]) +
	( 15'sd 9666) * $signed(input_fmap_106[15:0]) +
	( 15'sd 14400) * $signed(input_fmap_107[15:0]) +
	( 16'sd 22702) * $signed(input_fmap_108[15:0]) +
	( 15'sd 15086) * $signed(input_fmap_109[15:0]) +
	( 15'sd 8577) * $signed(input_fmap_110[15:0]) +
	( 16'sd 29262) * $signed(input_fmap_111[15:0]) +
	( 16'sd 21959) * $signed(input_fmap_112[15:0]) +
	( 16'sd 23145) * $signed(input_fmap_113[15:0]) +
	( 15'sd 8228) * $signed(input_fmap_114[15:0]) +
	( 14'sd 8176) * $signed(input_fmap_115[15:0]) +
	( 14'sd 4275) * $signed(input_fmap_116[15:0]) +
	( 15'sd 9917) * $signed(input_fmap_117[15:0]) +
	( 16'sd 32429) * $signed(input_fmap_118[15:0]) +
	( 16'sd 31634) * $signed(input_fmap_119[15:0]) +
	( 15'sd 13569) * $signed(input_fmap_120[15:0]) +
	( 12'sd 1083) * $signed(input_fmap_121[15:0]) +
	( 14'sd 4530) * $signed(input_fmap_122[15:0]) +
	( 16'sd 18365) * $signed(input_fmap_123[15:0]) +
	( 11'sd 970) * $signed(input_fmap_124[15:0]) +
	( 15'sd 10714) * $signed(input_fmap_125[15:0]) +
	( 16'sd 25441) * $signed(input_fmap_126[15:0]) +
	( 13'sd 2851) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 16'sd 25610) * $signed(input_fmap_0[15:0]) +
	( 13'sd 2549) * $signed(input_fmap_1[15:0]) +
	( 12'sd 1580) * $signed(input_fmap_2[15:0]) +
	( 16'sd 19489) * $signed(input_fmap_3[15:0]) +
	( 14'sd 5866) * $signed(input_fmap_4[15:0]) +
	( 15'sd 10726) * $signed(input_fmap_5[15:0]) +
	( 15'sd 9099) * $signed(input_fmap_6[15:0]) +
	( 15'sd 9058) * $signed(input_fmap_7[15:0]) +
	( 15'sd 9050) * $signed(input_fmap_8[15:0]) +
	( 15'sd 12172) * $signed(input_fmap_9[15:0]) +
	( 16'sd 19410) * $signed(input_fmap_10[15:0]) +
	( 16'sd 18203) * $signed(input_fmap_11[15:0]) +
	( 16'sd 19331) * $signed(input_fmap_12[15:0]) +
	( 16'sd 18255) * $signed(input_fmap_13[15:0]) +
	( 16'sd 21320) * $signed(input_fmap_14[15:0]) +
	( 16'sd 29865) * $signed(input_fmap_15[15:0]) +
	( 16'sd 22485) * $signed(input_fmap_16[15:0]) +
	( 14'sd 7789) * $signed(input_fmap_17[15:0]) +
	( 15'sd 10027) * $signed(input_fmap_18[15:0]) +
	( 16'sd 24311) * $signed(input_fmap_19[15:0]) +
	( 16'sd 22845) * $signed(input_fmap_20[15:0]) +
	( 16'sd 26168) * $signed(input_fmap_21[15:0]) +
	( 15'sd 9799) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24182) * $signed(input_fmap_23[15:0]) +
	( 14'sd 5497) * $signed(input_fmap_24[15:0]) +
	( 16'sd 30431) * $signed(input_fmap_25[15:0]) +
	( 14'sd 7842) * $signed(input_fmap_26[15:0]) +
	( 14'sd 5031) * $signed(input_fmap_27[15:0]) +
	( 16'sd 19082) * $signed(input_fmap_28[15:0]) +
	( 15'sd 15667) * $signed(input_fmap_29[15:0]) +
	( 16'sd 26826) * $signed(input_fmap_30[15:0]) +
	( 9'sd 241) * $signed(input_fmap_31[15:0]) +
	( 15'sd 11956) * $signed(input_fmap_32[15:0]) +
	( 16'sd 18196) * $signed(input_fmap_33[15:0]) +
	( 16'sd 30674) * $signed(input_fmap_34[15:0]) +
	( 16'sd 20933) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11616) * $signed(input_fmap_36[15:0]) +
	( 13'sd 3798) * $signed(input_fmap_37[15:0]) +
	( 12'sd 1049) * $signed(input_fmap_38[15:0]) +
	( 16'sd 26372) * $signed(input_fmap_39[15:0]) +
	( 14'sd 7665) * $signed(input_fmap_40[15:0]) +
	( 15'sd 11236) * $signed(input_fmap_41[15:0]) +
	( 15'sd 14056) * $signed(input_fmap_42[15:0]) +
	( 16'sd 31482) * $signed(input_fmap_43[15:0]) +
	( 15'sd 9592) * $signed(input_fmap_44[15:0]) +
	( 16'sd 19418) * $signed(input_fmap_45[15:0]) +
	( 16'sd 16625) * $signed(input_fmap_46[15:0]) +
	( 16'sd 21185) * $signed(input_fmap_47[15:0]) +
	( 16'sd 25434) * $signed(input_fmap_48[15:0]) +
	( 15'sd 11104) * $signed(input_fmap_49[15:0]) +
	( 16'sd 21664) * $signed(input_fmap_50[15:0]) +
	( 15'sd 8654) * $signed(input_fmap_51[15:0]) +
	( 16'sd 23997) * $signed(input_fmap_52[15:0]) +
	( 16'sd 18277) * $signed(input_fmap_53[15:0]) +
	( 16'sd 22360) * $signed(input_fmap_54[15:0]) +
	( 15'sd 8651) * $signed(input_fmap_55[15:0]) +
	( 16'sd 17706) * $signed(input_fmap_56[15:0]) +
	( 16'sd 31445) * $signed(input_fmap_57[15:0]) +
	( 13'sd 4012) * $signed(input_fmap_58[15:0]) +
	( 11'sd 981) * $signed(input_fmap_59[15:0]) +
	( 15'sd 14538) * $signed(input_fmap_60[15:0]) +
	( 14'sd 8088) * $signed(input_fmap_61[15:0]) +
	( 16'sd 22635) * $signed(input_fmap_62[15:0]) +
	( 15'sd 9777) * $signed(input_fmap_63[15:0]) +
	( 16'sd 19577) * $signed(input_fmap_64[15:0]) +
	( 16'sd 23712) * $signed(input_fmap_65[15:0]) +
	( 16'sd 24361) * $signed(input_fmap_66[15:0]) +
	( 11'sd 873) * $signed(input_fmap_67[15:0]) +
	( 10'sd 264) * $signed(input_fmap_68[15:0]) +
	( 15'sd 14027) * $signed(input_fmap_69[15:0]) +
	( 16'sd 19551) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31207) * $signed(input_fmap_71[15:0]) +
	( 16'sd 28189) * $signed(input_fmap_72[15:0]) +
	( 10'sd 333) * $signed(input_fmap_73[15:0]) +
	( 16'sd 29430) * $signed(input_fmap_74[15:0]) +
	( 16'sd 25930) * $signed(input_fmap_75[15:0]) +
	( 15'sd 9091) * $signed(input_fmap_76[15:0]) +
	( 16'sd 22640) * $signed(input_fmap_77[15:0]) +
	( 15'sd 10496) * $signed(input_fmap_78[15:0]) +
	( 16'sd 30269) * $signed(input_fmap_79[15:0]) +
	( 15'sd 9273) * $signed(input_fmap_80[15:0]) +
	( 15'sd 11635) * $signed(input_fmap_81[15:0]) +
	( 15'sd 12774) * $signed(input_fmap_82[15:0]) +
	( 15'sd 13787) * $signed(input_fmap_83[15:0]) +
	( 16'sd 20258) * $signed(input_fmap_84[15:0]) +
	( 16'sd 19551) * $signed(input_fmap_85[15:0]) +
	( 15'sd 11074) * $signed(input_fmap_86[15:0]) +
	( 14'sd 7583) * $signed(input_fmap_87[15:0]) +
	( 16'sd 25059) * $signed(input_fmap_88[15:0]) +
	( 16'sd 24443) * $signed(input_fmap_89[15:0]) +
	( 15'sd 12865) * $signed(input_fmap_90[15:0]) +
	( 16'sd 29495) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25208) * $signed(input_fmap_92[15:0]) +
	( 16'sd 30332) * $signed(input_fmap_93[15:0]) +
	( 16'sd 21461) * $signed(input_fmap_94[15:0]) +
	( 14'sd 8143) * $signed(input_fmap_95[15:0]) +
	( 16'sd 28557) * $signed(input_fmap_96[15:0]) +
	( 15'sd 16320) * $signed(input_fmap_97[15:0]) +
	( 16'sd 29140) * $signed(input_fmap_98[15:0]) +
	( 16'sd 27201) * $signed(input_fmap_99[15:0]) +
	( 13'sd 3931) * $signed(input_fmap_100[15:0]) +
	( 16'sd 17122) * $signed(input_fmap_101[15:0]) +
	( 15'sd 10625) * $signed(input_fmap_102[15:0]) +
	( 16'sd 21167) * $signed(input_fmap_103[15:0]) +
	( 16'sd 20767) * $signed(input_fmap_104[15:0]) +
	( 16'sd 20380) * $signed(input_fmap_105[15:0]) +
	( 16'sd 29219) * $signed(input_fmap_106[15:0]) +
	( 13'sd 3299) * $signed(input_fmap_107[15:0]) +
	( 14'sd 4617) * $signed(input_fmap_108[15:0]) +
	( 16'sd 18372) * $signed(input_fmap_109[15:0]) +
	( 13'sd 4026) * $signed(input_fmap_110[15:0]) +
	( 15'sd 15706) * $signed(input_fmap_111[15:0]) +
	( 15'sd 9035) * $signed(input_fmap_112[15:0]) +
	( 12'sd 1465) * $signed(input_fmap_113[15:0]) +
	( 16'sd 31421) * $signed(input_fmap_114[15:0]) +
	( 15'sd 15170) * $signed(input_fmap_115[15:0]) +
	( 16'sd 19585) * $signed(input_fmap_116[15:0]) +
	( 14'sd 5582) * $signed(input_fmap_117[15:0]) +
	( 16'sd 17843) * $signed(input_fmap_118[15:0]) +
	( 16'sd 26560) * $signed(input_fmap_119[15:0]) +
	( 16'sd 16658) * $signed(input_fmap_120[15:0]) +
	( 13'sd 2260) * $signed(input_fmap_121[15:0]) +
	( 16'sd 27607) * $signed(input_fmap_122[15:0]) +
	( 16'sd 32403) * $signed(input_fmap_123[15:0]) +
	( 16'sd 17095) * $signed(input_fmap_124[15:0]) +
	( 15'sd 13170) * $signed(input_fmap_125[15:0]) +
	( 15'sd 10829) * $signed(input_fmap_126[15:0]) +
	( 15'sd 14288) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 16'sd 27607) * $signed(input_fmap_0[15:0]) +
	( 15'sd 12645) * $signed(input_fmap_1[15:0]) +
	( 16'sd 28406) * $signed(input_fmap_2[15:0]) +
	( 12'sd 2008) * $signed(input_fmap_3[15:0]) +
	( 15'sd 12649) * $signed(input_fmap_4[15:0]) +
	( 15'sd 13122) * $signed(input_fmap_5[15:0]) +
	( 15'sd 16285) * $signed(input_fmap_6[15:0]) +
	( 16'sd 21909) * $signed(input_fmap_7[15:0]) +
	( 16'sd 23324) * $signed(input_fmap_8[15:0]) +
	( 14'sd 6354) * $signed(input_fmap_9[15:0]) +
	( 16'sd 27913) * $signed(input_fmap_10[15:0]) +
	( 14'sd 5357) * $signed(input_fmap_11[15:0]) +
	( 16'sd 16821) * $signed(input_fmap_12[15:0]) +
	( 13'sd 3083) * $signed(input_fmap_13[15:0]) +
	( 16'sd 19540) * $signed(input_fmap_14[15:0]) +
	( 16'sd 18991) * $signed(input_fmap_15[15:0]) +
	( 16'sd 26509) * $signed(input_fmap_16[15:0]) +
	( 15'sd 8368) * $signed(input_fmap_17[15:0]) +
	( 16'sd 19615) * $signed(input_fmap_18[15:0]) +
	( 15'sd 10609) * $signed(input_fmap_19[15:0]) +
	( 16'sd 24303) * $signed(input_fmap_20[15:0]) +
	( 16'sd 22045) * $signed(input_fmap_21[15:0]) +
	( 16'sd 32417) * $signed(input_fmap_22[15:0]) +
	( 15'sd 9927) * $signed(input_fmap_23[15:0]) +
	( 16'sd 29338) * $signed(input_fmap_24[15:0]) +
	( 16'sd 24806) * $signed(input_fmap_25[15:0]) +
	( 15'sd 12970) * $signed(input_fmap_26[15:0]) +
	( 16'sd 30597) * $signed(input_fmap_27[15:0]) +
	( 13'sd 3869) * $signed(input_fmap_28[15:0]) +
	( 15'sd 14057) * $signed(input_fmap_29[15:0]) +
	( 16'sd 19675) * $signed(input_fmap_30[15:0]) +
	( 16'sd 21166) * $signed(input_fmap_31[15:0]) +
	( 15'sd 15821) * $signed(input_fmap_32[15:0]) +
	( 16'sd 16556) * $signed(input_fmap_33[15:0]) +
	( 16'sd 22739) * $signed(input_fmap_34[15:0]) +
	( 11'sd 868) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2078) * $signed(input_fmap_36[15:0]) +
	( 15'sd 8593) * $signed(input_fmap_37[15:0]) +
	( 11'sd 927) * $signed(input_fmap_38[15:0]) +
	( 15'sd 11634) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6961) * $signed(input_fmap_40[15:0]) +
	( 14'sd 4750) * $signed(input_fmap_41[15:0]) +
	( 15'sd 10333) * $signed(input_fmap_42[15:0]) +
	( 15'sd 8728) * $signed(input_fmap_43[15:0]) +
	( 16'sd 28803) * $signed(input_fmap_44[15:0]) +
	( 15'sd 11441) * $signed(input_fmap_45[15:0]) +
	( 16'sd 22794) * $signed(input_fmap_46[15:0]) +
	( 14'sd 4515) * $signed(input_fmap_47[15:0]) +
	( 16'sd 27112) * $signed(input_fmap_48[15:0]) +
	( 14'sd 7584) * $signed(input_fmap_49[15:0]) +
	( 15'sd 12783) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15072) * $signed(input_fmap_51[15:0]) +
	( 15'sd 8958) * $signed(input_fmap_52[15:0]) +
	( 16'sd 28619) * $signed(input_fmap_53[15:0]) +
	( 14'sd 5302) * $signed(input_fmap_54[15:0]) +
	( 14'sd 5490) * $signed(input_fmap_55[15:0]) +
	( 13'sd 3249) * $signed(input_fmap_56[15:0]) +
	( 16'sd 30544) * $signed(input_fmap_57[15:0]) +
	( 16'sd 20781) * $signed(input_fmap_58[15:0]) +
	( 16'sd 26524) * $signed(input_fmap_59[15:0]) +
	( 15'sd 14628) * $signed(input_fmap_60[15:0]) +
	( 16'sd 18608) * $signed(input_fmap_61[15:0]) +
	( 16'sd 25951) * $signed(input_fmap_62[15:0]) +
	( 16'sd 16654) * $signed(input_fmap_63[15:0]) +
	( 13'sd 2356) * $signed(input_fmap_64[15:0]) +
	( 15'sd 12706) * $signed(input_fmap_65[15:0]) +
	( 16'sd 27652) * $signed(input_fmap_66[15:0]) +
	( 11'sd 678) * $signed(input_fmap_67[15:0]) +
	( 16'sd 32429) * $signed(input_fmap_68[15:0]) +
	( 12'sd 1412) * $signed(input_fmap_69[15:0]) +
	( 14'sd 5582) * $signed(input_fmap_70[15:0]) +
	( 15'sd 8617) * $signed(input_fmap_71[15:0]) +
	( 16'sd 20072) * $signed(input_fmap_72[15:0]) +
	( 12'sd 1588) * $signed(input_fmap_73[15:0]) +
	( 16'sd 24429) * $signed(input_fmap_74[15:0]) +
	( 11'sd 928) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19520) * $signed(input_fmap_76[15:0]) +
	( 15'sd 10995) * $signed(input_fmap_77[15:0]) +
	( 15'sd 12822) * $signed(input_fmap_78[15:0]) +
	( 15'sd 14554) * $signed(input_fmap_79[15:0]) +
	( 15'sd 10725) * $signed(input_fmap_80[15:0]) +
	( 14'sd 7036) * $signed(input_fmap_81[15:0]) +
	( 14'sd 7244) * $signed(input_fmap_82[15:0]) +
	( 16'sd 17695) * $signed(input_fmap_83[15:0]) +
	( 16'sd 16623) * $signed(input_fmap_84[15:0]) +
	( 16'sd 20329) * $signed(input_fmap_85[15:0]) +
	( 16'sd 25713) * $signed(input_fmap_86[15:0]) +
	( 16'sd 25777) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6216) * $signed(input_fmap_88[15:0]) +
	( 16'sd 30432) * $signed(input_fmap_89[15:0]) +
	( 16'sd 32049) * $signed(input_fmap_90[15:0]) +
	( 14'sd 5814) * $signed(input_fmap_91[15:0]) +
	( 15'sd 14686) * $signed(input_fmap_92[15:0]) +
	( 15'sd 11679) * $signed(input_fmap_93[15:0]) +
	( 15'sd 10623) * $signed(input_fmap_94[15:0]) +
	( 15'sd 10424) * $signed(input_fmap_95[15:0]) +
	( 16'sd 23270) * $signed(input_fmap_96[15:0]) +
	( 16'sd 28250) * $signed(input_fmap_97[15:0]) +
	( 14'sd 4563) * $signed(input_fmap_98[15:0]) +
	( 16'sd 24339) * $signed(input_fmap_99[15:0]) +
	( 16'sd 21521) * $signed(input_fmap_100[15:0]) +
	( 16'sd 29834) * $signed(input_fmap_101[15:0]) +
	( 16'sd 27077) * $signed(input_fmap_102[15:0]) +
	( 15'sd 14997) * $signed(input_fmap_103[15:0]) +
	( 13'sd 2123) * $signed(input_fmap_104[15:0]) +
	( 16'sd 17304) * $signed(input_fmap_105[15:0]) +
	( 16'sd 29877) * $signed(input_fmap_106[15:0]) +
	( 16'sd 24443) * $signed(input_fmap_107[15:0]) +
	( 16'sd 28692) * $signed(input_fmap_108[15:0]) +
	( 15'sd 10636) * $signed(input_fmap_109[15:0]) +
	( 13'sd 2462) * $signed(input_fmap_110[15:0]) +
	( 16'sd 26522) * $signed(input_fmap_111[15:0]) +
	( 14'sd 7642) * $signed(input_fmap_112[15:0]) +
	( 15'sd 14863) * $signed(input_fmap_113[15:0]) +
	( 16'sd 27482) * $signed(input_fmap_114[15:0]) +
	( 16'sd 20824) * $signed(input_fmap_115[15:0]) +
	( 16'sd 17158) * $signed(input_fmap_116[15:0]) +
	( 14'sd 7076) * $signed(input_fmap_117[15:0]) +
	( 15'sd 15836) * $signed(input_fmap_118[15:0]) +
	( 16'sd 25232) * $signed(input_fmap_119[15:0]) +
	( 9'sd 253) * $signed(input_fmap_120[15:0]) +
	( 14'sd 4723) * $signed(input_fmap_121[15:0]) +
	( 16'sd 20487) * $signed(input_fmap_122[15:0]) +
	( 16'sd 27031) * $signed(input_fmap_123[15:0]) +
	( 15'sd 11063) * $signed(input_fmap_124[15:0]) +
	( 16'sd 27686) * $signed(input_fmap_125[15:0]) +
	( 13'sd 3298) * $signed(input_fmap_126[15:0]) +
	( 15'sd 12134) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 14'sd 5584) * $signed(input_fmap_0[15:0]) +
	( 16'sd 16733) * $signed(input_fmap_1[15:0]) +
	( 16'sd 20476) * $signed(input_fmap_2[15:0]) +
	( 15'sd 11019) * $signed(input_fmap_3[15:0]) +
	( 15'sd 11957) * $signed(input_fmap_4[15:0]) +
	( 14'sd 6256) * $signed(input_fmap_5[15:0]) +
	( 14'sd 6184) * $signed(input_fmap_6[15:0]) +
	( 16'sd 29202) * $signed(input_fmap_7[15:0]) +
	( 15'sd 12836) * $signed(input_fmap_8[15:0]) +
	( 16'sd 24520) * $signed(input_fmap_9[15:0]) +
	( 15'sd 14667) * $signed(input_fmap_10[15:0]) +
	( 16'sd 18744) * $signed(input_fmap_11[15:0]) +
	( 16'sd 17659) * $signed(input_fmap_12[15:0]) +
	( 16'sd 18475) * $signed(input_fmap_13[15:0]) +
	( 15'sd 10273) * $signed(input_fmap_14[15:0]) +
	( 15'sd 13335) * $signed(input_fmap_15[15:0]) +
	( 14'sd 8118) * $signed(input_fmap_16[15:0]) +
	( 15'sd 13003) * $signed(input_fmap_17[15:0]) +
	( 16'sd 16701) * $signed(input_fmap_18[15:0]) +
	( 16'sd 24829) * $signed(input_fmap_19[15:0]) +
	( 16'sd 27551) * $signed(input_fmap_20[15:0]) +
	( 15'sd 13394) * $signed(input_fmap_21[15:0]) +
	( 11'sd 885) * $signed(input_fmap_22[15:0]) +
	( 16'sd 19092) * $signed(input_fmap_23[15:0]) +
	( 16'sd 30522) * $signed(input_fmap_24[15:0]) +
	( 15'sd 14707) * $signed(input_fmap_25[15:0]) +
	( 15'sd 12454) * $signed(input_fmap_26[15:0]) +
	( 16'sd 19445) * $signed(input_fmap_27[15:0]) +
	( 16'sd 18358) * $signed(input_fmap_28[15:0]) +
	( 16'sd 26650) * $signed(input_fmap_29[15:0]) +
	( 16'sd 23521) * $signed(input_fmap_30[15:0]) +
	( 13'sd 3535) * $signed(input_fmap_31[15:0]) +
	( 16'sd 19240) * $signed(input_fmap_32[15:0]) +
	( 16'sd 29877) * $signed(input_fmap_33[15:0]) +
	( 13'sd 3832) * $signed(input_fmap_34[15:0]) +
	( 16'sd 18634) * $signed(input_fmap_35[15:0]) +
	( 14'sd 5619) * $signed(input_fmap_36[15:0]) +
	( 15'sd 13862) * $signed(input_fmap_37[15:0]) +
	( 16'sd 28264) * $signed(input_fmap_38[15:0]) +
	( 14'sd 7864) * $signed(input_fmap_39[15:0]) +
	( 16'sd 30092) * $signed(input_fmap_40[15:0]) +
	( 16'sd 22506) * $signed(input_fmap_41[15:0]) +
	( 16'sd 26552) * $signed(input_fmap_42[15:0]) +
	( 15'sd 8719) * $signed(input_fmap_43[15:0]) +
	( 16'sd 21169) * $signed(input_fmap_44[15:0]) +
	( 16'sd 29286) * $signed(input_fmap_45[15:0]) +
	( 13'sd 2805) * $signed(input_fmap_46[15:0]) +
	( 13'sd 2195) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13814) * $signed(input_fmap_48[15:0]) +
	( 16'sd 17482) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26364) * $signed(input_fmap_50[15:0]) +
	( 15'sd 13549) * $signed(input_fmap_51[15:0]) +
	( 16'sd 31837) * $signed(input_fmap_52[15:0]) +
	( 16'sd 31394) * $signed(input_fmap_53[15:0]) +
	( 16'sd 25756) * $signed(input_fmap_54[15:0]) +
	( 16'sd 28659) * $signed(input_fmap_55[15:0]) +
	( 15'sd 15661) * $signed(input_fmap_56[15:0]) +
	( 16'sd 18637) * $signed(input_fmap_57[15:0]) +
	( 14'sd 6403) * $signed(input_fmap_58[15:0]) +
	( 16'sd 19971) * $signed(input_fmap_59[15:0]) +
	( 16'sd 30720) * $signed(input_fmap_60[15:0]) +
	( 16'sd 21394) * $signed(input_fmap_61[15:0]) +
	( 12'sd 1333) * $signed(input_fmap_62[15:0]) +
	( 15'sd 10618) * $signed(input_fmap_63[15:0]) +
	( 11'sd 660) * $signed(input_fmap_64[15:0]) +
	( 16'sd 29085) * $signed(input_fmap_65[15:0]) +
	( 11'sd 583) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28232) * $signed(input_fmap_67[15:0]) +
	( 15'sd 16193) * $signed(input_fmap_68[15:0]) +
	( 15'sd 11381) * $signed(input_fmap_69[15:0]) +
	( 16'sd 19970) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31564) * $signed(input_fmap_71[15:0]) +
	( 16'sd 23482) * $signed(input_fmap_72[15:0]) +
	( 13'sd 3842) * $signed(input_fmap_73[15:0]) +
	( 16'sd 17165) * $signed(input_fmap_74[15:0]) +
	( 14'sd 7306) * $signed(input_fmap_75[15:0]) +
	( 14'sd 5049) * $signed(input_fmap_76[15:0]) +
	( 16'sd 22561) * $signed(input_fmap_77[15:0]) +
	( 16'sd 32384) * $signed(input_fmap_78[15:0]) +
	( 16'sd 16841) * $signed(input_fmap_79[15:0]) +
	( 16'sd 26651) * $signed(input_fmap_80[15:0]) +
	( 14'sd 5619) * $signed(input_fmap_81[15:0]) +
	( 16'sd 18382) * $signed(input_fmap_82[15:0]) +
	( 16'sd 18109) * $signed(input_fmap_83[15:0]) +
	( 16'sd 19824) * $signed(input_fmap_84[15:0]) +
	( 16'sd 29470) * $signed(input_fmap_85[15:0]) +
	( 15'sd 12974) * $signed(input_fmap_86[15:0]) +
	( 15'sd 11111) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6852) * $signed(input_fmap_88[15:0]) +
	( 15'sd 15872) * $signed(input_fmap_89[15:0]) +
	( 16'sd 26664) * $signed(input_fmap_90[15:0]) +
	( 16'sd 20979) * $signed(input_fmap_91[15:0]) +
	( 13'sd 2648) * $signed(input_fmap_92[15:0]) +
	( 16'sd 16870) * $signed(input_fmap_93[15:0]) +
	( 12'sd 1740) * $signed(input_fmap_94[15:0]) +
	( 14'sd 6487) * $signed(input_fmap_95[15:0]) +
	( 16'sd 26137) * $signed(input_fmap_96[15:0]) +
	( 13'sd 4019) * $signed(input_fmap_97[15:0]) +
	( 16'sd 27218) * $signed(input_fmap_98[15:0]) +
	( 14'sd 5492) * $signed(input_fmap_99[15:0]) +
	( 16'sd 28899) * $signed(input_fmap_100[15:0]) +
	( 11'sd 696) * $signed(input_fmap_101[15:0]) +
	( 16'sd 17241) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28336) * $signed(input_fmap_103[15:0]) +
	( 16'sd 32002) * $signed(input_fmap_104[15:0]) +
	( 16'sd 26810) * $signed(input_fmap_105[15:0]) +
	( 15'sd 14984) * $signed(input_fmap_106[15:0]) +
	( 16'sd 19129) * $signed(input_fmap_107[15:0]) +
	( 16'sd 27384) * $signed(input_fmap_108[15:0]) +
	( 16'sd 32748) * $signed(input_fmap_109[15:0]) +
	( 16'sd 27935) * $signed(input_fmap_110[15:0]) +
	( 16'sd 27781) * $signed(input_fmap_111[15:0]) +
	( 16'sd 30509) * $signed(input_fmap_112[15:0]) +
	( 16'sd 31427) * $signed(input_fmap_113[15:0]) +
	( 16'sd 22613) * $signed(input_fmap_114[15:0]) +
	( 16'sd 26619) * $signed(input_fmap_115[15:0]) +
	( 16'sd 30556) * $signed(input_fmap_116[15:0]) +
	( 14'sd 6394) * $signed(input_fmap_117[15:0]) +
	( 15'sd 13315) * $signed(input_fmap_118[15:0]) +
	( 15'sd 11170) * $signed(input_fmap_119[15:0]) +
	( 15'sd 14836) * $signed(input_fmap_120[15:0]) +
	( 15'sd 11028) * $signed(input_fmap_121[15:0]) +
	( 16'sd 29879) * $signed(input_fmap_122[15:0]) +
	( 16'sd 17495) * $signed(input_fmap_123[15:0]) +
	( 16'sd 21518) * $signed(input_fmap_124[15:0]) +
	( 16'sd 28193) * $signed(input_fmap_125[15:0]) +
	( 16'sd 18600) * $signed(input_fmap_126[15:0]) +
	( 16'sd 24920) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 15'sd 12361) * $signed(input_fmap_0[15:0]) +
	( 16'sd 25343) * $signed(input_fmap_1[15:0]) +
	( 16'sd 28120) * $signed(input_fmap_2[15:0]) +
	( 15'sd 11051) * $signed(input_fmap_3[15:0]) +
	( 13'sd 2513) * $signed(input_fmap_4[15:0]) +
	( 13'sd 2419) * $signed(input_fmap_5[15:0]) +
	( 15'sd 15258) * $signed(input_fmap_6[15:0]) +
	( 14'sd 6210) * $signed(input_fmap_7[15:0]) +
	( 13'sd 3424) * $signed(input_fmap_8[15:0]) +
	( 16'sd 30195) * $signed(input_fmap_9[15:0]) +
	( 14'sd 7263) * $signed(input_fmap_10[15:0]) +
	( 14'sd 6833) * $signed(input_fmap_11[15:0]) +
	( 16'sd 32436) * $signed(input_fmap_12[15:0]) +
	( 16'sd 27455) * $signed(input_fmap_13[15:0]) +
	( 14'sd 7830) * $signed(input_fmap_14[15:0]) +
	( 15'sd 10608) * $signed(input_fmap_15[15:0]) +
	( 13'sd 2566) * $signed(input_fmap_16[15:0]) +
	( 15'sd 14578) * $signed(input_fmap_17[15:0]) +
	( 15'sd 8326) * $signed(input_fmap_18[15:0]) +
	( 15'sd 13254) * $signed(input_fmap_19[15:0]) +
	( 14'sd 7120) * $signed(input_fmap_20[15:0]) +
	( 15'sd 12176) * $signed(input_fmap_21[15:0]) +
	( 15'sd 11053) * $signed(input_fmap_22[15:0]) +
	( 15'sd 14956) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17278) * $signed(input_fmap_24[15:0]) +
	( 13'sd 2368) * $signed(input_fmap_25[15:0]) +
	( 16'sd 18686) * $signed(input_fmap_26[15:0]) +
	( 16'sd 28887) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24404) * $signed(input_fmap_28[15:0]) +
	( 16'sd 27206) * $signed(input_fmap_29[15:0]) +
	( 15'sd 9325) * $signed(input_fmap_30[15:0]) +
	( 16'sd 24121) * $signed(input_fmap_31[15:0]) +
	( 16'sd 20756) * $signed(input_fmap_32[15:0]) +
	( 16'sd 25251) * $signed(input_fmap_33[15:0]) +
	( 15'sd 10323) * $signed(input_fmap_34[15:0]) +
	( 16'sd 32201) * $signed(input_fmap_35[15:0]) +
	( 16'sd 30664) * $signed(input_fmap_36[15:0]) +
	( 16'sd 29695) * $signed(input_fmap_37[15:0]) +
	( 15'sd 15344) * $signed(input_fmap_38[15:0]) +
	( 15'sd 10645) * $signed(input_fmap_39[15:0]) +
	( 16'sd 20093) * $signed(input_fmap_40[15:0]) +
	( 13'sd 3198) * $signed(input_fmap_41[15:0]) +
	( 13'sd 3594) * $signed(input_fmap_42[15:0]) +
	( 16'sd 24063) * $signed(input_fmap_43[15:0]) +
	( 16'sd 30722) * $signed(input_fmap_44[15:0]) +
	( 13'sd 3616) * $signed(input_fmap_45[15:0]) +
	( 9'sd 217) * $signed(input_fmap_46[15:0]) +
	( 13'sd 3341) * $signed(input_fmap_47[15:0]) +
	( 13'sd 3356) * $signed(input_fmap_48[15:0]) +
	( 16'sd 27213) * $signed(input_fmap_49[15:0]) +
	( 16'sd 32408) * $signed(input_fmap_50[15:0]) +
	( 16'sd 23383) * $signed(input_fmap_51[15:0]) +
	( 16'sd 25021) * $signed(input_fmap_52[15:0]) +
	( 13'sd 3530) * $signed(input_fmap_53[15:0]) +
	( 16'sd 20186) * $signed(input_fmap_54[15:0]) +
	( 16'sd 23235) * $signed(input_fmap_55[15:0]) +
	( 14'sd 6181) * $signed(input_fmap_56[15:0]) +
	( 15'sd 15113) * $signed(input_fmap_57[15:0]) +
	( 13'sd 2114) * $signed(input_fmap_58[15:0]) +
	( 16'sd 21097) * $signed(input_fmap_59[15:0]) +
	( 16'sd 18881) * $signed(input_fmap_60[15:0]) +
	( 16'sd 20180) * $signed(input_fmap_61[15:0]) +
	( 16'sd 28331) * $signed(input_fmap_62[15:0]) +
	( 16'sd 19480) * $signed(input_fmap_63[15:0]) +
	( 16'sd 28206) * $signed(input_fmap_64[15:0]) +
	( 16'sd 21063) * $signed(input_fmap_65[15:0]) +
	( 15'sd 14521) * $signed(input_fmap_66[15:0]) +
	( 13'sd 3619) * $signed(input_fmap_67[15:0]) +
	( 16'sd 28873) * $signed(input_fmap_68[15:0]) +
	( 15'sd 11502) * $signed(input_fmap_69[15:0]) +
	( 16'sd 17750) * $signed(input_fmap_70[15:0]) +
	( 16'sd 29518) * $signed(input_fmap_71[15:0]) +
	( 16'sd 16862) * $signed(input_fmap_72[15:0]) +
	( 13'sd 2825) * $signed(input_fmap_73[15:0]) +
	( 15'sd 11775) * $signed(input_fmap_74[15:0]) +
	( 14'sd 6045) * $signed(input_fmap_75[15:0]) +
	( 15'sd 13225) * $signed(input_fmap_76[15:0]) +
	( 15'sd 10141) * $signed(input_fmap_77[15:0]) +
	( 16'sd 30363) * $signed(input_fmap_78[15:0]) +
	( 13'sd 2755) * $signed(input_fmap_79[15:0]) +
	( 8'sd 108) * $signed(input_fmap_80[15:0]) +
	( 15'sd 11051) * $signed(input_fmap_81[15:0]) +
	( 14'sd 7274) * $signed(input_fmap_82[15:0]) +
	( 15'sd 14113) * $signed(input_fmap_83[15:0]) +
	( 16'sd 26850) * $signed(input_fmap_84[15:0]) +
	( 15'sd 15428) * $signed(input_fmap_85[15:0]) +
	( 14'sd 5439) * $signed(input_fmap_86[15:0]) +
	( 16'sd 18296) * $signed(input_fmap_87[15:0]) +
	( 16'sd 30710) * $signed(input_fmap_88[15:0]) +
	( 15'sd 12780) * $signed(input_fmap_89[15:0]) +
	( 14'sd 5265) * $signed(input_fmap_90[15:0]) +
	( 15'sd 12277) * $signed(input_fmap_91[15:0]) +
	( 16'sd 16605) * $signed(input_fmap_92[15:0]) +
	( 14'sd 5029) * $signed(input_fmap_93[15:0]) +
	( 15'sd 15169) * $signed(input_fmap_94[15:0]) +
	( 15'sd 10442) * $signed(input_fmap_95[15:0]) +
	( 16'sd 30384) * $signed(input_fmap_96[15:0]) +
	( 16'sd 18201) * $signed(input_fmap_97[15:0]) +
	( 13'sd 2901) * $signed(input_fmap_98[15:0]) +
	( 16'sd 31644) * $signed(input_fmap_99[15:0]) +
	( 15'sd 8987) * $signed(input_fmap_100[15:0]) +
	( 16'sd 19467) * $signed(input_fmap_101[15:0]) +
	( 13'sd 4089) * $signed(input_fmap_102[15:0]) +
	( 12'sd 1788) * $signed(input_fmap_103[15:0]) +
	( 16'sd 21611) * $signed(input_fmap_104[15:0]) +
	( 15'sd 13825) * $signed(input_fmap_105[15:0]) +
	( 14'sd 7774) * $signed(input_fmap_106[15:0]) +
	( 13'sd 2417) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15626) * $signed(input_fmap_108[15:0]) +
	( 16'sd 17893) * $signed(input_fmap_109[15:0]) +
	( 15'sd 14747) * $signed(input_fmap_110[15:0]) +
	( 15'sd 16278) * $signed(input_fmap_111[15:0]) +
	( 12'sd 1205) * $signed(input_fmap_112[15:0]) +
	( 16'sd 20239) * $signed(input_fmap_113[15:0]) +
	( 16'sd 24982) * $signed(input_fmap_114[15:0]) +
	( 16'sd 30201) * $signed(input_fmap_115[15:0]) +
	( 16'sd 17913) * $signed(input_fmap_116[15:0]) +
	( 15'sd 11813) * $signed(input_fmap_117[15:0]) +
	( 16'sd 27875) * $signed(input_fmap_118[15:0]) +
	( 16'sd 17265) * $signed(input_fmap_119[15:0]) +
	( 15'sd 16056) * $signed(input_fmap_120[15:0]) +
	( 16'sd 30488) * $signed(input_fmap_121[15:0]) +
	( 14'sd 6563) * $signed(input_fmap_122[15:0]) +
	( 16'sd 22309) * $signed(input_fmap_123[15:0]) +
	( 16'sd 26271) * $signed(input_fmap_124[15:0]) +
	( 13'sd 2084) * $signed(input_fmap_125[15:0]) +
	( 14'sd 7487) * $signed(input_fmap_126[15:0]) +
	( 16'sd 26909) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 15'sd 12603) * $signed(input_fmap_0[15:0]) +
	( 16'sd 30349) * $signed(input_fmap_1[15:0]) +
	( 16'sd 31555) * $signed(input_fmap_2[15:0]) +
	( 12'sd 1654) * $signed(input_fmap_3[15:0]) +
	( 16'sd 27130) * $signed(input_fmap_4[15:0]) +
	( 16'sd 32487) * $signed(input_fmap_5[15:0]) +
	( 14'sd 5102) * $signed(input_fmap_6[15:0]) +
	( 16'sd 22013) * $signed(input_fmap_7[15:0]) +
	( 16'sd 30928) * $signed(input_fmap_8[15:0]) +
	( 14'sd 4739) * $signed(input_fmap_9[15:0]) +
	( 11'sd 639) * $signed(input_fmap_10[15:0]) +
	( 14'sd 7519) * $signed(input_fmap_11[15:0]) +
	( 14'sd 4748) * $signed(input_fmap_12[15:0]) +
	( 16'sd 25598) * $signed(input_fmap_13[15:0]) +
	( 16'sd 24796) * $signed(input_fmap_14[15:0]) +
	( 15'sd 9839) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10977) * $signed(input_fmap_16[15:0]) +
	( 15'sd 15581) * $signed(input_fmap_17[15:0]) +
	( 16'sd 29974) * $signed(input_fmap_18[15:0]) +
	( 15'sd 16251) * $signed(input_fmap_19[15:0]) +
	( 14'sd 8152) * $signed(input_fmap_20[15:0]) +
	( 15'sd 14420) * $signed(input_fmap_21[15:0]) +
	( 14'sd 4146) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24631) * $signed(input_fmap_23[15:0]) +
	( 16'sd 27574) * $signed(input_fmap_24[15:0]) +
	( 15'sd 12437) * $signed(input_fmap_25[15:0]) +
	( 14'sd 7133) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1246) * $signed(input_fmap_27[15:0]) +
	( 15'sd 13197) * $signed(input_fmap_28[15:0]) +
	( 9'sd 235) * $signed(input_fmap_29[15:0]) +
	( 15'sd 10941) * $signed(input_fmap_30[15:0]) +
	( 16'sd 30063) * $signed(input_fmap_31[15:0]) +
	( 16'sd 32340) * $signed(input_fmap_32[15:0]) +
	( 14'sd 5133) * $signed(input_fmap_33[15:0]) +
	( 16'sd 24993) * $signed(input_fmap_34[15:0]) +
	( 16'sd 29770) * $signed(input_fmap_35[15:0]) +
	( 16'sd 28665) * $signed(input_fmap_36[15:0]) +
	( 10'sd 478) * $signed(input_fmap_37[15:0]) +
	( 15'sd 13914) * $signed(input_fmap_38[15:0]) +
	( 16'sd 22163) * $signed(input_fmap_39[15:0]) +
	( 10'sd 326) * $signed(input_fmap_40[15:0]) +
	( 13'sd 3768) * $signed(input_fmap_41[15:0]) +
	( 16'sd 17169) * $signed(input_fmap_42[15:0]) +
	( 16'sd 31280) * $signed(input_fmap_43[15:0]) +
	( 14'sd 7271) * $signed(input_fmap_44[15:0]) +
	( 15'sd 9816) * $signed(input_fmap_45[15:0]) +
	( 14'sd 7004) * $signed(input_fmap_46[15:0]) +
	( 16'sd 24353) * $signed(input_fmap_47[15:0]) +
	( 16'sd 21304) * $signed(input_fmap_48[15:0]) +
	( 16'sd 23203) * $signed(input_fmap_49[15:0]) +
	( 16'sd 30698) * $signed(input_fmap_50[15:0]) +
	( 10'sd 322) * $signed(input_fmap_51[15:0]) +
	( 15'sd 8784) * $signed(input_fmap_52[15:0]) +
	( 15'sd 15601) * $signed(input_fmap_53[15:0]) +
	( 16'sd 29114) * $signed(input_fmap_54[15:0]) +
	( 15'sd 12094) * $signed(input_fmap_55[15:0]) +
	( 16'sd 22396) * $signed(input_fmap_56[15:0]) +
	( 14'sd 5782) * $signed(input_fmap_57[15:0]) +
	( 15'sd 9452) * $signed(input_fmap_58[15:0]) +
	( 16'sd 22123) * $signed(input_fmap_59[15:0]) +
	( 15'sd 16124) * $signed(input_fmap_60[15:0]) +
	( 15'sd 13947) * $signed(input_fmap_61[15:0]) +
	( 16'sd 17918) * $signed(input_fmap_62[15:0]) +
	( 16'sd 17863) * $signed(input_fmap_63[15:0]) +
	( 16'sd 18137) * $signed(input_fmap_64[15:0]) +
	( 16'sd 21195) * $signed(input_fmap_65[15:0]) +
	( 15'sd 12105) * $signed(input_fmap_66[15:0]) +
	( 13'sd 3331) * $signed(input_fmap_67[15:0]) +
	( 15'sd 12123) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31774) * $signed(input_fmap_69[15:0]) +
	( 14'sd 4562) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11781) * $signed(input_fmap_71[15:0]) +
	( 16'sd 24372) * $signed(input_fmap_72[15:0]) +
	( 15'sd 8523) * $signed(input_fmap_73[15:0]) +
	( 14'sd 6352) * $signed(input_fmap_74[15:0]) +
	( 16'sd 29522) * $signed(input_fmap_75[15:0]) +
	( 16'sd 18816) * $signed(input_fmap_76[15:0]) +
	( 14'sd 7935) * $signed(input_fmap_77[15:0]) +
	( 16'sd 22228) * $signed(input_fmap_78[15:0]) +
	( 12'sd 2029) * $signed(input_fmap_79[15:0]) +
	( 16'sd 23189) * $signed(input_fmap_80[15:0]) +
	( 16'sd 29404) * $signed(input_fmap_81[15:0]) +
	( 15'sd 8312) * $signed(input_fmap_82[15:0]) +
	( 16'sd 19229) * $signed(input_fmap_83[15:0]) +
	( 15'sd 12676) * $signed(input_fmap_84[15:0]) +
	( 12'sd 1474) * $signed(input_fmap_85[15:0]) +
	( 16'sd 29330) * $signed(input_fmap_86[15:0]) +
	( 16'sd 20509) * $signed(input_fmap_87[15:0]) +
	( 16'sd 27718) * $signed(input_fmap_88[15:0]) +
	( 14'sd 4818) * $signed(input_fmap_89[15:0]) +
	( 16'sd 21111) * $signed(input_fmap_90[15:0]) +
	( 14'sd 4343) * $signed(input_fmap_91[15:0]) +
	( 13'sd 3267) * $signed(input_fmap_92[15:0]) +
	( 16'sd 32340) * $signed(input_fmap_93[15:0]) +
	( 16'sd 22952) * $signed(input_fmap_94[15:0]) +
	( 15'sd 9748) * $signed(input_fmap_95[15:0]) +
	( 13'sd 3529) * $signed(input_fmap_96[15:0]) +
	( 16'sd 20085) * $signed(input_fmap_97[15:0]) +
	( 15'sd 14894) * $signed(input_fmap_98[15:0]) +
	( 13'sd 2546) * $signed(input_fmap_99[15:0]) +
	( 16'sd 21052) * $signed(input_fmap_100[15:0]) +
	( 16'sd 17403) * $signed(input_fmap_101[15:0]) +
	( 16'sd 18970) * $signed(input_fmap_102[15:0]) +
	( 16'sd 27904) * $signed(input_fmap_103[15:0]) +
	( 15'sd 14039) * $signed(input_fmap_104[15:0]) +
	( 16'sd 32737) * $signed(input_fmap_105[15:0]) +
	( 15'sd 11656) * $signed(input_fmap_106[15:0]) +
	( 16'sd 17648) * $signed(input_fmap_107[15:0]) +
	( 16'sd 22486) * $signed(input_fmap_108[15:0]) +
	( 16'sd 20537) * $signed(input_fmap_109[15:0]) +
	( 16'sd 21363) * $signed(input_fmap_110[15:0]) +
	( 16'sd 19491) * $signed(input_fmap_111[15:0]) +
	( 14'sd 4829) * $signed(input_fmap_112[15:0]) +
	( 16'sd 30248) * $signed(input_fmap_113[15:0]) +
	( 16'sd 16476) * $signed(input_fmap_114[15:0]) +
	( 15'sd 11748) * $signed(input_fmap_115[15:0]) +
	( 12'sd 1032) * $signed(input_fmap_116[15:0]) +
	( 14'sd 7143) * $signed(input_fmap_117[15:0]) +
	( 16'sd 21728) * $signed(input_fmap_118[15:0]) +
	( 13'sd 3647) * $signed(input_fmap_119[15:0]) +
	( 14'sd 5422) * $signed(input_fmap_120[15:0]) +
	( 16'sd 20152) * $signed(input_fmap_121[15:0]) +
	( 16'sd 31474) * $signed(input_fmap_122[15:0]) +
	( 14'sd 6783) * $signed(input_fmap_123[15:0]) +
	( 12'sd 1271) * $signed(input_fmap_124[15:0]) +
	( 16'sd 23975) * $signed(input_fmap_125[15:0]) +
	( 8'sd 112) * $signed(input_fmap_126[15:0]) +
	( 16'sd 32228) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 14'sd 7726) * $signed(input_fmap_0[15:0]) +
	( 16'sd 18272) * $signed(input_fmap_1[15:0]) +
	( 16'sd 26149) * $signed(input_fmap_2[15:0]) +
	( 11'sd 916) * $signed(input_fmap_3[15:0]) +
	( 15'sd 15463) * $signed(input_fmap_4[15:0]) +
	( 16'sd 19101) * $signed(input_fmap_5[15:0]) +
	( 16'sd 29093) * $signed(input_fmap_6[15:0]) +
	( 14'sd 7598) * $signed(input_fmap_7[15:0]) +
	( 15'sd 9254) * $signed(input_fmap_8[15:0]) +
	( 16'sd 20024) * $signed(input_fmap_9[15:0]) +
	( 16'sd 30923) * $signed(input_fmap_10[15:0]) +
	( 16'sd 26356) * $signed(input_fmap_11[15:0]) +
	( 14'sd 6104) * $signed(input_fmap_12[15:0]) +
	( 16'sd 23054) * $signed(input_fmap_13[15:0]) +
	( 13'sd 2181) * $signed(input_fmap_14[15:0]) +
	( 12'sd 1336) * $signed(input_fmap_15[15:0]) +
	( 12'sd 1714) * $signed(input_fmap_16[15:0]) +
	( 13'sd 3468) * $signed(input_fmap_17[15:0]) +
	( 16'sd 28001) * $signed(input_fmap_18[15:0]) +
	( 16'sd 16555) * $signed(input_fmap_19[15:0]) +
	( 13'sd 2664) * $signed(input_fmap_20[15:0]) +
	( 16'sd 29347) * $signed(input_fmap_21[15:0]) +
	( 16'sd 24995) * $signed(input_fmap_22[15:0]) +
	( 16'sd 19225) * $signed(input_fmap_23[15:0]) +
	( 16'sd 26760) * $signed(input_fmap_24[15:0]) +
	( 16'sd 20446) * $signed(input_fmap_25[15:0]) +
	( 16'sd 31623) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9944) * $signed(input_fmap_27[15:0]) +
	( 11'sd 973) * $signed(input_fmap_28[15:0]) +
	( 16'sd 30765) * $signed(input_fmap_29[15:0]) +
	( 16'sd 19619) * $signed(input_fmap_30[15:0]) +
	( 14'sd 6840) * $signed(input_fmap_31[15:0]) +
	( 15'sd 9763) * $signed(input_fmap_32[15:0]) +
	( 16'sd 28275) * $signed(input_fmap_33[15:0]) +
	( 16'sd 23302) * $signed(input_fmap_34[15:0]) +
	( 16'sd 17221) * $signed(input_fmap_35[15:0]) +
	( 15'sd 12774) * $signed(input_fmap_36[15:0]) +
	( 16'sd 22729) * $signed(input_fmap_37[15:0]) +
	( 15'sd 12676) * $signed(input_fmap_38[15:0]) +
	( 16'sd 19820) * $signed(input_fmap_39[15:0]) +
	( 16'sd 31098) * $signed(input_fmap_40[15:0]) +
	( 15'sd 12974) * $signed(input_fmap_41[15:0]) +
	( 16'sd 16947) * $signed(input_fmap_42[15:0]) +
	( 11'sd 675) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31905) * $signed(input_fmap_44[15:0]) +
	( 10'sd 346) * $signed(input_fmap_45[15:0]) +
	( 14'sd 4239) * $signed(input_fmap_46[15:0]) +
	( 12'sd 1587) * $signed(input_fmap_47[15:0]) +
	( 8'sd 93) * $signed(input_fmap_48[15:0]) +
	( 14'sd 5936) * $signed(input_fmap_49[15:0]) +
	( 14'sd 7913) * $signed(input_fmap_50[15:0]) +
	( 16'sd 31564) * $signed(input_fmap_51[15:0]) +
	( 16'sd 17435) * $signed(input_fmap_52[15:0]) +
	( 11'sd 912) * $signed(input_fmap_53[15:0]) +
	( 15'sd 14967) * $signed(input_fmap_54[15:0]) +
	( 16'sd 22353) * $signed(input_fmap_55[15:0]) +
	( 15'sd 14555) * $signed(input_fmap_56[15:0]) +
	( 16'sd 32271) * $signed(input_fmap_57[15:0]) +
	( 14'sd 4279) * $signed(input_fmap_58[15:0]) +
	( 15'sd 10017) * $signed(input_fmap_59[15:0]) +
	( 15'sd 11600) * $signed(input_fmap_60[15:0]) +
	( 16'sd 32080) * $signed(input_fmap_61[15:0]) +
	( 16'sd 22288) * $signed(input_fmap_62[15:0]) +
	( 16'sd 16421) * $signed(input_fmap_63[15:0]) +
	( 13'sd 3865) * $signed(input_fmap_64[15:0]) +
	( 15'sd 10975) * $signed(input_fmap_65[15:0]) +
	( 16'sd 19772) * $signed(input_fmap_66[15:0]) +
	( 15'sd 10230) * $signed(input_fmap_67[15:0]) +
	( 16'sd 17247) * $signed(input_fmap_68[15:0]) +
	( 8'sd 113) * $signed(input_fmap_69[15:0]) +
	( 15'sd 15460) * $signed(input_fmap_70[15:0]) +
	( 16'sd 24614) * $signed(input_fmap_71[15:0]) +
	( 16'sd 22177) * $signed(input_fmap_72[15:0]) +
	( 16'sd 19856) * $signed(input_fmap_73[15:0]) +
	( 16'sd 20078) * $signed(input_fmap_74[15:0]) +
	( 16'sd 23863) * $signed(input_fmap_75[15:0]) +
	( 16'sd 30279) * $signed(input_fmap_76[15:0]) +
	( 16'sd 25837) * $signed(input_fmap_77[15:0]) +
	( 16'sd 16452) * $signed(input_fmap_78[15:0]) +
	( 15'sd 16352) * $signed(input_fmap_79[15:0]) +
	( 16'sd 27219) * $signed(input_fmap_80[15:0]) +
	( 15'sd 10518) * $signed(input_fmap_81[15:0]) +
	( 15'sd 10364) * $signed(input_fmap_82[15:0]) +
	( 14'sd 7993) * $signed(input_fmap_83[15:0]) +
	( 15'sd 8215) * $signed(input_fmap_84[15:0]) +
	( 16'sd 21201) * $signed(input_fmap_85[15:0]) +
	( 15'sd 9445) * $signed(input_fmap_86[15:0]) +
	( 12'sd 1071) * $signed(input_fmap_87[15:0]) +
	( 14'sd 4419) * $signed(input_fmap_88[15:0]) +
	( 15'sd 8509) * $signed(input_fmap_89[15:0]) +
	( 15'sd 14086) * $signed(input_fmap_90[15:0]) +
	( 14'sd 7977) * $signed(input_fmap_91[15:0]) +
	( 15'sd 10737) * $signed(input_fmap_92[15:0]) +
	( 16'sd 23898) * $signed(input_fmap_93[15:0]) +
	( 16'sd 25783) * $signed(input_fmap_94[15:0]) +
	( 14'sd 4746) * $signed(input_fmap_95[15:0]) +
	( 16'sd 30379) * $signed(input_fmap_96[15:0]) +
	( 16'sd 29262) * $signed(input_fmap_97[15:0]) +
	( 15'sd 9892) * $signed(input_fmap_98[15:0]) +
	( 15'sd 12809) * $signed(input_fmap_99[15:0]) +
	( 15'sd 9062) * $signed(input_fmap_100[15:0]) +
	( 16'sd 25947) * $signed(input_fmap_101[15:0]) +
	( 15'sd 8455) * $signed(input_fmap_102[15:0]) +
	( 16'sd 19100) * $signed(input_fmap_103[15:0]) +
	( 10'sd 415) * $signed(input_fmap_104[15:0]) +
	( 14'sd 4781) * $signed(input_fmap_105[15:0]) +
	( 15'sd 15337) * $signed(input_fmap_106[15:0]) +
	( 14'sd 6136) * $signed(input_fmap_107[15:0]) +
	( 10'sd 421) * $signed(input_fmap_108[15:0]) +
	( 14'sd 5180) * $signed(input_fmap_109[15:0]) +
	( 15'sd 14584) * $signed(input_fmap_110[15:0]) +
	( 14'sd 7755) * $signed(input_fmap_111[15:0]) +
	( 16'sd 19689) * $signed(input_fmap_112[15:0]) +
	( 16'sd 20179) * $signed(input_fmap_113[15:0]) +
	( 16'sd 16843) * $signed(input_fmap_114[15:0]) +
	( 16'sd 26185) * $signed(input_fmap_115[15:0]) +
	( 16'sd 21230) * $signed(input_fmap_116[15:0]) +
	( 16'sd 30702) * $signed(input_fmap_117[15:0]) +
	( 15'sd 13040) * $signed(input_fmap_118[15:0]) +
	( 13'sd 3141) * $signed(input_fmap_119[15:0]) +
	( 16'sd 26066) * $signed(input_fmap_120[15:0]) +
	( 16'sd 17324) * $signed(input_fmap_121[15:0]) +
	( 16'sd 23709) * $signed(input_fmap_122[15:0]) +
	( 16'sd 30231) * $signed(input_fmap_123[15:0]) +
	( 13'sd 3910) * $signed(input_fmap_124[15:0]) +
	( 14'sd 4337) * $signed(input_fmap_125[15:0]) +
	( 15'sd 11160) * $signed(input_fmap_126[15:0]) +
	( 16'sd 16568) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 16'sd 23282) * $signed(input_fmap_0[15:0]) +
	( 15'sd 12635) * $signed(input_fmap_1[15:0]) +
	( 15'sd 15531) * $signed(input_fmap_2[15:0]) +
	( 16'sd 31698) * $signed(input_fmap_3[15:0]) +
	( 15'sd 15481) * $signed(input_fmap_4[15:0]) +
	( 12'sd 1238) * $signed(input_fmap_5[15:0]) +
	( 16'sd 31211) * $signed(input_fmap_6[15:0]) +
	( 13'sd 2434) * $signed(input_fmap_7[15:0]) +
	( 14'sd 7286) * $signed(input_fmap_8[15:0]) +
	( 14'sd 8144) * $signed(input_fmap_9[15:0]) +
	( 15'sd 8572) * $signed(input_fmap_10[15:0]) +
	( 15'sd 15366) * $signed(input_fmap_11[15:0]) +
	( 15'sd 15737) * $signed(input_fmap_12[15:0]) +
	( 14'sd 8134) * $signed(input_fmap_13[15:0]) +
	( 16'sd 31584) * $signed(input_fmap_14[15:0]) +
	( 16'sd 25440) * $signed(input_fmap_15[15:0]) +
	( 16'sd 29778) * $signed(input_fmap_16[15:0]) +
	( 16'sd 23862) * $signed(input_fmap_17[15:0]) +
	( 16'sd 24922) * $signed(input_fmap_18[15:0]) +
	( 16'sd 18782) * $signed(input_fmap_19[15:0]) +
	( 16'sd 30255) * $signed(input_fmap_20[15:0]) +
	( 12'sd 1411) * $signed(input_fmap_21[15:0]) +
	( 16'sd 23305) * $signed(input_fmap_22[15:0]) +
	( 16'sd 23736) * $signed(input_fmap_23[15:0]) +
	( 16'sd 16506) * $signed(input_fmap_24[15:0]) +
	( 12'sd 1071) * $signed(input_fmap_25[15:0]) +
	( 16'sd 26186) * $signed(input_fmap_26[15:0]) +
	( 16'sd 26445) * $signed(input_fmap_27[15:0]) +
	( 13'sd 2076) * $signed(input_fmap_28[15:0]) +
	( 15'sd 13285) * $signed(input_fmap_29[15:0]) +
	( 16'sd 24512) * $signed(input_fmap_30[15:0]) +
	( 13'sd 2150) * $signed(input_fmap_31[15:0]) +
	( 16'sd 29840) * $signed(input_fmap_32[15:0]) +
	( 12'sd 1505) * $signed(input_fmap_33[15:0]) +
	( 14'sd 7193) * $signed(input_fmap_34[15:0]) +
	( 15'sd 16370) * $signed(input_fmap_35[15:0]) +
	( 13'sd 3441) * $signed(input_fmap_36[15:0]) +
	( 13'sd 3767) * $signed(input_fmap_37[15:0]) +
	( 13'sd 3112) * $signed(input_fmap_38[15:0]) +
	( 14'sd 7743) * $signed(input_fmap_39[15:0]) +
	( 16'sd 23429) * $signed(input_fmap_40[15:0]) +
	( 16'sd 19756) * $signed(input_fmap_41[15:0]) +
	( 16'sd 22136) * $signed(input_fmap_42[15:0]) +
	( 15'sd 12745) * $signed(input_fmap_43[15:0]) +
	( 16'sd 23816) * $signed(input_fmap_44[15:0]) +
	( 14'sd 6037) * $signed(input_fmap_45[15:0]) +
	( 15'sd 13862) * $signed(input_fmap_46[15:0]) +
	( 14'sd 4893) * $signed(input_fmap_47[15:0]) +
	( 16'sd 22653) * $signed(input_fmap_48[15:0]) +
	( 16'sd 24169) * $signed(input_fmap_49[15:0]) +
	( 16'sd 23795) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15690) * $signed(input_fmap_51[15:0]) +
	( 15'sd 11142) * $signed(input_fmap_52[15:0]) +
	( 15'sd 13955) * $signed(input_fmap_53[15:0]) +
	( 14'sd 4345) * $signed(input_fmap_54[15:0]) +
	( 15'sd 11567) * $signed(input_fmap_55[15:0]) +
	( 16'sd 25555) * $signed(input_fmap_56[15:0]) +
	( 15'sd 15941) * $signed(input_fmap_57[15:0]) +
	( 16'sd 24952) * $signed(input_fmap_58[15:0]) +
	( 14'sd 5867) * $signed(input_fmap_59[15:0]) +
	( 16'sd 30155) * $signed(input_fmap_60[15:0]) +
	( 16'sd 23518) * $signed(input_fmap_61[15:0]) +
	( 15'sd 10202) * $signed(input_fmap_62[15:0]) +
	( 16'sd 32475) * $signed(input_fmap_63[15:0]) +
	( 12'sd 1673) * $signed(input_fmap_64[15:0]) +
	( 14'sd 7032) * $signed(input_fmap_65[15:0]) +
	( 16'sd 16784) * $signed(input_fmap_66[15:0]) +
	( 16'sd 32761) * $signed(input_fmap_67[15:0]) +
	( 16'sd 29594) * $signed(input_fmap_68[15:0]) +
	( 16'sd 30512) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31618) * $signed(input_fmap_70[15:0]) +
	( 16'sd 21842) * $signed(input_fmap_71[15:0]) +
	( 13'sd 2463) * $signed(input_fmap_72[15:0]) +
	( 16'sd 24455) * $signed(input_fmap_73[15:0]) +
	( 16'sd 28937) * $signed(input_fmap_74[15:0]) +
	( 14'sd 4278) * $signed(input_fmap_75[15:0]) +
	( 16'sd 26644) * $signed(input_fmap_76[15:0]) +
	( 16'sd 25240) * $signed(input_fmap_77[15:0]) +
	( 15'sd 11049) * $signed(input_fmap_78[15:0]) +
	( 15'sd 12549) * $signed(input_fmap_79[15:0]) +
	( 15'sd 8984) * $signed(input_fmap_80[15:0]) +
	( 16'sd 19208) * $signed(input_fmap_81[15:0]) +
	( 16'sd 28621) * $signed(input_fmap_82[15:0]) +
	( 13'sd 3566) * $signed(input_fmap_83[15:0]) +
	( 13'sd 2444) * $signed(input_fmap_84[15:0]) +
	( 16'sd 18637) * $signed(input_fmap_85[15:0]) +
	( 16'sd 31800) * $signed(input_fmap_86[15:0]) +
	( 16'sd 22271) * $signed(input_fmap_87[15:0]) +
	( 14'sd 4226) * $signed(input_fmap_88[15:0]) +
	( 13'sd 4076) * $signed(input_fmap_89[15:0]) +
	( 13'sd 3283) * $signed(input_fmap_90[15:0]) +
	( 16'sd 30111) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25291) * $signed(input_fmap_92[15:0]) +
	( 14'sd 4524) * $signed(input_fmap_93[15:0]) +
	( 16'sd 30430) * $signed(input_fmap_94[15:0]) +
	( 12'sd 1970) * $signed(input_fmap_95[15:0]) +
	( 15'sd 8293) * $signed(input_fmap_96[15:0]) +
	( 15'sd 14868) * $signed(input_fmap_97[15:0]) +
	( 16'sd 24562) * $signed(input_fmap_98[15:0]) +
	( 15'sd 11960) * $signed(input_fmap_99[15:0]) +
	( 16'sd 19716) * $signed(input_fmap_100[15:0]) +
	( 14'sd 6486) * $signed(input_fmap_101[15:0]) +
	( 15'sd 10629) * $signed(input_fmap_102[15:0]) +
	( 12'sd 1459) * $signed(input_fmap_103[15:0]) +
	( 15'sd 11618) * $signed(input_fmap_104[15:0]) +
	( 15'sd 15900) * $signed(input_fmap_105[15:0]) +
	( 15'sd 8444) * $signed(input_fmap_106[15:0]) +
	( 16'sd 16860) * $signed(input_fmap_107[15:0]) +
	( 16'sd 24999) * $signed(input_fmap_108[15:0]) +
	( 15'sd 13361) * $signed(input_fmap_109[15:0]) +
	( 16'sd 26929) * $signed(input_fmap_110[15:0]) +
	( 16'sd 16834) * $signed(input_fmap_111[15:0]) +
	( 16'sd 21356) * $signed(input_fmap_112[15:0]) +
	( 16'sd 29687) * $signed(input_fmap_113[15:0]) +
	( 12'sd 1482) * $signed(input_fmap_114[15:0]) +
	( 15'sd 13751) * $signed(input_fmap_115[15:0]) +
	( 15'sd 11209) * $signed(input_fmap_116[15:0]) +
	( 14'sd 7017) * $signed(input_fmap_117[15:0]) +
	( 16'sd 22085) * $signed(input_fmap_118[15:0]) +
	( 14'sd 6603) * $signed(input_fmap_119[15:0]) +
	( 13'sd 2307) * $signed(input_fmap_120[15:0]) +
	( 15'sd 15074) * $signed(input_fmap_121[15:0]) +
	( 16'sd 32414) * $signed(input_fmap_122[15:0]) +
	( 15'sd 9085) * $signed(input_fmap_123[15:0]) +
	( 16'sd 18295) * $signed(input_fmap_124[15:0]) +
	( 16'sd 32325) * $signed(input_fmap_125[15:0]) +
	( 16'sd 28620) * $signed(input_fmap_126[15:0]) +
	( 16'sd 23407) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 15'sd 13732) * $signed(input_fmap_0[15:0]) +
	( 16'sd 19413) * $signed(input_fmap_1[15:0]) +
	( 13'sd 2451) * $signed(input_fmap_2[15:0]) +
	( 14'sd 7746) * $signed(input_fmap_3[15:0]) +
	( 15'sd 11734) * $signed(input_fmap_4[15:0]) +
	( 15'sd 14243) * $signed(input_fmap_5[15:0]) +
	( 16'sd 26451) * $signed(input_fmap_6[15:0]) +
	( 12'sd 2042) * $signed(input_fmap_7[15:0]) +
	( 16'sd 25144) * $signed(input_fmap_8[15:0]) +
	( 16'sd 18283) * $signed(input_fmap_9[15:0]) +
	( 16'sd 25615) * $signed(input_fmap_10[15:0]) +
	( 15'sd 11983) * $signed(input_fmap_11[15:0]) +
	( 16'sd 25927) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24334) * $signed(input_fmap_13[15:0]) +
	( 15'sd 10269) * $signed(input_fmap_14[15:0]) +
	( 16'sd 19228) * $signed(input_fmap_15[15:0]) +
	( 16'sd 21993) * $signed(input_fmap_16[15:0]) +
	( 15'sd 14350) * $signed(input_fmap_17[15:0]) +
	( 15'sd 16375) * $signed(input_fmap_18[15:0]) +
	( 14'sd 5955) * $signed(input_fmap_19[15:0]) +
	( 13'sd 4090) * $signed(input_fmap_20[15:0]) +
	( 14'sd 4646) * $signed(input_fmap_21[15:0]) +
	( 15'sd 13793) * $signed(input_fmap_22[15:0]) +
	( 15'sd 11686) * $signed(input_fmap_23[15:0]) +
	( 16'sd 22370) * $signed(input_fmap_24[15:0]) +
	( 15'sd 10336) * $signed(input_fmap_25[15:0]) +
	( 15'sd 9400) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9051) * $signed(input_fmap_27[15:0]) +
	( 16'sd 30502) * $signed(input_fmap_28[15:0]) +
	( 15'sd 8750) * $signed(input_fmap_29[15:0]) +
	( 14'sd 4372) * $signed(input_fmap_30[15:0]) +
	( 13'sd 4027) * $signed(input_fmap_31[15:0]) +
	( 15'sd 13170) * $signed(input_fmap_32[15:0]) +
	( 15'sd 9078) * $signed(input_fmap_33[15:0]) +
	( 16'sd 21472) * $signed(input_fmap_34[15:0]) +
	( 16'sd 24670) * $signed(input_fmap_35[15:0]) +
	( 15'sd 14879) * $signed(input_fmap_36[15:0]) +
	( 14'sd 7774) * $signed(input_fmap_37[15:0]) +
	( 14'sd 7797) * $signed(input_fmap_38[15:0]) +
	( 16'sd 17252) * $signed(input_fmap_39[15:0]) +
	( 16'sd 27940) * $signed(input_fmap_40[15:0]) +
	( 16'sd 23999) * $signed(input_fmap_41[15:0]) +
	( 14'sd 7894) * $signed(input_fmap_42[15:0]) +
	( 13'sd 2831) * $signed(input_fmap_43[15:0]) +
	( 16'sd 25677) * $signed(input_fmap_44[15:0]) +
	( 15'sd 9388) * $signed(input_fmap_45[15:0]) +
	( 15'sd 13539) * $signed(input_fmap_46[15:0]) +
	( 16'sd 18326) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13031) * $signed(input_fmap_48[15:0]) +
	( 16'sd 25958) * $signed(input_fmap_49[15:0]) +
	( 16'sd 31907) * $signed(input_fmap_50[15:0]) +
	( 16'sd 22264) * $signed(input_fmap_51[15:0]) +
	( 15'sd 15461) * $signed(input_fmap_52[15:0]) +
	( 15'sd 10563) * $signed(input_fmap_53[15:0]) +
	( 14'sd 5881) * $signed(input_fmap_54[15:0]) +
	( 15'sd 14489) * $signed(input_fmap_55[15:0]) +
	( 15'sd 10868) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17713) * $signed(input_fmap_57[15:0]) +
	( 16'sd 27051) * $signed(input_fmap_58[15:0]) +
	( 14'sd 4363) * $signed(input_fmap_59[15:0]) +
	( 15'sd 11870) * $signed(input_fmap_60[15:0]) +
	( 16'sd 26120) * $signed(input_fmap_61[15:0]) +
	( 16'sd 19689) * $signed(input_fmap_62[15:0]) +
	( 13'sd 3996) * $signed(input_fmap_63[15:0]) +
	( 14'sd 6262) * $signed(input_fmap_64[15:0]) +
	( 15'sd 14576) * $signed(input_fmap_65[15:0]) +
	( 15'sd 9204) * $signed(input_fmap_66[15:0]) +
	( 10'sd 508) * $signed(input_fmap_67[15:0]) +
	( 16'sd 31624) * $signed(input_fmap_68[15:0]) +
	( 14'sd 4678) * $signed(input_fmap_69[15:0]) +
	( 14'sd 5859) * $signed(input_fmap_70[15:0]) +
	( 16'sd 30555) * $signed(input_fmap_71[15:0]) +
	( 15'sd 9633) * $signed(input_fmap_72[15:0]) +
	( 12'sd 1085) * $signed(input_fmap_73[15:0]) +
	( 16'sd 31670) * $signed(input_fmap_74[15:0]) +
	( 15'sd 12024) * $signed(input_fmap_75[15:0]) +
	( 16'sd 27751) * $signed(input_fmap_76[15:0]) +
	( 16'sd 29532) * $signed(input_fmap_77[15:0]) +
	( 15'sd 15051) * $signed(input_fmap_78[15:0]) +
	( 16'sd 20309) * $signed(input_fmap_79[15:0]) +
	( 16'sd 18546) * $signed(input_fmap_80[15:0]) +
	( 14'sd 6986) * $signed(input_fmap_81[15:0]) +
	( 10'sd 306) * $signed(input_fmap_82[15:0]) +
	( 16'sd 19703) * $signed(input_fmap_83[15:0]) +
	( 16'sd 27539) * $signed(input_fmap_84[15:0]) +
	( 14'sd 5194) * $signed(input_fmap_85[15:0]) +
	( 16'sd 23759) * $signed(input_fmap_86[15:0]) +
	( 16'sd 24066) * $signed(input_fmap_87[15:0]) +
	( 16'sd 28477) * $signed(input_fmap_88[15:0]) +
	( 14'sd 8153) * $signed(input_fmap_89[15:0]) +
	( 16'sd 27607) * $signed(input_fmap_90[15:0]) +
	( 12'sd 1898) * $signed(input_fmap_91[15:0]) +
	( 16'sd 21985) * $signed(input_fmap_92[15:0]) +
	( 16'sd 28232) * $signed(input_fmap_93[15:0]) +
	( 14'sd 6772) * $signed(input_fmap_94[15:0]) +
	( 16'sd 28251) * $signed(input_fmap_95[15:0]) +
	( 16'sd 25171) * $signed(input_fmap_96[15:0]) +
	( 16'sd 22442) * $signed(input_fmap_97[15:0]) +
	( 16'sd 19623) * $signed(input_fmap_98[15:0]) +
	( 16'sd 23159) * $signed(input_fmap_99[15:0]) +
	( 15'sd 8362) * $signed(input_fmap_100[15:0]) +
	( 16'sd 21678) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5664) * $signed(input_fmap_102[15:0]) +
	( 15'sd 14856) * $signed(input_fmap_103[15:0]) +
	( 12'sd 1543) * $signed(input_fmap_104[15:0]) +
	( 16'sd 18067) * $signed(input_fmap_105[15:0]) +
	( 16'sd 24311) * $signed(input_fmap_106[15:0]) +
	( 15'sd 15291) * $signed(input_fmap_107[15:0]) +
	( 15'sd 13490) * $signed(input_fmap_108[15:0]) +
	( 15'sd 12630) * $signed(input_fmap_109[15:0]) +
	( 15'sd 10989) * $signed(input_fmap_110[15:0]) +
	( 15'sd 12706) * $signed(input_fmap_111[15:0]) +
	( 16'sd 18575) * $signed(input_fmap_112[15:0]) +
	( 15'sd 15412) * $signed(input_fmap_113[15:0]) +
	( 16'sd 30170) * $signed(input_fmap_114[15:0]) +
	( 16'sd 24368) * $signed(input_fmap_115[15:0]) +
	( 16'sd 22713) * $signed(input_fmap_116[15:0]) +
	( 13'sd 3158) * $signed(input_fmap_117[15:0]) +
	( 15'sd 9609) * $signed(input_fmap_118[15:0]) +
	( 16'sd 27279) * $signed(input_fmap_119[15:0]) +
	( 15'sd 10494) * $signed(input_fmap_120[15:0]) +
	( 16'sd 17064) * $signed(input_fmap_121[15:0]) +
	( 16'sd 21508) * $signed(input_fmap_122[15:0]) +
	( 10'sd 437) * $signed(input_fmap_123[15:0]) +
	( 16'sd 19583) * $signed(input_fmap_124[15:0]) +
	( 13'sd 2392) * $signed(input_fmap_125[15:0]) +
	( 14'sd 4527) * $signed(input_fmap_126[15:0]) +
	( 15'sd 12433) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 13'sd 3655) * $signed(input_fmap_0[15:0]) +
	( 15'sd 15982) * $signed(input_fmap_1[15:0]) +
	( 15'sd 13429) * $signed(input_fmap_2[15:0]) +
	( 13'sd 3583) * $signed(input_fmap_3[15:0]) +
	( 16'sd 32391) * $signed(input_fmap_4[15:0]) +
	( 16'sd 19845) * $signed(input_fmap_5[15:0]) +
	( 16'sd 29821) * $signed(input_fmap_6[15:0]) +
	( 15'sd 12407) * $signed(input_fmap_7[15:0]) +
	( 12'sd 1692) * $signed(input_fmap_8[15:0]) +
	( 13'sd 2750) * $signed(input_fmap_9[15:0]) +
	( 16'sd 30911) * $signed(input_fmap_10[15:0]) +
	( 16'sd 27275) * $signed(input_fmap_11[15:0]) +
	( 15'sd 9478) * $signed(input_fmap_12[15:0]) +
	( 14'sd 6045) * $signed(input_fmap_13[15:0]) +
	( 16'sd 28411) * $signed(input_fmap_14[15:0]) +
	( 16'sd 17590) * $signed(input_fmap_15[15:0]) +
	( 16'sd 20725) * $signed(input_fmap_16[15:0]) +
	( 16'sd 27292) * $signed(input_fmap_17[15:0]) +
	( 14'sd 6576) * $signed(input_fmap_18[15:0]) +
	( 15'sd 10996) * $signed(input_fmap_19[15:0]) +
	( 12'sd 1649) * $signed(input_fmap_20[15:0]) +
	( 16'sd 28580) * $signed(input_fmap_21[15:0]) +
	( 15'sd 14724) * $signed(input_fmap_22[15:0]) +
	( 15'sd 14886) * $signed(input_fmap_23[15:0]) +
	( 15'sd 10212) * $signed(input_fmap_24[15:0]) +
	( 16'sd 25032) * $signed(input_fmap_25[15:0]) +
	( 16'sd 24929) * $signed(input_fmap_26[15:0]) +
	( 14'sd 5978) * $signed(input_fmap_27[15:0]) +
	( 13'sd 3913) * $signed(input_fmap_28[15:0]) +
	( 15'sd 11902) * $signed(input_fmap_29[15:0]) +
	( 16'sd 19641) * $signed(input_fmap_30[15:0]) +
	( 16'sd 17409) * $signed(input_fmap_31[15:0]) +
	( 15'sd 8410) * $signed(input_fmap_32[15:0]) +
	( 16'sd 30368) * $signed(input_fmap_33[15:0]) +
	( 16'sd 25190) * $signed(input_fmap_34[15:0]) +
	( 16'sd 23223) * $signed(input_fmap_35[15:0]) +
	( 16'sd 28430) * $signed(input_fmap_36[15:0]) +
	( 16'sd 17721) * $signed(input_fmap_37[15:0]) +
	( 16'sd 24524) * $signed(input_fmap_38[15:0]) +
	( 16'sd 31258) * $signed(input_fmap_39[15:0]) +
	( 16'sd 24779) * $signed(input_fmap_40[15:0]) +
	( 16'sd 20693) * $signed(input_fmap_41[15:0]) +
	( 15'sd 10200) * $signed(input_fmap_42[15:0]) +
	( 16'sd 20778) * $signed(input_fmap_43[15:0]) +
	( 16'sd 28442) * $signed(input_fmap_44[15:0]) +
	( 15'sd 15800) * $signed(input_fmap_45[15:0]) +
	( 16'sd 24782) * $signed(input_fmap_46[15:0]) +
	( 16'sd 22362) * $signed(input_fmap_47[15:0]) +
	( 16'sd 29725) * $signed(input_fmap_48[15:0]) +
	( 15'sd 13042) * $signed(input_fmap_49[15:0]) +
	( 16'sd 30053) * $signed(input_fmap_50[15:0]) +
	( 16'sd 27265) * $signed(input_fmap_51[15:0]) +
	( 16'sd 26003) * $signed(input_fmap_52[15:0]) +
	( 16'sd 19568) * $signed(input_fmap_53[15:0]) +
	( 15'sd 14865) * $signed(input_fmap_54[15:0]) +
	( 14'sd 7821) * $signed(input_fmap_55[15:0]) +
	( 16'sd 28806) * $signed(input_fmap_56[15:0]) +
	( 15'sd 9738) * $signed(input_fmap_57[15:0]) +
	( 14'sd 6696) * $signed(input_fmap_58[15:0]) +
	( 16'sd 27706) * $signed(input_fmap_59[15:0]) +
	( 16'sd 24470) * $signed(input_fmap_60[15:0]) +
	( 16'sd 30694) * $signed(input_fmap_61[15:0]) +
	( 15'sd 11965) * $signed(input_fmap_62[15:0]) +
	( 14'sd 4393) * $signed(input_fmap_63[15:0]) +
	( 16'sd 26849) * $signed(input_fmap_64[15:0]) +
	( 16'sd 31362) * $signed(input_fmap_65[15:0]) +
	( 14'sd 5907) * $signed(input_fmap_66[15:0]) +
	( 11'sd 521) * $signed(input_fmap_67[15:0]) +
	( 14'sd 4816) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31624) * $signed(input_fmap_69[15:0]) +
	( 14'sd 6068) * $signed(input_fmap_70[15:0]) +
	( 16'sd 23088) * $signed(input_fmap_71[15:0]) +
	( 16'sd 21223) * $signed(input_fmap_72[15:0]) +
	( 16'sd 30675) * $signed(input_fmap_73[15:0]) +
	( 14'sd 6700) * $signed(input_fmap_74[15:0]) +
	( 12'sd 1697) * $signed(input_fmap_75[15:0]) +
	( 16'sd 26491) * $signed(input_fmap_76[15:0]) +
	( 15'sd 14299) * $signed(input_fmap_77[15:0]) +
	( 15'sd 13449) * $signed(input_fmap_78[15:0]) +
	( 15'sd 10048) * $signed(input_fmap_79[15:0]) +
	( 15'sd 13848) * $signed(input_fmap_80[15:0]) +
	( 16'sd 22325) * $signed(input_fmap_81[15:0]) +
	( 16'sd 30775) * $signed(input_fmap_82[15:0]) +
	( 15'sd 15259) * $signed(input_fmap_83[15:0]) +
	( 16'sd 26100) * $signed(input_fmap_84[15:0]) +
	( 14'sd 4702) * $signed(input_fmap_85[15:0]) +
	( 15'sd 11048) * $signed(input_fmap_86[15:0]) +
	( 14'sd 6331) * $signed(input_fmap_87[15:0]) +
	( 16'sd 28435) * $signed(input_fmap_88[15:0]) +
	( 13'sd 3415) * $signed(input_fmap_89[15:0]) +
	( 16'sd 16842) * $signed(input_fmap_90[15:0]) +
	( 13'sd 3611) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25806) * $signed(input_fmap_92[15:0]) +
	( 14'sd 4106) * $signed(input_fmap_93[15:0]) +
	( 16'sd 20842) * $signed(input_fmap_94[15:0]) +
	( 15'sd 8214) * $signed(input_fmap_95[15:0]) +
	( 16'sd 20195) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27683) * $signed(input_fmap_97[15:0]) +
	( 16'sd 24965) * $signed(input_fmap_98[15:0]) +
	( 16'sd 24186) * $signed(input_fmap_99[15:0]) +
	( 15'sd 13620) * $signed(input_fmap_100[15:0]) +
	( 15'sd 12826) * $signed(input_fmap_101[15:0]) +
	( 16'sd 26213) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28320) * $signed(input_fmap_103[15:0]) +
	( 14'sd 6681) * $signed(input_fmap_104[15:0]) +
	( 15'sd 13126) * $signed(input_fmap_105[15:0]) +
	( 16'sd 24120) * $signed(input_fmap_106[15:0]) +
	( 16'sd 22814) * $signed(input_fmap_107[15:0]) +
	( 16'sd 16415) * $signed(input_fmap_108[15:0]) +
	( 16'sd 28366) * $signed(input_fmap_109[15:0]) +
	( 16'sd 25182) * $signed(input_fmap_110[15:0]) +
	( 15'sd 10511) * $signed(input_fmap_111[15:0]) +
	( 14'sd 6250) * $signed(input_fmap_112[15:0]) +
	( 16'sd 22763) * $signed(input_fmap_113[15:0]) +
	( 16'sd 18219) * $signed(input_fmap_114[15:0]) +
	( 16'sd 25703) * $signed(input_fmap_115[15:0]) +
	( 13'sd 2428) * $signed(input_fmap_116[15:0]) +
	( 16'sd 25108) * $signed(input_fmap_117[15:0]) +
	( 16'sd 23378) * $signed(input_fmap_118[15:0]) +
	( 16'sd 29951) * $signed(input_fmap_119[15:0]) +
	( 16'sd 30160) * $signed(input_fmap_120[15:0]) +
	( 15'sd 9300) * $signed(input_fmap_121[15:0]) +
	( 16'sd 17166) * $signed(input_fmap_122[15:0]) +
	( 16'sd 29675) * $signed(input_fmap_123[15:0]) +
	( 16'sd 17848) * $signed(input_fmap_124[15:0]) +
	( 14'sd 5624) * $signed(input_fmap_125[15:0]) +
	( 16'sd 23072) * $signed(input_fmap_126[15:0]) +
	( 16'sd 17402) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 15'sd 12802) * $signed(input_fmap_0[15:0]) +
	( 16'sd 22958) * $signed(input_fmap_1[15:0]) +
	( 15'sd 13070) * $signed(input_fmap_2[15:0]) +
	( 15'sd 9435) * $signed(input_fmap_3[15:0]) +
	( 14'sd 6324) * $signed(input_fmap_4[15:0]) +
	( 16'sd 30032) * $signed(input_fmap_5[15:0]) +
	( 16'sd 17879) * $signed(input_fmap_6[15:0]) +
	( 16'sd 26010) * $signed(input_fmap_7[15:0]) +
	( 16'sd 19955) * $signed(input_fmap_8[15:0]) +
	( 16'sd 30564) * $signed(input_fmap_9[15:0]) +
	( 15'sd 16371) * $signed(input_fmap_10[15:0]) +
	( 13'sd 4063) * $signed(input_fmap_11[15:0]) +
	( 16'sd 24759) * $signed(input_fmap_12[15:0]) +
	( 16'sd 30537) * $signed(input_fmap_13[15:0]) +
	( 15'sd 11431) * $signed(input_fmap_14[15:0]) +
	( 15'sd 10872) * $signed(input_fmap_15[15:0]) +
	( 16'sd 30380) * $signed(input_fmap_16[15:0]) +
	( 16'sd 27786) * $signed(input_fmap_17[15:0]) +
	( 15'sd 12223) * $signed(input_fmap_18[15:0]) +
	( 15'sd 10343) * $signed(input_fmap_19[15:0]) +
	( 15'sd 8921) * $signed(input_fmap_20[15:0]) +
	( 16'sd 18251) * $signed(input_fmap_21[15:0]) +
	( 16'sd 19730) * $signed(input_fmap_22[15:0]) +
	( 16'sd 32511) * $signed(input_fmap_23[15:0]) +
	( 15'sd 8583) * $signed(input_fmap_24[15:0]) +
	( 16'sd 17320) * $signed(input_fmap_25[15:0]) +
	( 16'sd 20066) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9207) * $signed(input_fmap_27[15:0]) +
	( 15'sd 8814) * $signed(input_fmap_28[15:0]) +
	( 16'sd 31260) * $signed(input_fmap_29[15:0]) +
	( 14'sd 4902) * $signed(input_fmap_30[15:0]) +
	( 14'sd 5331) * $signed(input_fmap_31[15:0]) +
	( 16'sd 27389) * $signed(input_fmap_32[15:0]) +
	( 16'sd 32061) * $signed(input_fmap_33[15:0]) +
	( 16'sd 22187) * $signed(input_fmap_34[15:0]) +
	( 15'sd 12598) * $signed(input_fmap_35[15:0]) +
	( 16'sd 23547) * $signed(input_fmap_36[15:0]) +
	( 16'sd 24827) * $signed(input_fmap_37[15:0]) +
	( 15'sd 8260) * $signed(input_fmap_38[15:0]) +
	( 16'sd 18583) * $signed(input_fmap_39[15:0]) +
	( 16'sd 29751) * $signed(input_fmap_40[15:0]) +
	( 16'sd 28433) * $signed(input_fmap_41[15:0]) +
	( 16'sd 21980) * $signed(input_fmap_42[15:0]) +
	( 12'sd 1149) * $signed(input_fmap_43[15:0]) +
	( 15'sd 8796) * $signed(input_fmap_44[15:0]) +
	( 16'sd 20177) * $signed(input_fmap_45[15:0]) +
	( 16'sd 18589) * $signed(input_fmap_46[15:0]) +
	( 12'sd 1973) * $signed(input_fmap_47[15:0]) +
	( 16'sd 24416) * $signed(input_fmap_48[15:0]) +
	( 15'sd 10598) * $signed(input_fmap_49[15:0]) +
	( 15'sd 10028) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15112) * $signed(input_fmap_51[15:0]) +
	( 15'sd 14420) * $signed(input_fmap_52[15:0]) +
	( 16'sd 20015) * $signed(input_fmap_53[15:0]) +
	( 15'sd 14764) * $signed(input_fmap_54[15:0]) +
	( 15'sd 10007) * $signed(input_fmap_55[15:0]) +
	( 16'sd 24904) * $signed(input_fmap_56[15:0]) +
	( 16'sd 24386) * $signed(input_fmap_57[15:0]) +
	( 15'sd 9365) * $signed(input_fmap_58[15:0]) +
	( 16'sd 26041) * $signed(input_fmap_59[15:0]) +
	( 16'sd 24103) * $signed(input_fmap_60[15:0]) +
	( 16'sd 23577) * $signed(input_fmap_61[15:0]) +
	( 15'sd 15892) * $signed(input_fmap_62[15:0]) +
	( 15'sd 14915) * $signed(input_fmap_63[15:0]) +
	( 12'sd 1951) * $signed(input_fmap_64[15:0]) +
	( 16'sd 29354) * $signed(input_fmap_65[15:0]) +
	( 13'sd 3881) * $signed(input_fmap_66[15:0]) +
	( 12'sd 1446) * $signed(input_fmap_67[15:0]) +
	( 16'sd 22922) * $signed(input_fmap_68[15:0]) +
	( 16'sd 25477) * $signed(input_fmap_69[15:0]) +
	( 15'sd 9938) * $signed(input_fmap_70[15:0]) +
	( 16'sd 26898) * $signed(input_fmap_71[15:0]) +
	( 16'sd 21153) * $signed(input_fmap_72[15:0]) +
	( 16'sd 31018) * $signed(input_fmap_73[15:0]) +
	( 15'sd 16198) * $signed(input_fmap_74[15:0]) +
	( 15'sd 15898) * $signed(input_fmap_75[15:0]) +
	( 16'sd 21085) * $signed(input_fmap_76[15:0]) +
	( 15'sd 15441) * $signed(input_fmap_77[15:0]) +
	( 16'sd 26288) * $signed(input_fmap_78[15:0]) +
	( 12'sd 1886) * $signed(input_fmap_79[15:0]) +
	( 16'sd 23004) * $signed(input_fmap_80[15:0]) +
	( 15'sd 11682) * $signed(input_fmap_81[15:0]) +
	( 16'sd 21651) * $signed(input_fmap_82[15:0]) +
	( 16'sd 30903) * $signed(input_fmap_83[15:0]) +
	( 16'sd 30468) * $signed(input_fmap_84[15:0]) +
	( 16'sd 17470) * $signed(input_fmap_85[15:0]) +
	( 15'sd 8672) * $signed(input_fmap_86[15:0]) +
	( 16'sd 31333) * $signed(input_fmap_87[15:0]) +
	( 15'sd 14157) * $signed(input_fmap_88[15:0]) +
	( 13'sd 2674) * $signed(input_fmap_89[15:0]) +
	( 16'sd 17060) * $signed(input_fmap_90[15:0]) +
	( 16'sd 31863) * $signed(input_fmap_91[15:0]) +
	( 15'sd 11180) * $signed(input_fmap_92[15:0]) +
	( 16'sd 22112) * $signed(input_fmap_93[15:0]) +
	( 14'sd 6398) * $signed(input_fmap_94[15:0]) +
	( 16'sd 27991) * $signed(input_fmap_95[15:0]) +
	( 16'sd 27153) * $signed(input_fmap_96[15:0]) +
	( 15'sd 10347) * $signed(input_fmap_97[15:0]) +
	( 15'sd 12644) * $signed(input_fmap_98[15:0]) +
	( 16'sd 18108) * $signed(input_fmap_99[15:0]) +
	( 16'sd 17710) * $signed(input_fmap_100[15:0]) +
	( 16'sd 24278) * $signed(input_fmap_101[15:0]) +
	( 16'sd 23769) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28276) * $signed(input_fmap_103[15:0]) +
	( 14'sd 7573) * $signed(input_fmap_104[15:0]) +
	( 16'sd 25456) * $signed(input_fmap_105[15:0]) +
	( 16'sd 29672) * $signed(input_fmap_106[15:0]) +
	( 16'sd 31034) * $signed(input_fmap_107[15:0]) +
	( 16'sd 26548) * $signed(input_fmap_108[15:0]) +
	( 16'sd 22179) * $signed(input_fmap_109[15:0]) +
	( 16'sd 31393) * $signed(input_fmap_110[15:0]) +
	( 13'sd 3075) * $signed(input_fmap_111[15:0]) +
	( 16'sd 30340) * $signed(input_fmap_112[15:0]) +
	( 16'sd 19772) * $signed(input_fmap_113[15:0]) +
	( 9'sd 204) * $signed(input_fmap_114[15:0]) +
	( 13'sd 3438) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26210) * $signed(input_fmap_116[15:0]) +
	( 15'sd 14439) * $signed(input_fmap_117[15:0]) +
	( 16'sd 18588) * $signed(input_fmap_118[15:0]) +
	( 16'sd 21091) * $signed(input_fmap_119[15:0]) +
	( 13'sd 3098) * $signed(input_fmap_120[15:0]) +
	( 15'sd 12700) * $signed(input_fmap_121[15:0]) +
	( 16'sd 27133) * $signed(input_fmap_122[15:0]) +
	( 12'sd 1790) * $signed(input_fmap_123[15:0]) +
	( 15'sd 13059) * $signed(input_fmap_124[15:0]) +
	( 16'sd 28973) * $signed(input_fmap_125[15:0]) +
	( 16'sd 25682) * $signed(input_fmap_126[15:0]) +
	( 13'sd 2827) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 16'sd 20350) * $signed(input_fmap_0[15:0]) +
	( 15'sd 12976) * $signed(input_fmap_1[15:0]) +
	( 16'sd 31835) * $signed(input_fmap_2[15:0]) +
	( 15'sd 14000) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30737) * $signed(input_fmap_4[15:0]) +
	( 11'sd 551) * $signed(input_fmap_5[15:0]) +
	( 14'sd 4951) * $signed(input_fmap_6[15:0]) +
	( 16'sd 30164) * $signed(input_fmap_7[15:0]) +
	( 16'sd 24045) * $signed(input_fmap_8[15:0]) +
	( 15'sd 10890) * $signed(input_fmap_9[15:0]) +
	( 16'sd 17620) * $signed(input_fmap_10[15:0]) +
	( 15'sd 14320) * $signed(input_fmap_11[15:0]) +
	( 14'sd 4399) * $signed(input_fmap_12[15:0]) +
	( 16'sd 22290) * $signed(input_fmap_13[15:0]) +
	( 16'sd 28837) * $signed(input_fmap_14[15:0]) +
	( 14'sd 5805) * $signed(input_fmap_15[15:0]) +
	( 14'sd 7044) * $signed(input_fmap_16[15:0]) +
	( 13'sd 4007) * $signed(input_fmap_17[15:0]) +
	( 16'sd 25107) * $signed(input_fmap_18[15:0]) +
	( 15'sd 13903) * $signed(input_fmap_19[15:0]) +
	( 14'sd 6785) * $signed(input_fmap_20[15:0]) +
	( 16'sd 23546) * $signed(input_fmap_21[15:0]) +
	( 16'sd 23498) * $signed(input_fmap_22[15:0]) +
	( 15'sd 14243) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17219) * $signed(input_fmap_24[15:0]) +
	( 16'sd 16837) * $signed(input_fmap_25[15:0]) +
	( 15'sd 14520) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2443) * $signed(input_fmap_27[15:0]) +
	( 16'sd 27805) * $signed(input_fmap_28[15:0]) +
	( 15'sd 8656) * $signed(input_fmap_29[15:0]) +
	( 15'sd 10633) * $signed(input_fmap_30[15:0]) +
	( 16'sd 22973) * $signed(input_fmap_31[15:0]) +
	( 16'sd 18645) * $signed(input_fmap_32[15:0]) +
	( 13'sd 2799) * $signed(input_fmap_33[15:0]) +
	( 11'sd 714) * $signed(input_fmap_34[15:0]) +
	( 16'sd 25323) * $signed(input_fmap_35[15:0]) +
	( 16'sd 25902) * $signed(input_fmap_36[15:0]) +
	( 16'sd 32213) * $signed(input_fmap_37[15:0]) +
	( 11'sd 1011) * $signed(input_fmap_38[15:0]) +
	( 13'sd 2197) * $signed(input_fmap_39[15:0]) +
	( 15'sd 13689) * $signed(input_fmap_40[15:0]) +
	( 15'sd 11138) * $signed(input_fmap_41[15:0]) +
	( 16'sd 17789) * $signed(input_fmap_42[15:0]) +
	( 15'sd 14682) * $signed(input_fmap_43[15:0]) +
	( 14'sd 5328) * $signed(input_fmap_44[15:0]) +
	( 12'sd 1765) * $signed(input_fmap_45[15:0]) +
	( 13'sd 3389) * $signed(input_fmap_46[15:0]) +
	( 16'sd 17795) * $signed(input_fmap_47[15:0]) +
	( 13'sd 2359) * $signed(input_fmap_48[15:0]) +
	( 16'sd 24676) * $signed(input_fmap_49[15:0]) +
	( 16'sd 30957) * $signed(input_fmap_50[15:0]) +
	( 16'sd 27472) * $signed(input_fmap_51[15:0]) +
	( 16'sd 32735) * $signed(input_fmap_52[15:0]) +
	( 15'sd 10153) * $signed(input_fmap_53[15:0]) +
	( 16'sd 29713) * $signed(input_fmap_54[15:0]) +
	( 16'sd 32171) * $signed(input_fmap_55[15:0]) +
	( 16'sd 17534) * $signed(input_fmap_56[15:0]) +
	( 15'sd 10380) * $signed(input_fmap_57[15:0]) +
	( 16'sd 30297) * $signed(input_fmap_58[15:0]) +
	( 16'sd 20114) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1992) * $signed(input_fmap_60[15:0]) +
	( 15'sd 10638) * $signed(input_fmap_61[15:0]) +
	( 15'sd 15783) * $signed(input_fmap_62[15:0]) +
	( 16'sd 29352) * $signed(input_fmap_63[15:0]) +
	( 15'sd 13519) * $signed(input_fmap_64[15:0]) +
	( 16'sd 31810) * $signed(input_fmap_65[15:0]) +
	( 16'sd 29989) * $signed(input_fmap_66[15:0]) +
	( 16'sd 27660) * $signed(input_fmap_67[15:0]) +
	( 15'sd 14682) * $signed(input_fmap_68[15:0]) +
	( 16'sd 30123) * $signed(input_fmap_69[15:0]) +
	( 13'sd 2884) * $signed(input_fmap_70[15:0]) +
	( 13'sd 2503) * $signed(input_fmap_71[15:0]) +
	( 16'sd 28316) * $signed(input_fmap_72[15:0]) +
	( 16'sd 30202) * $signed(input_fmap_73[15:0]) +
	( 10'sd 318) * $signed(input_fmap_74[15:0]) +
	( 14'sd 5719) * $signed(input_fmap_75[15:0]) +
	( 16'sd 18795) * $signed(input_fmap_76[15:0]) +
	( 14'sd 7531) * $signed(input_fmap_77[15:0]) +
	( 16'sd 32672) * $signed(input_fmap_78[15:0]) +
	( 15'sd 8965) * $signed(input_fmap_79[15:0]) +
	( 15'sd 11943) * $signed(input_fmap_80[15:0]) +
	( 16'sd 25076) * $signed(input_fmap_81[15:0]) +
	( 16'sd 20911) * $signed(input_fmap_82[15:0]) +
	( 14'sd 7555) * $signed(input_fmap_83[15:0]) +
	( 15'sd 10756) * $signed(input_fmap_84[15:0]) +
	( 16'sd 27331) * $signed(input_fmap_85[15:0]) +
	( 14'sd 7109) * $signed(input_fmap_86[15:0]) +
	( 16'sd 21037) * $signed(input_fmap_87[15:0]) +
	( 15'sd 14172) * $signed(input_fmap_88[15:0]) +
	( 16'sd 17790) * $signed(input_fmap_89[15:0]) +
	( 16'sd 18970) * $signed(input_fmap_90[15:0]) +
	( 16'sd 20909) * $signed(input_fmap_91[15:0]) +
	( 15'sd 9506) * $signed(input_fmap_92[15:0]) +
	( 15'sd 12051) * $signed(input_fmap_93[15:0]) +
	( 16'sd 28950) * $signed(input_fmap_94[15:0]) +
	( 15'sd 14320) * $signed(input_fmap_95[15:0]) +
	( 16'sd 18038) * $signed(input_fmap_96[15:0]) +
	( 15'sd 11507) * $signed(input_fmap_97[15:0]) +
	( 15'sd 13102) * $signed(input_fmap_98[15:0]) +
	( 14'sd 5290) * $signed(input_fmap_99[15:0]) +
	( 15'sd 14818) * $signed(input_fmap_100[15:0]) +
	( 16'sd 23672) * $signed(input_fmap_101[15:0]) +
	( 15'sd 9895) * $signed(input_fmap_102[15:0]) +
	( 16'sd 26492) * $signed(input_fmap_103[15:0]) +
	( 15'sd 13449) * $signed(input_fmap_104[15:0]) +
	( 12'sd 1123) * $signed(input_fmap_105[15:0]) +
	( 16'sd 19169) * $signed(input_fmap_106[15:0]) +
	( 16'sd 32509) * $signed(input_fmap_107[15:0]) +
	( 16'sd 22030) * $signed(input_fmap_108[15:0]) +
	( 16'sd 23511) * $signed(input_fmap_109[15:0]) +
	( 14'sd 7927) * $signed(input_fmap_110[15:0]) +
	( 16'sd 21822) * $signed(input_fmap_111[15:0]) +
	( 14'sd 7021) * $signed(input_fmap_112[15:0]) +
	( 16'sd 25835) * $signed(input_fmap_113[15:0]) +
	( 16'sd 16734) * $signed(input_fmap_114[15:0]) +
	( 14'sd 6567) * $signed(input_fmap_115[15:0]) +
	( 16'sd 23764) * $signed(input_fmap_116[15:0]) +
	( 15'sd 9684) * $signed(input_fmap_117[15:0]) +
	( 16'sd 20194) * $signed(input_fmap_118[15:0]) +
	( 16'sd 29053) * $signed(input_fmap_119[15:0]) +
	( 14'sd 8161) * $signed(input_fmap_120[15:0]) +
	( 16'sd 17138) * $signed(input_fmap_121[15:0]) +
	( 16'sd 22708) * $signed(input_fmap_122[15:0]) +
	( 16'sd 27921) * $signed(input_fmap_123[15:0]) +
	( 16'sd 20795) * $signed(input_fmap_124[15:0]) +
	( 15'sd 12763) * $signed(input_fmap_125[15:0]) +
	( 16'sd 22146) * $signed(input_fmap_126[15:0]) +
	( 14'sd 5700) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 15'sd 8658) * $signed(input_fmap_0[15:0]) +
	( 14'sd 6291) * $signed(input_fmap_1[15:0]) +
	( 16'sd 22335) * $signed(input_fmap_2[15:0]) +
	( 15'sd 13540) * $signed(input_fmap_3[15:0]) +
	( 16'sd 18605) * $signed(input_fmap_4[15:0]) +
	( 15'sd 11603) * $signed(input_fmap_5[15:0]) +
	( 16'sd 25061) * $signed(input_fmap_6[15:0]) +
	( 16'sd 32750) * $signed(input_fmap_7[15:0]) +
	( 14'sd 6443) * $signed(input_fmap_8[15:0]) +
	( 16'sd 28929) * $signed(input_fmap_9[15:0]) +
	( 16'sd 25576) * $signed(input_fmap_10[15:0]) +
	( 16'sd 23893) * $signed(input_fmap_11[15:0]) +
	( 16'sd 24492) * $signed(input_fmap_12[15:0]) +
	( 13'sd 4053) * $signed(input_fmap_13[15:0]) +
	( 16'sd 28480) * $signed(input_fmap_14[15:0]) +
	( 16'sd 27639) * $signed(input_fmap_15[15:0]) +
	( 16'sd 16764) * $signed(input_fmap_16[15:0]) +
	( 16'sd 31295) * $signed(input_fmap_17[15:0]) +
	( 16'sd 30458) * $signed(input_fmap_18[15:0]) +
	( 16'sd 21726) * $signed(input_fmap_19[15:0]) +
	( 16'sd 21421) * $signed(input_fmap_20[15:0]) +
	( 15'sd 12026) * $signed(input_fmap_21[15:0]) +
	( 16'sd 18695) * $signed(input_fmap_22[15:0]) +
	( 14'sd 6335) * $signed(input_fmap_23[15:0]) +
	( 16'sd 26732) * $signed(input_fmap_24[15:0]) +
	( 16'sd 18243) * $signed(input_fmap_25[15:0]) +
	( 16'sd 18002) * $signed(input_fmap_26[15:0]) +
	( 2'sd 1) * $signed(input_fmap_27[15:0]) +
	( 16'sd 21309) * $signed(input_fmap_28[15:0]) +
	( 15'sd 15525) * $signed(input_fmap_29[15:0]) +
	( 16'sd 28498) * $signed(input_fmap_30[15:0]) +
	( 15'sd 10651) * $signed(input_fmap_31[15:0]) +
	( 16'sd 22765) * $signed(input_fmap_32[15:0]) +
	( 15'sd 13709) * $signed(input_fmap_33[15:0]) +
	( 11'sd 892) * $signed(input_fmap_34[15:0]) +
	( 16'sd 27931) * $signed(input_fmap_35[15:0]) +
	( 16'sd 28947) * $signed(input_fmap_36[15:0]) +
	( 11'sd 568) * $signed(input_fmap_37[15:0]) +
	( 12'sd 1327) * $signed(input_fmap_38[15:0]) +
	( 16'sd 29066) * $signed(input_fmap_39[15:0]) +
	( 16'sd 23691) * $signed(input_fmap_40[15:0]) +
	( 13'sd 2457) * $signed(input_fmap_41[15:0]) +
	( 16'sd 25828) * $signed(input_fmap_42[15:0]) +
	( 15'sd 9383) * $signed(input_fmap_43[15:0]) +
	( 12'sd 1359) * $signed(input_fmap_44[15:0]) +
	( 13'sd 2106) * $signed(input_fmap_45[15:0]) +
	( 16'sd 16586) * $signed(input_fmap_46[15:0]) +
	( 16'sd 29114) * $signed(input_fmap_47[15:0]) +
	( 14'sd 6915) * $signed(input_fmap_48[15:0]) +
	( 16'sd 22101) * $signed(input_fmap_49[15:0]) +
	( 13'sd 2148) * $signed(input_fmap_50[15:0]) +
	( 15'sd 12257) * $signed(input_fmap_51[15:0]) +
	( 15'sd 13899) * $signed(input_fmap_52[15:0]) +
	( 16'sd 22964) * $signed(input_fmap_53[15:0]) +
	( 15'sd 13963) * $signed(input_fmap_54[15:0]) +
	( 15'sd 12410) * $signed(input_fmap_55[15:0]) +
	( 16'sd 20597) * $signed(input_fmap_56[15:0]) +
	( 11'sd 512) * $signed(input_fmap_57[15:0]) +
	( 15'sd 9504) * $signed(input_fmap_58[15:0]) +
	( 16'sd 17285) * $signed(input_fmap_59[15:0]) +
	( 16'sd 27631) * $signed(input_fmap_60[15:0]) +
	( 15'sd 11676) * $signed(input_fmap_61[15:0]) +
	( 16'sd 28020) * $signed(input_fmap_62[15:0]) +
	( 16'sd 21062) * $signed(input_fmap_63[15:0]) +
	( 16'sd 26244) * $signed(input_fmap_64[15:0]) +
	( 12'sd 1078) * $signed(input_fmap_65[15:0]) +
	( 16'sd 30947) * $signed(input_fmap_66[15:0]) +
	( 16'sd 26341) * $signed(input_fmap_67[15:0]) +
	( 16'sd 23511) * $signed(input_fmap_68[15:0]) +
	( 15'sd 10279) * $signed(input_fmap_69[15:0]) +
	( 16'sd 27980) * $signed(input_fmap_70[15:0]) +
	( 16'sd 27353) * $signed(input_fmap_71[15:0]) +
	( 16'sd 22524) * $signed(input_fmap_72[15:0]) +
	( 14'sd 7472) * $signed(input_fmap_73[15:0]) +
	( 16'sd 25662) * $signed(input_fmap_74[15:0]) +
	( 16'sd 27724) * $signed(input_fmap_75[15:0]) +
	( 15'sd 12712) * $signed(input_fmap_76[15:0]) +
	( 16'sd 19407) * $signed(input_fmap_77[15:0]) +
	( 16'sd 27239) * $signed(input_fmap_78[15:0]) +
	( 15'sd 16314) * $signed(input_fmap_79[15:0]) +
	( 16'sd 24793) * $signed(input_fmap_80[15:0]) +
	( 15'sd 12723) * $signed(input_fmap_81[15:0]) +
	( 15'sd 10549) * $signed(input_fmap_82[15:0]) +
	( 15'sd 14792) * $signed(input_fmap_83[15:0]) +
	( 16'sd 25317) * $signed(input_fmap_84[15:0]) +
	( 16'sd 25064) * $signed(input_fmap_85[15:0]) +
	( 16'sd 17132) * $signed(input_fmap_86[15:0]) +
	( 15'sd 15940) * $signed(input_fmap_87[15:0]) +
	( 15'sd 13880) * $signed(input_fmap_88[15:0]) +
	( 14'sd 6626) * $signed(input_fmap_89[15:0]) +
	( 15'sd 14151) * $signed(input_fmap_90[15:0]) +
	( 15'sd 12736) * $signed(input_fmap_91[15:0]) +
	( 16'sd 23807) * $signed(input_fmap_92[15:0]) +
	( 16'sd 21170) * $signed(input_fmap_93[15:0]) +
	( 16'sd 18879) * $signed(input_fmap_94[15:0]) +
	( 15'sd 9127) * $signed(input_fmap_95[15:0]) +
	( 16'sd 28436) * $signed(input_fmap_96[15:0]) +
	( 15'sd 10896) * $signed(input_fmap_97[15:0]) +
	( 14'sd 4888) * $signed(input_fmap_98[15:0]) +
	( 16'sd 28131) * $signed(input_fmap_99[15:0]) +
	( 16'sd 19708) * $signed(input_fmap_100[15:0]) +
	( 14'sd 4945) * $signed(input_fmap_101[15:0]) +
	( 15'sd 11746) * $signed(input_fmap_102[15:0]) +
	( 16'sd 29098) * $signed(input_fmap_103[15:0]) +
	( 15'sd 15344) * $signed(input_fmap_104[15:0]) +
	( 16'sd 32003) * $signed(input_fmap_105[15:0]) +
	( 16'sd 30887) * $signed(input_fmap_106[15:0]) +
	( 16'sd 28004) * $signed(input_fmap_107[15:0]) +
	( 16'sd 27740) * $signed(input_fmap_108[15:0]) +
	( 16'sd 30668) * $signed(input_fmap_109[15:0]) +
	( 14'sd 5712) * $signed(input_fmap_110[15:0]) +
	( 15'sd 9905) * $signed(input_fmap_111[15:0]) +
	( 16'sd 27043) * $signed(input_fmap_112[15:0]) +
	( 16'sd 27440) * $signed(input_fmap_113[15:0]) +
	( 13'sd 3922) * $signed(input_fmap_114[15:0]) +
	( 15'sd 10757) * $signed(input_fmap_115[15:0]) +
	( 16'sd 31005) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27594) * $signed(input_fmap_117[15:0]) +
	( 16'sd 27771) * $signed(input_fmap_118[15:0]) +
	( 16'sd 17560) * $signed(input_fmap_119[15:0]) +
	( 16'sd 27986) * $signed(input_fmap_120[15:0]) +
	( 15'sd 12637) * $signed(input_fmap_121[15:0]) +
	( 16'sd 20839) * $signed(input_fmap_122[15:0]) +
	( 15'sd 15337) * $signed(input_fmap_123[15:0]) +
	( 15'sd 15695) * $signed(input_fmap_124[15:0]) +
	( 15'sd 14131) * $signed(input_fmap_125[15:0]) +
	( 16'sd 22604) * $signed(input_fmap_126[15:0]) +
	( 16'sd 30767) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 15'sd 11316) * $signed(input_fmap_0[15:0]) +
	( 14'sd 4648) * $signed(input_fmap_1[15:0]) +
	( 15'sd 13244) * $signed(input_fmap_2[15:0]) +
	( 16'sd 27672) * $signed(input_fmap_3[15:0]) +
	( 16'sd 20809) * $signed(input_fmap_4[15:0]) +
	( 16'sd 17390) * $signed(input_fmap_5[15:0]) +
	( 16'sd 18166) * $signed(input_fmap_6[15:0]) +
	( 15'sd 8474) * $signed(input_fmap_7[15:0]) +
	( 15'sd 15244) * $signed(input_fmap_8[15:0]) +
	( 15'sd 11720) * $signed(input_fmap_9[15:0]) +
	( 14'sd 4247) * $signed(input_fmap_10[15:0]) +
	( 14'sd 4563) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20899) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24646) * $signed(input_fmap_13[15:0]) +
	( 16'sd 30867) * $signed(input_fmap_14[15:0]) +
	( 16'sd 24797) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10514) * $signed(input_fmap_16[15:0]) +
	( 16'sd 21294) * $signed(input_fmap_17[15:0]) +
	( 14'sd 6623) * $signed(input_fmap_18[15:0]) +
	( 16'sd 25840) * $signed(input_fmap_19[15:0]) +
	( 15'sd 13730) * $signed(input_fmap_20[15:0]) +
	( 16'sd 21199) * $signed(input_fmap_21[15:0]) +
	( 16'sd 30000) * $signed(input_fmap_22[15:0]) +
	( 15'sd 10634) * $signed(input_fmap_23[15:0]) +
	( 15'sd 10113) * $signed(input_fmap_24[15:0]) +
	( 14'sd 4205) * $signed(input_fmap_25[15:0]) +
	( 16'sd 31863) * $signed(input_fmap_26[15:0]) +
	( 15'sd 10490) * $signed(input_fmap_27[15:0]) +
	( 10'sd 369) * $signed(input_fmap_28[15:0]) +
	( 16'sd 22498) * $signed(input_fmap_29[15:0]) +
	( 16'sd 24495) * $signed(input_fmap_30[15:0]) +
	( 16'sd 23451) * $signed(input_fmap_31[15:0]) +
	( 15'sd 12562) * $signed(input_fmap_32[15:0]) +
	( 16'sd 22337) * $signed(input_fmap_33[15:0]) +
	( 16'sd 27277) * $signed(input_fmap_34[15:0]) +
	( 14'sd 5299) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11179) * $signed(input_fmap_36[15:0]) +
	( 15'sd 13954) * $signed(input_fmap_37[15:0]) +
	( 16'sd 29491) * $signed(input_fmap_38[15:0]) +
	( 15'sd 14777) * $signed(input_fmap_39[15:0]) +
	( 14'sd 5841) * $signed(input_fmap_40[15:0]) +
	( 16'sd 29713) * $signed(input_fmap_41[15:0]) +
	( 16'sd 19585) * $signed(input_fmap_42[15:0]) +
	( 14'sd 6063) * $signed(input_fmap_43[15:0]) +
	( 15'sd 11038) * $signed(input_fmap_44[15:0]) +
	( 13'sd 2660) * $signed(input_fmap_45[15:0]) +
	( 13'sd 3112) * $signed(input_fmap_46[15:0]) +
	( 16'sd 17689) * $signed(input_fmap_47[15:0]) +
	( 16'sd 22759) * $signed(input_fmap_48[15:0]) +
	( 16'sd 23255) * $signed(input_fmap_49[15:0]) +
	( 16'sd 25204) * $signed(input_fmap_50[15:0]) +
	( 16'sd 32077) * $signed(input_fmap_51[15:0]) +
	( 14'sd 4634) * $signed(input_fmap_52[15:0]) +
	( 16'sd 25003) * $signed(input_fmap_53[15:0]) +
	( 16'sd 17351) * $signed(input_fmap_54[15:0]) +
	( 16'sd 16810) * $signed(input_fmap_55[15:0]) +
	( 13'sd 3590) * $signed(input_fmap_56[15:0]) +
	( 16'sd 18459) * $signed(input_fmap_57[15:0]) +
	( 15'sd 15818) * $signed(input_fmap_58[15:0]) +
	( 16'sd 32049) * $signed(input_fmap_59[15:0]) +
	( 16'sd 23846) * $signed(input_fmap_60[15:0]) +
	( 14'sd 8018) * $signed(input_fmap_61[15:0]) +
	( 11'sd 596) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20949) * $signed(input_fmap_63[15:0]) +
	( 16'sd 26460) * $signed(input_fmap_64[15:0]) +
	( 16'sd 19947) * $signed(input_fmap_65[15:0]) +
	( 16'sd 27887) * $signed(input_fmap_66[15:0]) +
	( 15'sd 8476) * $signed(input_fmap_67[15:0]) +
	( 12'sd 1629) * $signed(input_fmap_68[15:0]) +
	( 14'sd 6803) * $signed(input_fmap_69[15:0]) +
	( 16'sd 20641) * $signed(input_fmap_70[15:0]) +
	( 13'sd 2488) * $signed(input_fmap_71[15:0]) +
	( 13'sd 2668) * $signed(input_fmap_72[15:0]) +
	( 16'sd 31494) * $signed(input_fmap_73[15:0]) +
	( 14'sd 5641) * $signed(input_fmap_74[15:0]) +
	( 16'sd 18077) * $signed(input_fmap_75[15:0]) +
	( 15'sd 15673) * $signed(input_fmap_76[15:0]) +
	( 15'sd 15594) * $signed(input_fmap_77[15:0]) +
	( 16'sd 25571) * $signed(input_fmap_78[15:0]) +
	( 16'sd 30752) * $signed(input_fmap_79[15:0]) +
	( 15'sd 13133) * $signed(input_fmap_80[15:0]) +
	( 15'sd 9046) * $signed(input_fmap_81[15:0]) +
	( 16'sd 25575) * $signed(input_fmap_82[15:0]) +
	( 14'sd 4106) * $signed(input_fmap_83[15:0]) +
	( 16'sd 25054) * $signed(input_fmap_84[15:0]) +
	( 16'sd 32093) * $signed(input_fmap_85[15:0]) +
	( 16'sd 28259) * $signed(input_fmap_86[15:0]) +
	( 16'sd 18526) * $signed(input_fmap_87[15:0]) +
	( 16'sd 30909) * $signed(input_fmap_88[15:0]) +
	( 14'sd 6935) * $signed(input_fmap_89[15:0]) +
	( 11'sd 889) * $signed(input_fmap_90[15:0]) +
	( 16'sd 29647) * $signed(input_fmap_91[15:0]) +
	( 16'sd 17569) * $signed(input_fmap_92[15:0]) +
	( 15'sd 15339) * $signed(input_fmap_93[15:0]) +
	( 15'sd 14838) * $signed(input_fmap_94[15:0]) +
	( 15'sd 16024) * $signed(input_fmap_95[15:0]) +
	( 16'sd 24574) * $signed(input_fmap_96[15:0]) +
	( 16'sd 29880) * $signed(input_fmap_97[15:0]) +
	( 16'sd 19323) * $signed(input_fmap_98[15:0]) +
	( 14'sd 5897) * $signed(input_fmap_99[15:0]) +
	( 15'sd 13624) * $signed(input_fmap_100[15:0]) +
	( 16'sd 30677) * $signed(input_fmap_101[15:0]) +
	( 13'sd 2181) * $signed(input_fmap_102[15:0]) +
	( 15'sd 10725) * $signed(input_fmap_103[15:0]) +
	( 16'sd 17114) * $signed(input_fmap_104[15:0]) +
	( 10'sd 467) * $signed(input_fmap_105[15:0]) +
	( 16'sd 26030) * $signed(input_fmap_106[15:0]) +
	( 16'sd 29363) * $signed(input_fmap_107[15:0]) +
	( 15'sd 11806) * $signed(input_fmap_108[15:0]) +
	( 16'sd 31564) * $signed(input_fmap_109[15:0]) +
	( 15'sd 13442) * $signed(input_fmap_110[15:0]) +
	( 15'sd 15117) * $signed(input_fmap_111[15:0]) +
	( 12'sd 1670) * $signed(input_fmap_112[15:0]) +
	( 10'sd 318) * $signed(input_fmap_113[15:0]) +
	( 8'sd 110) * $signed(input_fmap_114[15:0]) +
	( 16'sd 30254) * $signed(input_fmap_115[15:0]) +
	( 13'sd 3395) * $signed(input_fmap_116[15:0]) +
	( 16'sd 19200) * $signed(input_fmap_117[15:0]) +
	( 15'sd 13719) * $signed(input_fmap_118[15:0]) +
	( 16'sd 19396) * $signed(input_fmap_119[15:0]) +
	( 12'sd 1611) * $signed(input_fmap_120[15:0]) +
	( 16'sd 19246) * $signed(input_fmap_121[15:0]) +
	( 15'sd 14546) * $signed(input_fmap_122[15:0]) +
	( 13'sd 2206) * $signed(input_fmap_123[15:0]) +
	( 16'sd 19509) * $signed(input_fmap_124[15:0]) +
	( 16'sd 20710) * $signed(input_fmap_125[15:0]) +
	( 16'sd 24589) * $signed(input_fmap_126[15:0]) +
	( 16'sd 18237) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 16'sd 25786) * $signed(input_fmap_0[15:0]) +
	( 16'sd 25490) * $signed(input_fmap_1[15:0]) +
	( 16'sd 25078) * $signed(input_fmap_2[15:0]) +
	( 16'sd 23535) * $signed(input_fmap_3[15:0]) +
	( 14'sd 4732) * $signed(input_fmap_4[15:0]) +
	( 16'sd 29867) * $signed(input_fmap_5[15:0]) +
	( 16'sd 16680) * $signed(input_fmap_6[15:0]) +
	( 15'sd 12326) * $signed(input_fmap_7[15:0]) +
	( 15'sd 8365) * $signed(input_fmap_8[15:0]) +
	( 15'sd 15166) * $signed(input_fmap_9[15:0]) +
	( 15'sd 14910) * $signed(input_fmap_10[15:0]) +
	( 14'sd 6013) * $signed(input_fmap_11[15:0]) +
	( 14'sd 8105) * $signed(input_fmap_12[15:0]) +
	( 16'sd 21541) * $signed(input_fmap_13[15:0]) +
	( 15'sd 9541) * $signed(input_fmap_14[15:0]) +
	( 15'sd 14983) * $signed(input_fmap_15[15:0]) +
	( 16'sd 30362) * $signed(input_fmap_16[15:0]) +
	( 14'sd 4337) * $signed(input_fmap_17[15:0]) +
	( 16'sd 17418) * $signed(input_fmap_18[15:0]) +
	( 16'sd 23807) * $signed(input_fmap_19[15:0]) +
	( 16'sd 29631) * $signed(input_fmap_20[15:0]) +
	( 16'sd 30407) * $signed(input_fmap_21[15:0]) +
	( 14'sd 8137) * $signed(input_fmap_22[15:0]) +
	( 15'sd 15859) * $signed(input_fmap_23[15:0]) +
	( 15'sd 12954) * $signed(input_fmap_24[15:0]) +
	( 13'sd 3954) * $signed(input_fmap_25[15:0]) +
	( 14'sd 4975) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1539) * $signed(input_fmap_27[15:0]) +
	( 16'sd 21292) * $signed(input_fmap_28[15:0]) +
	( 13'sd 3833) * $signed(input_fmap_29[15:0]) +
	( 14'sd 7089) * $signed(input_fmap_30[15:0]) +
	( 15'sd 12133) * $signed(input_fmap_31[15:0]) +
	( 16'sd 24770) * $signed(input_fmap_32[15:0]) +
	( 16'sd 17745) * $signed(input_fmap_33[15:0]) +
	( 16'sd 29022) * $signed(input_fmap_34[15:0]) +
	( 16'sd 21014) * $signed(input_fmap_35[15:0]) +
	( 15'sd 15399) * $signed(input_fmap_36[15:0]) +
	( 14'sd 6307) * $signed(input_fmap_37[15:0]) +
	( 16'sd 30127) * $signed(input_fmap_38[15:0]) +
	( 16'sd 25744) * $signed(input_fmap_39[15:0]) +
	( 16'sd 30257) * $signed(input_fmap_40[15:0]) +
	( 16'sd 22047) * $signed(input_fmap_41[15:0]) +
	( 16'sd 25221) * $signed(input_fmap_42[15:0]) +
	( 15'sd 14567) * $signed(input_fmap_43[15:0]) +
	( 16'sd 18479) * $signed(input_fmap_44[15:0]) +
	( 15'sd 12219) * $signed(input_fmap_45[15:0]) +
	( 15'sd 8291) * $signed(input_fmap_46[15:0]) +
	( 16'sd 23861) * $signed(input_fmap_47[15:0]) +
	( 15'sd 9810) * $signed(input_fmap_48[15:0]) +
	( 16'sd 23514) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26051) * $signed(input_fmap_50[15:0]) +
	( 16'sd 31070) * $signed(input_fmap_51[15:0]) +
	( 14'sd 7532) * $signed(input_fmap_52[15:0]) +
	( 14'sd 5756) * $signed(input_fmap_53[15:0]) +
	( 16'sd 22718) * $signed(input_fmap_54[15:0]) +
	( 13'sd 2067) * $signed(input_fmap_55[15:0]) +
	( 16'sd 27770) * $signed(input_fmap_56[15:0]) +
	( 16'sd 30017) * $signed(input_fmap_57[15:0]) +
	( 11'sd 773) * $signed(input_fmap_58[15:0]) +
	( 16'sd 18446) * $signed(input_fmap_59[15:0]) +
	( 16'sd 19662) * $signed(input_fmap_60[15:0]) +
	( 12'sd 1455) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29544) * $signed(input_fmap_62[15:0]) +
	( 15'sd 9118) * $signed(input_fmap_63[15:0]) +
	( 16'sd 21733) * $signed(input_fmap_64[15:0]) +
	( 15'sd 15237) * $signed(input_fmap_65[15:0]) +
	( 12'sd 1808) * $signed(input_fmap_66[15:0]) +
	( 16'sd 17814) * $signed(input_fmap_67[15:0]) +
	( 16'sd 20625) * $signed(input_fmap_68[15:0]) +
	( 10'sd 281) * $signed(input_fmap_69[15:0]) +
	( 16'sd 20982) * $signed(input_fmap_70[15:0]) +
	( 15'sd 15558) * $signed(input_fmap_71[15:0]) +
	( 16'sd 32343) * $signed(input_fmap_72[15:0]) +
	( 14'sd 5105) * $signed(input_fmap_73[15:0]) +
	( 16'sd 30073) * $signed(input_fmap_74[15:0]) +
	( 15'sd 13863) * $signed(input_fmap_75[15:0]) +
	( 16'sd 18002) * $signed(input_fmap_76[15:0]) +
	( 13'sd 3877) * $signed(input_fmap_77[15:0]) +
	( 13'sd 3221) * $signed(input_fmap_78[15:0]) +
	( 15'sd 13944) * $signed(input_fmap_79[15:0]) +
	( 16'sd 30679) * $signed(input_fmap_80[15:0]) +
	( 16'sd 17007) * $signed(input_fmap_81[15:0]) +
	( 9'sd 207) * $signed(input_fmap_82[15:0]) +
	( 16'sd 22832) * $signed(input_fmap_83[15:0]) +
	( 16'sd 29686) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24726) * $signed(input_fmap_85[15:0]) +
	( 16'sd 29421) * $signed(input_fmap_86[15:0]) +
	( 14'sd 4171) * $signed(input_fmap_87[15:0]) +
	( 15'sd 8648) * $signed(input_fmap_88[15:0]) +
	( 13'sd 4035) * $signed(input_fmap_89[15:0]) +
	( 15'sd 12602) * $signed(input_fmap_90[15:0]) +
	( 16'sd 18075) * $signed(input_fmap_91[15:0]) +
	( 12'sd 1865) * $signed(input_fmap_92[15:0]) +
	( 16'sd 16461) * $signed(input_fmap_93[15:0]) +
	( 16'sd 31463) * $signed(input_fmap_94[15:0]) +
	( 15'sd 15241) * $signed(input_fmap_95[15:0]) +
	( 15'sd 11807) * $signed(input_fmap_96[15:0]) +
	( 15'sd 13232) * $signed(input_fmap_97[15:0]) +
	( 15'sd 15379) * $signed(input_fmap_98[15:0]) +
	( 16'sd 26315) * $signed(input_fmap_99[15:0]) +
	( 15'sd 8952) * $signed(input_fmap_100[15:0]) +
	( 10'sd 272) * $signed(input_fmap_101[15:0]) +
	( 14'sd 7628) * $signed(input_fmap_102[15:0]) +
	( 16'sd 27933) * $signed(input_fmap_103[15:0]) +
	( 16'sd 30836) * $signed(input_fmap_104[15:0]) +
	( 16'sd 22307) * $signed(input_fmap_105[15:0]) +
	( 16'sd 21231) * $signed(input_fmap_106[15:0]) +
	( 16'sd 30822) * $signed(input_fmap_107[15:0]) +
	( 15'sd 16225) * $signed(input_fmap_108[15:0]) +
	( 15'sd 13384) * $signed(input_fmap_109[15:0]) +
	( 14'sd 7567) * $signed(input_fmap_110[15:0]) +
	( 15'sd 16278) * $signed(input_fmap_111[15:0]) +
	( 16'sd 19288) * $signed(input_fmap_112[15:0]) +
	( 14'sd 6443) * $signed(input_fmap_113[15:0]) +
	( 12'sd 1517) * $signed(input_fmap_114[15:0]) +
	( 15'sd 14781) * $signed(input_fmap_115[15:0]) +
	( 16'sd 16692) * $signed(input_fmap_116[15:0]) +
	( 16'sd 28502) * $signed(input_fmap_117[15:0]) +
	( 16'sd 26976) * $signed(input_fmap_118[15:0]) +
	( 16'sd 17335) * $signed(input_fmap_119[15:0]) +
	( 15'sd 11936) * $signed(input_fmap_120[15:0]) +
	( 13'sd 3837) * $signed(input_fmap_121[15:0]) +
	( 15'sd 15000) * $signed(input_fmap_122[15:0]) +
	( 14'sd 5704) * $signed(input_fmap_123[15:0]) +
	( 15'sd 9375) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24141) * $signed(input_fmap_125[15:0]) +
	( 14'sd 4331) * $signed(input_fmap_126[15:0]) +
	( 15'sd 10124) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 14'sd 4192) * $signed(input_fmap_0[15:0]) +
	( 16'sd 29303) * $signed(input_fmap_1[15:0]) +
	( 16'sd 17082) * $signed(input_fmap_2[15:0]) +
	( 13'sd 3829) * $signed(input_fmap_3[15:0]) +
	( 16'sd 29188) * $signed(input_fmap_4[15:0]) +
	( 13'sd 2617) * $signed(input_fmap_5[15:0]) +
	( 16'sd 25914) * $signed(input_fmap_6[15:0]) +
	( 16'sd 31896) * $signed(input_fmap_7[15:0]) +
	( 16'sd 27513) * $signed(input_fmap_8[15:0]) +
	( 14'sd 4639) * $signed(input_fmap_9[15:0]) +
	( 15'sd 10207) * $signed(input_fmap_10[15:0]) +
	( 16'sd 24060) * $signed(input_fmap_11[15:0]) +
	( 16'sd 27404) * $signed(input_fmap_12[15:0]) +
	( 16'sd 25532) * $signed(input_fmap_13[15:0]) +
	( 16'sd 17684) * $signed(input_fmap_14[15:0]) +
	( 16'sd 16772) * $signed(input_fmap_15[15:0]) +
	( 15'sd 9261) * $signed(input_fmap_16[15:0]) +
	( 15'sd 11866) * $signed(input_fmap_17[15:0]) +
	( 16'sd 24063) * $signed(input_fmap_18[15:0]) +
	( 14'sd 5543) * $signed(input_fmap_19[15:0]) +
	( 15'sd 10393) * $signed(input_fmap_20[15:0]) +
	( 16'sd 19999) * $signed(input_fmap_21[15:0]) +
	( 15'sd 14300) * $signed(input_fmap_22[15:0]) +
	( 13'sd 3810) * $signed(input_fmap_23[15:0]) +
	( 16'sd 29866) * $signed(input_fmap_24[15:0]) +
	( 16'sd 27840) * $signed(input_fmap_25[15:0]) +
	( 16'sd 28025) * $signed(input_fmap_26[15:0]) +
	( 16'sd 22649) * $signed(input_fmap_27[15:0]) +
	( 14'sd 8178) * $signed(input_fmap_28[15:0]) +
	( 16'sd 25948) * $signed(input_fmap_29[15:0]) +
	( 14'sd 4990) * $signed(input_fmap_30[15:0]) +
	( 16'sd 31111) * $signed(input_fmap_31[15:0]) +
	( 12'sd 1852) * $signed(input_fmap_32[15:0]) +
	( 14'sd 4181) * $signed(input_fmap_33[15:0]) +
	( 16'sd 31849) * $signed(input_fmap_34[15:0]) +
	( 16'sd 17671) * $signed(input_fmap_35[15:0]) +
	( 14'sd 7271) * $signed(input_fmap_36[15:0]) +
	( 16'sd 23410) * $signed(input_fmap_37[15:0]) +
	( 14'sd 5395) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24635) * $signed(input_fmap_39[15:0]) +
	( 16'sd 27595) * $signed(input_fmap_40[15:0]) +
	( 16'sd 19713) * $signed(input_fmap_41[15:0]) +
	( 16'sd 24681) * $signed(input_fmap_42[15:0]) +
	( 16'sd 29113) * $signed(input_fmap_43[15:0]) +
	( 15'sd 8929) * $signed(input_fmap_44[15:0]) +
	( 14'sd 6796) * $signed(input_fmap_45[15:0]) +
	( 15'sd 12018) * $signed(input_fmap_46[15:0]) +
	( 16'sd 19344) * $signed(input_fmap_47[15:0]) +
	( 15'sd 9538) * $signed(input_fmap_48[15:0]) +
	( 15'sd 9719) * $signed(input_fmap_49[15:0]) +
	( 16'sd 18318) * $signed(input_fmap_50[15:0]) +
	( 14'sd 6787) * $signed(input_fmap_51[15:0]) +
	( 15'sd 16341) * $signed(input_fmap_52[15:0]) +
	( 16'sd 23871) * $signed(input_fmap_53[15:0]) +
	( 15'sd 12823) * $signed(input_fmap_54[15:0]) +
	( 15'sd 15396) * $signed(input_fmap_55[15:0]) +
	( 16'sd 27989) * $signed(input_fmap_56[15:0]) +
	( 16'sd 26503) * $signed(input_fmap_57[15:0]) +
	( 16'sd 25841) * $signed(input_fmap_58[15:0]) +
	( 16'sd 27860) * $signed(input_fmap_59[15:0]) +
	( 13'sd 2248) * $signed(input_fmap_60[15:0]) +
	( 15'sd 9491) * $signed(input_fmap_61[15:0]) +
	( 14'sd 5342) * $signed(input_fmap_62[15:0]) +
	( 13'sd 2226) * $signed(input_fmap_63[15:0]) +
	( 15'sd 13812) * $signed(input_fmap_64[15:0]) +
	( 15'sd 14177) * $signed(input_fmap_65[15:0]) +
	( 16'sd 17916) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28020) * $signed(input_fmap_67[15:0]) +
	( 15'sd 10547) * $signed(input_fmap_68[15:0]) +
	( 13'sd 4093) * $signed(input_fmap_69[15:0]) +
	( 16'sd 25178) * $signed(input_fmap_70[15:0]) +
	( 16'sd 29060) * $signed(input_fmap_71[15:0]) +
	( 16'sd 23739) * $signed(input_fmap_72[15:0]) +
	( 13'sd 2247) * $signed(input_fmap_73[15:0]) +
	( 16'sd 27907) * $signed(input_fmap_74[15:0]) +
	( 16'sd 26279) * $signed(input_fmap_75[15:0]) +
	( 16'sd 28554) * $signed(input_fmap_76[15:0]) +
	( 16'sd 27309) * $signed(input_fmap_77[15:0]) +
	( 9'sd 238) * $signed(input_fmap_78[15:0]) +
	( 15'sd 13926) * $signed(input_fmap_79[15:0]) +
	( 16'sd 30847) * $signed(input_fmap_80[15:0]) +
	( 15'sd 16122) * $signed(input_fmap_81[15:0]) +
	( 16'sd 27465) * $signed(input_fmap_82[15:0]) +
	( 15'sd 9282) * $signed(input_fmap_83[15:0]) +
	( 16'sd 29878) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24175) * $signed(input_fmap_85[15:0]) +
	( 16'sd 23943) * $signed(input_fmap_86[15:0]) +
	( 16'sd 20246) * $signed(input_fmap_87[15:0]) +
	( 16'sd 22320) * $signed(input_fmap_88[15:0]) +
	( 16'sd 31565) * $signed(input_fmap_89[15:0]) +
	( 15'sd 14045) * $signed(input_fmap_90[15:0]) +
	( 15'sd 9569) * $signed(input_fmap_91[15:0]) +
	( 15'sd 14565) * $signed(input_fmap_92[15:0]) +
	( 16'sd 21413) * $signed(input_fmap_93[15:0]) +
	( 14'sd 5104) * $signed(input_fmap_94[15:0]) +
	( 15'sd 10604) * $signed(input_fmap_95[15:0]) +
	( 14'sd 8188) * $signed(input_fmap_96[15:0]) +
	( 13'sd 2438) * $signed(input_fmap_97[15:0]) +
	( 16'sd 32281) * $signed(input_fmap_98[15:0]) +
	( 14'sd 4255) * $signed(input_fmap_99[15:0]) +
	( 15'sd 15934) * $signed(input_fmap_100[15:0]) +
	( 15'sd 16228) * $signed(input_fmap_101[15:0]) +
	( 14'sd 7271) * $signed(input_fmap_102[15:0]) +
	( 14'sd 7777) * $signed(input_fmap_103[15:0]) +
	( 16'sd 31825) * $signed(input_fmap_104[15:0]) +
	( 10'sd 267) * $signed(input_fmap_105[15:0]) +
	( 16'sd 32544) * $signed(input_fmap_106[15:0]) +
	( 16'sd 26518) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15536) * $signed(input_fmap_108[15:0]) +
	( 16'sd 26752) * $signed(input_fmap_109[15:0]) +
	( 16'sd 16695) * $signed(input_fmap_110[15:0]) +
	( 16'sd 32516) * $signed(input_fmap_111[15:0]) +
	( 14'sd 6647) * $signed(input_fmap_112[15:0]) +
	( 16'sd 19730) * $signed(input_fmap_113[15:0]) +
	( 15'sd 8224) * $signed(input_fmap_114[15:0]) +
	( 16'sd 25253) * $signed(input_fmap_115[15:0]) +
	( 16'sd 21150) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27200) * $signed(input_fmap_117[15:0]) +
	( 16'sd 16885) * $signed(input_fmap_118[15:0]) +
	( 16'sd 17833) * $signed(input_fmap_119[15:0]) +
	( 15'sd 8371) * $signed(input_fmap_120[15:0]) +
	( 15'sd 14660) * $signed(input_fmap_121[15:0]) +
	( 16'sd 17050) * $signed(input_fmap_122[15:0]) +
	( 16'sd 27367) * $signed(input_fmap_123[15:0]) +
	( 16'sd 25646) * $signed(input_fmap_124[15:0]) +
	( 14'sd 7120) * $signed(input_fmap_125[15:0]) +
	( 16'sd 24466) * $signed(input_fmap_126[15:0]) +
	( 16'sd 28597) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 16'sd 17100) * $signed(input_fmap_0[15:0]) +
	( 16'sd 16491) * $signed(input_fmap_1[15:0]) +
	( 16'sd 25896) * $signed(input_fmap_2[15:0]) +
	( 16'sd 18894) * $signed(input_fmap_3[15:0]) +
	( 16'sd 25868) * $signed(input_fmap_4[15:0]) +
	( 15'sd 8816) * $signed(input_fmap_5[15:0]) +
	( 16'sd 26020) * $signed(input_fmap_6[15:0]) +
	( 16'sd 27977) * $signed(input_fmap_7[15:0]) +
	( 15'sd 12065) * $signed(input_fmap_8[15:0]) +
	( 12'sd 1869) * $signed(input_fmap_9[15:0]) +
	( 15'sd 12902) * $signed(input_fmap_10[15:0]) +
	( 16'sd 20397) * $signed(input_fmap_11[15:0]) +
	( 13'sd 3513) * $signed(input_fmap_12[15:0]) +
	( 16'sd 27676) * $signed(input_fmap_13[15:0]) +
	( 15'sd 13086) * $signed(input_fmap_14[15:0]) +
	( 15'sd 12112) * $signed(input_fmap_15[15:0]) +
	( 13'sd 2413) * $signed(input_fmap_16[15:0]) +
	( 15'sd 9462) * $signed(input_fmap_17[15:0]) +
	( 16'sd 26309) * $signed(input_fmap_18[15:0]) +
	( 14'sd 5298) * $signed(input_fmap_19[15:0]) +
	( 16'sd 27148) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17868) * $signed(input_fmap_21[15:0]) +
	( 15'sd 14612) * $signed(input_fmap_22[15:0]) +
	( 16'sd 18396) * $signed(input_fmap_23[15:0]) +
	( 16'sd 24309) * $signed(input_fmap_24[15:0]) +
	( 12'sd 1661) * $signed(input_fmap_25[15:0]) +
	( 14'sd 4834) * $signed(input_fmap_26[15:0]) +
	( 15'sd 11706) * $signed(input_fmap_27[15:0]) +
	( 14'sd 6639) * $signed(input_fmap_28[15:0]) +
	( 15'sd 13766) * $signed(input_fmap_29[15:0]) +
	( 15'sd 10678) * $signed(input_fmap_30[15:0]) +
	( 8'sd 88) * $signed(input_fmap_31[15:0]) +
	( 14'sd 5740) * $signed(input_fmap_32[15:0]) +
	( 16'sd 27945) * $signed(input_fmap_33[15:0]) +
	( 16'sd 16753) * $signed(input_fmap_34[15:0]) +
	( 13'sd 3377) * $signed(input_fmap_35[15:0]) +
	( 15'sd 8289) * $signed(input_fmap_36[15:0]) +
	( 16'sd 31933) * $signed(input_fmap_37[15:0]) +
	( 14'sd 6426) * $signed(input_fmap_38[15:0]) +
	( 16'sd 22545) * $signed(input_fmap_39[15:0]) +
	( 16'sd 25693) * $signed(input_fmap_40[15:0]) +
	( 16'sd 19418) * $signed(input_fmap_41[15:0]) +
	( 15'sd 15738) * $signed(input_fmap_42[15:0]) +
	( 15'sd 14285) * $signed(input_fmap_43[15:0]) +
	( 16'sd 16946) * $signed(input_fmap_44[15:0]) +
	( 16'sd 18149) * $signed(input_fmap_45[15:0]) +
	( 11'sd 537) * $signed(input_fmap_46[15:0]) +
	( 15'sd 10308) * $signed(input_fmap_47[15:0]) +
	( 13'sd 3935) * $signed(input_fmap_48[15:0]) +
	( 15'sd 16223) * $signed(input_fmap_49[15:0]) +
	( 15'sd 14890) * $signed(input_fmap_50[15:0]) +
	( 16'sd 27213) * $signed(input_fmap_51[15:0]) +
	( 14'sd 7710) * $signed(input_fmap_52[15:0]) +
	( 16'sd 28926) * $signed(input_fmap_53[15:0]) +
	( 13'sd 2787) * $signed(input_fmap_54[15:0]) +
	( 16'sd 25279) * $signed(input_fmap_55[15:0]) +
	( 16'sd 18756) * $signed(input_fmap_56[15:0]) +
	( 16'sd 20405) * $signed(input_fmap_57[15:0]) +
	( 16'sd 32112) * $signed(input_fmap_58[15:0]) +
	( 12'sd 1575) * $signed(input_fmap_59[15:0]) +
	( 15'sd 14271) * $signed(input_fmap_60[15:0]) +
	( 12'sd 1739) * $signed(input_fmap_61[15:0]) +
	( 14'sd 7149) * $signed(input_fmap_62[15:0]) +
	( 16'sd 27939) * $signed(input_fmap_63[15:0]) +
	( 16'sd 32459) * $signed(input_fmap_64[15:0]) +
	( 16'sd 31716) * $signed(input_fmap_65[15:0]) +
	( 16'sd 26945) * $signed(input_fmap_66[15:0]) +
	( 16'sd 25215) * $signed(input_fmap_67[15:0]) +
	( 16'sd 30952) * $signed(input_fmap_68[15:0]) +
	( 16'sd 16742) * $signed(input_fmap_69[15:0]) +
	( 15'sd 8531) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11921) * $signed(input_fmap_71[15:0]) +
	( 14'sd 4612) * $signed(input_fmap_72[15:0]) +
	( 16'sd 21129) * $signed(input_fmap_73[15:0]) +
	( 14'sd 7094) * $signed(input_fmap_74[15:0]) +
	( 15'sd 8823) * $signed(input_fmap_75[15:0]) +
	( 16'sd 29053) * $signed(input_fmap_76[15:0]) +
	( 16'sd 32254) * $signed(input_fmap_77[15:0]) +
	( 16'sd 25864) * $signed(input_fmap_78[15:0]) +
	( 16'sd 32368) * $signed(input_fmap_79[15:0]) +
	( 13'sd 3299) * $signed(input_fmap_80[15:0]) +
	( 16'sd 20313) * $signed(input_fmap_81[15:0]) +
	( 16'sd 23482) * $signed(input_fmap_82[15:0]) +
	( 15'sd 8563) * $signed(input_fmap_83[15:0]) +
	( 15'sd 14400) * $signed(input_fmap_84[15:0]) +
	( 16'sd 28482) * $signed(input_fmap_85[15:0]) +
	( 12'sd 1076) * $signed(input_fmap_86[15:0]) +
	( 16'sd 26329) * $signed(input_fmap_87[15:0]) +
	( 15'sd 11249) * $signed(input_fmap_88[15:0]) +
	( 15'sd 14076) * $signed(input_fmap_89[15:0]) +
	( 16'sd 20940) * $signed(input_fmap_90[15:0]) +
	( 15'sd 9030) * $signed(input_fmap_91[15:0]) +
	( 14'sd 7734) * $signed(input_fmap_92[15:0]) +
	( 12'sd 1258) * $signed(input_fmap_93[15:0]) +
	( 16'sd 17716) * $signed(input_fmap_94[15:0]) +
	( 15'sd 14009) * $signed(input_fmap_95[15:0]) +
	( 12'sd 1463) * $signed(input_fmap_96[15:0]) +
	( 16'sd 18820) * $signed(input_fmap_97[15:0]) +
	( 14'sd 4289) * $signed(input_fmap_98[15:0]) +
	( 16'sd 17410) * $signed(input_fmap_99[15:0]) +
	( 16'sd 24891) * $signed(input_fmap_100[15:0]) +
	( 16'sd 24532) * $signed(input_fmap_101[15:0]) +
	( 16'sd 20071) * $signed(input_fmap_102[15:0]) +
	( 15'sd 9450) * $signed(input_fmap_103[15:0]) +
	( 16'sd 17819) * $signed(input_fmap_104[15:0]) +
	( 16'sd 30008) * $signed(input_fmap_105[15:0]) +
	( 16'sd 20042) * $signed(input_fmap_106[15:0]) +
	( 15'sd 10313) * $signed(input_fmap_107[15:0]) +
	( 16'sd 18589) * $signed(input_fmap_108[15:0]) +
	( 16'sd 18680) * $signed(input_fmap_109[15:0]) +
	( 16'sd 25026) * $signed(input_fmap_110[15:0]) +
	( 16'sd 31258) * $signed(input_fmap_111[15:0]) +
	( 14'sd 5200) * $signed(input_fmap_112[15:0]) +
	( 16'sd 19458) * $signed(input_fmap_113[15:0]) +
	( 16'sd 21872) * $signed(input_fmap_114[15:0]) +
	( 16'sd 27213) * $signed(input_fmap_115[15:0]) +
	( 15'sd 10924) * $signed(input_fmap_116[15:0]) +
	( 15'sd 14650) * $signed(input_fmap_117[15:0]) +
	( 14'sd 6808) * $signed(input_fmap_118[15:0]) +
	( 14'sd 4478) * $signed(input_fmap_119[15:0]) +
	( 16'sd 23248) * $signed(input_fmap_120[15:0]) +
	( 16'sd 18458) * $signed(input_fmap_121[15:0]) +
	( 15'sd 11211) * $signed(input_fmap_122[15:0]) +
	( 15'sd 11666) * $signed(input_fmap_123[15:0]) +
	( 15'sd 12145) * $signed(input_fmap_124[15:0]) +
	( 16'sd 32213) * $signed(input_fmap_125[15:0]) +
	( 12'sd 1357) * $signed(input_fmap_126[15:0]) +
	( 11'sd 785) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 16'sd 22721) * $signed(input_fmap_0[15:0]) +
	( 16'sd 21769) * $signed(input_fmap_1[15:0]) +
	( 14'sd 5562) * $signed(input_fmap_2[15:0]) +
	( 15'sd 15774) * $signed(input_fmap_3[15:0]) +
	( 15'sd 14945) * $signed(input_fmap_4[15:0]) +
	( 15'sd 14503) * $signed(input_fmap_5[15:0]) +
	( 16'sd 28133) * $signed(input_fmap_6[15:0]) +
	( 12'sd 1378) * $signed(input_fmap_7[15:0]) +
	( 15'sd 12153) * $signed(input_fmap_8[15:0]) +
	( 13'sd 2944) * $signed(input_fmap_9[15:0]) +
	( 13'sd 3980) * $signed(input_fmap_10[15:0]) +
	( 16'sd 19980) * $signed(input_fmap_11[15:0]) +
	( 16'sd 26654) * $signed(input_fmap_12[15:0]) +
	( 13'sd 2768) * $signed(input_fmap_13[15:0]) +
	( 16'sd 27130) * $signed(input_fmap_14[15:0]) +
	( 16'sd 23710) * $signed(input_fmap_15[15:0]) +
	( 15'sd 14272) * $signed(input_fmap_16[15:0]) +
	( 14'sd 6725) * $signed(input_fmap_17[15:0]) +
	( 15'sd 15192) * $signed(input_fmap_18[15:0]) +
	( 15'sd 10481) * $signed(input_fmap_19[15:0]) +
	( 16'sd 17566) * $signed(input_fmap_20[15:0]) +
	( 15'sd 13408) * $signed(input_fmap_21[15:0]) +
	( 15'sd 12838) * $signed(input_fmap_22[15:0]) +
	( 16'sd 27576) * $signed(input_fmap_23[15:0]) +
	( 16'sd 31952) * $signed(input_fmap_24[15:0]) +
	( 15'sd 8934) * $signed(input_fmap_25[15:0]) +
	( 16'sd 24608) * $signed(input_fmap_26[15:0]) +
	( 16'sd 18061) * $signed(input_fmap_27[15:0]) +
	( 14'sd 5214) * $signed(input_fmap_28[15:0]) +
	( 11'sd 783) * $signed(input_fmap_29[15:0]) +
	( 14'sd 6742) * $signed(input_fmap_30[15:0]) +
	( 15'sd 15058) * $signed(input_fmap_31[15:0]) +
	( 16'sd 25703) * $signed(input_fmap_32[15:0]) +
	( 15'sd 10478) * $signed(input_fmap_33[15:0]) +
	( 15'sd 8351) * $signed(input_fmap_34[15:0]) +
	( 15'sd 9450) * $signed(input_fmap_35[15:0]) +
	( 16'sd 19324) * $signed(input_fmap_36[15:0]) +
	( 14'sd 5494) * $signed(input_fmap_37[15:0]) +
	( 16'sd 21214) * $signed(input_fmap_38[15:0]) +
	( 15'sd 8469) * $signed(input_fmap_39[15:0]) +
	( 15'sd 12432) * $signed(input_fmap_40[15:0]) +
	( 15'sd 14590) * $signed(input_fmap_41[15:0]) +
	( 15'sd 15610) * $signed(input_fmap_42[15:0]) +
	( 16'sd 25345) * $signed(input_fmap_43[15:0]) +
	( 15'sd 9059) * $signed(input_fmap_44[15:0]) +
	( 15'sd 13362) * $signed(input_fmap_45[15:0]) +
	( 16'sd 25086) * $signed(input_fmap_46[15:0]) +
	( 15'sd 10254) * $signed(input_fmap_47[15:0]) +
	( 15'sd 12225) * $signed(input_fmap_48[15:0]) +
	( 14'sd 6344) * $signed(input_fmap_49[15:0]) +
	( 13'sd 2106) * $signed(input_fmap_50[15:0]) +
	( 16'sd 32238) * $signed(input_fmap_51[15:0]) +
	( 14'sd 5693) * $signed(input_fmap_52[15:0]) +
	( 11'sd 905) * $signed(input_fmap_53[15:0]) +
	( 14'sd 6363) * $signed(input_fmap_54[15:0]) +
	( 14'sd 6302) * $signed(input_fmap_55[15:0]) +
	( 16'sd 18015) * $signed(input_fmap_56[15:0]) +
	( 16'sd 21942) * $signed(input_fmap_57[15:0]) +
	( 16'sd 18193) * $signed(input_fmap_58[15:0]) +
	( 16'sd 31619) * $signed(input_fmap_59[15:0]) +
	( 16'sd 23313) * $signed(input_fmap_60[15:0]) +
	( 15'sd 11856) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29216) * $signed(input_fmap_62[15:0]) +
	( 15'sd 11986) * $signed(input_fmap_63[15:0]) +
	( 14'sd 5054) * $signed(input_fmap_64[15:0]) +
	( 16'sd 23054) * $signed(input_fmap_65[15:0]) +
	( 16'sd 17887) * $signed(input_fmap_66[15:0]) +
	( 16'sd 23618) * $signed(input_fmap_67[15:0]) +
	( 16'sd 29744) * $signed(input_fmap_68[15:0]) +
	( 14'sd 7046) * $signed(input_fmap_69[15:0]) +
	( 15'sd 15874) * $signed(input_fmap_70[15:0]) +
	( 15'sd 12472) * $signed(input_fmap_71[15:0]) +
	( 16'sd 31506) * $signed(input_fmap_72[15:0]) +
	( 16'sd 28130) * $signed(input_fmap_73[15:0]) +
	( 16'sd 19582) * $signed(input_fmap_74[15:0]) +
	( 16'sd 19731) * $signed(input_fmap_75[15:0]) +
	( 16'sd 23284) * $signed(input_fmap_76[15:0]) +
	( 16'sd 22131) * $signed(input_fmap_77[15:0]) +
	( 15'sd 10772) * $signed(input_fmap_78[15:0]) +
	( 14'sd 6436) * $signed(input_fmap_79[15:0]) +
	( 13'sd 2373) * $signed(input_fmap_80[15:0]) +
	( 12'sd 1323) * $signed(input_fmap_81[15:0]) +
	( 15'sd 8488) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25951) * $signed(input_fmap_83[15:0]) +
	( 15'sd 13921) * $signed(input_fmap_84[15:0]) +
	( 16'sd 32095) * $signed(input_fmap_85[15:0]) +
	( 16'sd 18827) * $signed(input_fmap_86[15:0]) +
	( 15'sd 8607) * $signed(input_fmap_87[15:0]) +
	( 15'sd 12538) * $signed(input_fmap_88[15:0]) +
	( 16'sd 26985) * $signed(input_fmap_89[15:0]) +
	( 15'sd 8706) * $signed(input_fmap_90[15:0]) +
	( 15'sd 14773) * $signed(input_fmap_91[15:0]) +
	( 15'sd 11524) * $signed(input_fmap_92[15:0]) +
	( 16'sd 23902) * $signed(input_fmap_93[15:0]) +
	( 8'sd 127) * $signed(input_fmap_94[15:0]) +
	( 16'sd 23710) * $signed(input_fmap_95[15:0]) +
	( 15'sd 11145) * $signed(input_fmap_96[15:0]) +
	( 16'sd 31969) * $signed(input_fmap_97[15:0]) +
	( 16'sd 29625) * $signed(input_fmap_98[15:0]) +
	( 15'sd 14161) * $signed(input_fmap_99[15:0]) +
	( 15'sd 16259) * $signed(input_fmap_100[15:0]) +
	( 15'sd 8494) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5475) * $signed(input_fmap_102[15:0]) +
	( 14'sd 6083) * $signed(input_fmap_103[15:0]) +
	( 15'sd 9484) * $signed(input_fmap_104[15:0]) +
	( 16'sd 19020) * $signed(input_fmap_105[15:0]) +
	( 14'sd 6910) * $signed(input_fmap_106[15:0]) +
	( 14'sd 5700) * $signed(input_fmap_107[15:0]) +
	( 15'sd 8837) * $signed(input_fmap_108[15:0]) +
	( 16'sd 29049) * $signed(input_fmap_109[15:0]) +
	( 16'sd 20740) * $signed(input_fmap_110[15:0]) +
	( 16'sd 18736) * $signed(input_fmap_111[15:0]) +
	( 16'sd 29665) * $signed(input_fmap_112[15:0]) +
	( 16'sd 16547) * $signed(input_fmap_113[15:0]) +
	( 16'sd 32117) * $signed(input_fmap_114[15:0]) +
	( 16'sd 16650) * $signed(input_fmap_115[15:0]) +
	( 15'sd 16202) * $signed(input_fmap_116[15:0]) +
	( 13'sd 2719) * $signed(input_fmap_117[15:0]) +
	( 15'sd 13592) * $signed(input_fmap_118[15:0]) +
	( 15'sd 8951) * $signed(input_fmap_119[15:0]) +
	( 15'sd 10457) * $signed(input_fmap_120[15:0]) +
	( 14'sd 6005) * $signed(input_fmap_121[15:0]) +
	( 16'sd 29037) * $signed(input_fmap_122[15:0]) +
	( 11'sd 669) * $signed(input_fmap_123[15:0]) +
	( 16'sd 27177) * $signed(input_fmap_124[15:0]) +
	( 13'sd 3134) * $signed(input_fmap_125[15:0]) +
	( 15'sd 8965) * $signed(input_fmap_126[15:0]) +
	( 16'sd 24683) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 16'sd 29210) * $signed(input_fmap_0[15:0]) +
	( 16'sd 25786) * $signed(input_fmap_1[15:0]) +
	( 16'sd 25972) * $signed(input_fmap_2[15:0]) +
	( 16'sd 32253) * $signed(input_fmap_3[15:0]) +
	( 16'sd 31793) * $signed(input_fmap_4[15:0]) +
	( 16'sd 27802) * $signed(input_fmap_5[15:0]) +
	( 14'sd 7148) * $signed(input_fmap_6[15:0]) +
	( 15'sd 9166) * $signed(input_fmap_7[15:0]) +
	( 15'sd 14193) * $signed(input_fmap_8[15:0]) +
	( 16'sd 30290) * $signed(input_fmap_9[15:0]) +
	( 16'sd 24847) * $signed(input_fmap_10[15:0]) +
	( 14'sd 4375) * $signed(input_fmap_11[15:0]) +
	( 15'sd 13854) * $signed(input_fmap_12[15:0]) +
	( 16'sd 28565) * $signed(input_fmap_13[15:0]) +
	( 16'sd 18965) * $signed(input_fmap_14[15:0]) +
	( 16'sd 25275) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10526) * $signed(input_fmap_16[15:0]) +
	( 15'sd 11830) * $signed(input_fmap_17[15:0]) +
	( 11'sd 544) * $signed(input_fmap_18[15:0]) +
	( 15'sd 12679) * $signed(input_fmap_19[15:0]) +
	( 15'sd 11015) * $signed(input_fmap_20[15:0]) +
	( 14'sd 8027) * $signed(input_fmap_21[15:0]) +
	( 14'sd 5091) * $signed(input_fmap_22[15:0]) +
	( 16'sd 26186) * $signed(input_fmap_23[15:0]) +
	( 16'sd 31726) * $signed(input_fmap_24[15:0]) +
	( 11'sd 973) * $signed(input_fmap_25[15:0]) +
	( 14'sd 6353) * $signed(input_fmap_26[15:0]) +
	( 13'sd 3251) * $signed(input_fmap_27[15:0]) +
	( 14'sd 5630) * $signed(input_fmap_28[15:0]) +
	( 16'sd 19456) * $signed(input_fmap_29[15:0]) +
	( 16'sd 18184) * $signed(input_fmap_30[15:0]) +
	( 13'sd 2291) * $signed(input_fmap_31[15:0]) +
	( 16'sd 27432) * $signed(input_fmap_32[15:0]) +
	( 15'sd 15280) * $signed(input_fmap_33[15:0]) +
	( 15'sd 9369) * $signed(input_fmap_34[15:0]) +
	( 15'sd 15321) * $signed(input_fmap_35[15:0]) +
	( 16'sd 18717) * $signed(input_fmap_36[15:0]) +
	( 14'sd 7341) * $signed(input_fmap_37[15:0]) +
	( 10'sd 366) * $signed(input_fmap_38[15:0]) +
	( 14'sd 7112) * $signed(input_fmap_39[15:0]) +
	( 10'sd 270) * $signed(input_fmap_40[15:0]) +
	( 16'sd 27068) * $signed(input_fmap_41[15:0]) +
	( 14'sd 6234) * $signed(input_fmap_42[15:0]) +
	( 16'sd 24399) * $signed(input_fmap_43[15:0]) +
	( 15'sd 11268) * $signed(input_fmap_44[15:0]) +
	( 14'sd 4936) * $signed(input_fmap_45[15:0]) +
	( 14'sd 4480) * $signed(input_fmap_46[15:0]) +
	( 13'sd 3295) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13411) * $signed(input_fmap_48[15:0]) +
	( 16'sd 22936) * $signed(input_fmap_49[15:0]) +
	( 14'sd 5571) * $signed(input_fmap_50[15:0]) +
	( 15'sd 8559) * $signed(input_fmap_51[15:0]) +
	( 15'sd 11261) * $signed(input_fmap_52[15:0]) +
	( 13'sd 2239) * $signed(input_fmap_53[15:0]) +
	( 15'sd 14816) * $signed(input_fmap_54[15:0]) +
	( 15'sd 13780) * $signed(input_fmap_55[15:0]) +
	( 15'sd 10640) * $signed(input_fmap_56[15:0]) +
	( 9'sd 130) * $signed(input_fmap_57[15:0]) +
	( 15'sd 10581) * $signed(input_fmap_58[15:0]) +
	( 13'sd 3816) * $signed(input_fmap_59[15:0]) +
	( 16'sd 30203) * $signed(input_fmap_60[15:0]) +
	( 13'sd 3602) * $signed(input_fmap_61[15:0]) +
	( 15'sd 15734) * $signed(input_fmap_62[15:0]) +
	( 15'sd 10118) * $signed(input_fmap_63[15:0]) +
	( 14'sd 7674) * $signed(input_fmap_64[15:0]) +
	( 15'sd 9608) * $signed(input_fmap_65[15:0]) +
	( 12'sd 1199) * $signed(input_fmap_66[15:0]) +
	( 16'sd 27597) * $signed(input_fmap_67[15:0]) +
	( 16'sd 18577) * $signed(input_fmap_68[15:0]) +
	( 15'sd 11161) * $signed(input_fmap_69[15:0]) +
	( 14'sd 7892) * $signed(input_fmap_70[15:0]) +
	( 15'sd 9638) * $signed(input_fmap_71[15:0]) +
	( 15'sd 8389) * $signed(input_fmap_72[15:0]) +
	( 16'sd 20538) * $signed(input_fmap_73[15:0]) +
	( 15'sd 14843) * $signed(input_fmap_74[15:0]) +
	( 16'sd 17709) * $signed(input_fmap_75[15:0]) +
	( 15'sd 10561) * $signed(input_fmap_76[15:0]) +
	( 16'sd 28522) * $signed(input_fmap_77[15:0]) +
	( 15'sd 9252) * $signed(input_fmap_78[15:0]) +
	( 15'sd 8656) * $signed(input_fmap_79[15:0]) +
	( 16'sd 25677) * $signed(input_fmap_80[15:0]) +
	( 14'sd 4157) * $signed(input_fmap_81[15:0]) +
	( 16'sd 24795) * $signed(input_fmap_82[15:0]) +
	( 16'sd 26884) * $signed(input_fmap_83[15:0]) +
	( 16'sd 20673) * $signed(input_fmap_84[15:0]) +
	( 15'sd 13254) * $signed(input_fmap_85[15:0]) +
	( 15'sd 12015) * $signed(input_fmap_86[15:0]) +
	( 16'sd 17152) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6014) * $signed(input_fmap_88[15:0]) +
	( 16'sd 22868) * $signed(input_fmap_89[15:0]) +
	( 14'sd 5259) * $signed(input_fmap_90[15:0]) +
	( 14'sd 6729) * $signed(input_fmap_91[15:0]) +
	( 16'sd 16755) * $signed(input_fmap_92[15:0]) +
	( 16'sd 27644) * $signed(input_fmap_93[15:0]) +
	( 15'sd 12524) * $signed(input_fmap_94[15:0]) +
	( 16'sd 21263) * $signed(input_fmap_95[15:0]) +
	( 16'sd 26457) * $signed(input_fmap_96[15:0]) +
	( 16'sd 26787) * $signed(input_fmap_97[15:0]) +
	( 16'sd 18470) * $signed(input_fmap_98[15:0]) +
	( 16'sd 29033) * $signed(input_fmap_99[15:0]) +
	( 16'sd 25266) * $signed(input_fmap_100[15:0]) +
	( 16'sd 18535) * $signed(input_fmap_101[15:0]) +
	( 16'sd 18616) * $signed(input_fmap_102[15:0]) +
	( 16'sd 22974) * $signed(input_fmap_103[15:0]) +
	( 14'sd 7156) * $signed(input_fmap_104[15:0]) +
	( 14'sd 4101) * $signed(input_fmap_105[15:0]) +
	( 16'sd 29571) * $signed(input_fmap_106[15:0]) +
	( 12'sd 1474) * $signed(input_fmap_107[15:0]) +
	( 16'sd 23079) * $signed(input_fmap_108[15:0]) +
	( 15'sd 8841) * $signed(input_fmap_109[15:0]) +
	( 16'sd 18474) * $signed(input_fmap_110[15:0]) +
	( 14'sd 6137) * $signed(input_fmap_111[15:0]) +
	( 16'sd 21287) * $signed(input_fmap_112[15:0]) +
	( 16'sd 23577) * $signed(input_fmap_113[15:0]) +
	( 14'sd 7917) * $signed(input_fmap_114[15:0]) +
	( 16'sd 32334) * $signed(input_fmap_115[15:0]) +
	( 16'sd 25121) * $signed(input_fmap_116[15:0]) +
	( 14'sd 4139) * $signed(input_fmap_117[15:0]) +
	( 16'sd 19736) * $signed(input_fmap_118[15:0]) +
	( 13'sd 3415) * $signed(input_fmap_119[15:0]) +
	( 15'sd 14913) * $signed(input_fmap_120[15:0]) +
	( 16'sd 28664) * $signed(input_fmap_121[15:0]) +
	( 15'sd 14700) * $signed(input_fmap_122[15:0]) +
	( 16'sd 22273) * $signed(input_fmap_123[15:0]) +
	( 16'sd 23816) * $signed(input_fmap_124[15:0]) +
	( 16'sd 18364) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6997) * $signed(input_fmap_126[15:0]) +
	( 15'sd 9076) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 15'sd 12145) * $signed(input_fmap_0[15:0]) +
	( 16'sd 21755) * $signed(input_fmap_1[15:0]) +
	( 16'sd 30062) * $signed(input_fmap_2[15:0]) +
	( 14'sd 5818) * $signed(input_fmap_3[15:0]) +
	( 15'sd 16199) * $signed(input_fmap_4[15:0]) +
	( 16'sd 17652) * $signed(input_fmap_5[15:0]) +
	( 16'sd 29761) * $signed(input_fmap_6[15:0]) +
	( 13'sd 4018) * $signed(input_fmap_7[15:0]) +
	( 16'sd 25340) * $signed(input_fmap_8[15:0]) +
	( 15'sd 10235) * $signed(input_fmap_9[15:0]) +
	( 16'sd 20928) * $signed(input_fmap_10[15:0]) +
	( 14'sd 5805) * $signed(input_fmap_11[15:0]) +
	( 16'sd 17819) * $signed(input_fmap_12[15:0]) +
	( 13'sd 2204) * $signed(input_fmap_13[15:0]) +
	( 15'sd 13957) * $signed(input_fmap_14[15:0]) +
	( 16'sd 17523) * $signed(input_fmap_15[15:0]) +
	( 16'sd 25010) * $signed(input_fmap_16[15:0]) +
	( 16'sd 23723) * $signed(input_fmap_17[15:0]) +
	( 15'sd 8346) * $signed(input_fmap_18[15:0]) +
	( 15'sd 11709) * $signed(input_fmap_19[15:0]) +
	( 14'sd 4516) * $signed(input_fmap_20[15:0]) +
	( 15'sd 16330) * $signed(input_fmap_21[15:0]) +
	( 14'sd 7232) * $signed(input_fmap_22[15:0]) +
	( 16'sd 31569) * $signed(input_fmap_23[15:0]) +
	( 16'sd 22828) * $signed(input_fmap_24[15:0]) +
	( 16'sd 21218) * $signed(input_fmap_25[15:0]) +
	( 10'sd 466) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1255) * $signed(input_fmap_27[15:0]) +
	( 16'sd 27050) * $signed(input_fmap_28[15:0]) +
	( 15'sd 13941) * $signed(input_fmap_29[15:0]) +
	( 15'sd 11498) * $signed(input_fmap_30[15:0]) +
	( 15'sd 11593) * $signed(input_fmap_31[15:0]) +
	( 16'sd 25144) * $signed(input_fmap_32[15:0]) +
	( 13'sd 2259) * $signed(input_fmap_33[15:0]) +
	( 13'sd 3769) * $signed(input_fmap_34[15:0]) +
	( 16'sd 32530) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11495) * $signed(input_fmap_36[15:0]) +
	( 16'sd 22921) * $signed(input_fmap_37[15:0]) +
	( 15'sd 10477) * $signed(input_fmap_38[15:0]) +
	( 13'sd 2304) * $signed(input_fmap_39[15:0]) +
	( 15'sd 14077) * $signed(input_fmap_40[15:0]) +
	( 11'sd 940) * $signed(input_fmap_41[15:0]) +
	( 16'sd 24932) * $signed(input_fmap_42[15:0]) +
	( 16'sd 30212) * $signed(input_fmap_43[15:0]) +
	( 14'sd 5163) * $signed(input_fmap_44[15:0]) +
	( 14'sd 5788) * $signed(input_fmap_45[15:0]) +
	( 15'sd 15189) * $signed(input_fmap_46[15:0]) +
	( 15'sd 10519) * $signed(input_fmap_47[15:0]) +
	( 14'sd 6024) * $signed(input_fmap_48[15:0]) +
	( 13'sd 2895) * $signed(input_fmap_49[15:0]) +
	( 16'sd 28195) * $signed(input_fmap_50[15:0]) +
	( 15'sd 10027) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19890) * $signed(input_fmap_52[15:0]) +
	( 16'sd 27855) * $signed(input_fmap_53[15:0]) +
	( 16'sd 29183) * $signed(input_fmap_54[15:0]) +
	( 16'sd 20278) * $signed(input_fmap_55[15:0]) +
	( 16'sd 27645) * $signed(input_fmap_56[15:0]) +
	( 16'sd 28848) * $signed(input_fmap_57[15:0]) +
	( 14'sd 5511) * $signed(input_fmap_58[15:0]) +
	( 15'sd 10149) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1967) * $signed(input_fmap_60[15:0]) +
	( 13'sd 4037) * $signed(input_fmap_61[15:0]) +
	( 16'sd 28068) * $signed(input_fmap_62[15:0]) +
	( 16'sd 31574) * $signed(input_fmap_63[15:0]) +
	( 15'sd 12700) * $signed(input_fmap_64[15:0]) +
	( 16'sd 19923) * $signed(input_fmap_65[15:0]) +
	( 16'sd 21111) * $signed(input_fmap_66[15:0]) +
	( 16'sd 18669) * $signed(input_fmap_67[15:0]) +
	( 14'sd 7614) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31011) * $signed(input_fmap_69[15:0]) +
	( 16'sd 32348) * $signed(input_fmap_70[15:0]) +
	( 16'sd 16976) * $signed(input_fmap_71[15:0]) +
	( 12'sd 1795) * $signed(input_fmap_72[15:0]) +
	( 16'sd 30088) * $signed(input_fmap_73[15:0]) +
	( 15'sd 14680) * $signed(input_fmap_74[15:0]) +
	( 14'sd 7592) * $signed(input_fmap_75[15:0]) +
	( 12'sd 1777) * $signed(input_fmap_76[15:0]) +
	( 14'sd 5589) * $signed(input_fmap_77[15:0]) +
	( 16'sd 16857) * $signed(input_fmap_78[15:0]) +
	( 16'sd 30156) * $signed(input_fmap_79[15:0]) +
	( 16'sd 20558) * $signed(input_fmap_80[15:0]) +
	( 13'sd 3180) * $signed(input_fmap_81[15:0]) +
	( 15'sd 13378) * $signed(input_fmap_82[15:0]) +
	( 15'sd 8934) * $signed(input_fmap_83[15:0]) +
	( 14'sd 7111) * $signed(input_fmap_84[15:0]) +
	( 13'sd 2396) * $signed(input_fmap_85[15:0]) +
	( 14'sd 6171) * $signed(input_fmap_86[15:0]) +
	( 15'sd 10635) * $signed(input_fmap_87[15:0]) +
	( 14'sd 5348) * $signed(input_fmap_88[15:0]) +
	( 16'sd 17500) * $signed(input_fmap_89[15:0]) +
	( 14'sd 7958) * $signed(input_fmap_90[15:0]) +
	( 16'sd 28981) * $signed(input_fmap_91[15:0]) +
	( 16'sd 28795) * $signed(input_fmap_92[15:0]) +
	( 16'sd 27429) * $signed(input_fmap_93[15:0]) +
	( 15'sd 13777) * $signed(input_fmap_94[15:0]) +
	( 14'sd 4421) * $signed(input_fmap_95[15:0]) +
	( 15'sd 12120) * $signed(input_fmap_96[15:0]) +
	( 12'sd 1088) * $signed(input_fmap_97[15:0]) +
	( 16'sd 28766) * $signed(input_fmap_98[15:0]) +
	( 15'sd 11860) * $signed(input_fmap_99[15:0]) +
	( 16'sd 16967) * $signed(input_fmap_100[15:0]) +
	( 13'sd 2150) * $signed(input_fmap_101[15:0]) +
	( 16'sd 22163) * $signed(input_fmap_102[15:0]) +
	( 15'sd 11617) * $signed(input_fmap_103[15:0]) +
	( 11'sd 565) * $signed(input_fmap_104[15:0]) +
	( 15'sd 8358) * $signed(input_fmap_105[15:0]) +
	( 16'sd 30810) * $signed(input_fmap_106[15:0]) +
	( 14'sd 4215) * $signed(input_fmap_107[15:0]) +
	( 16'sd 24927) * $signed(input_fmap_108[15:0]) +
	( 15'sd 12008) * $signed(input_fmap_109[15:0]) +
	( 13'sd 2876) * $signed(input_fmap_110[15:0]) +
	( 16'sd 31878) * $signed(input_fmap_111[15:0]) +
	( 14'sd 5657) * $signed(input_fmap_112[15:0]) +
	( 16'sd 25056) * $signed(input_fmap_113[15:0]) +
	( 16'sd 30482) * $signed(input_fmap_114[15:0]) +
	( 16'sd 22993) * $signed(input_fmap_115[15:0]) +
	( 16'sd 16969) * $signed(input_fmap_116[15:0]) +
	( 16'sd 26427) * $signed(input_fmap_117[15:0]) +
	( 16'sd 16837) * $signed(input_fmap_118[15:0]) +
	( 16'sd 24150) * $signed(input_fmap_119[15:0]) +
	( 11'sd 826) * $signed(input_fmap_120[15:0]) +
	( 15'sd 12127) * $signed(input_fmap_121[15:0]) +
	( 16'sd 29532) * $signed(input_fmap_122[15:0]) +
	( 15'sd 11634) * $signed(input_fmap_123[15:0]) +
	( 16'sd 24381) * $signed(input_fmap_124[15:0]) +
	( 14'sd 5039) * $signed(input_fmap_125[15:0]) +
	( 16'sd 23245) * $signed(input_fmap_126[15:0]) +
	( 14'sd 7602) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 14'sd 7419) * $signed(input_fmap_0[15:0]) +
	( 16'sd 17841) * $signed(input_fmap_1[15:0]) +
	( 13'sd 2248) * $signed(input_fmap_2[15:0]) +
	( 16'sd 28230) * $signed(input_fmap_3[15:0]) +
	( 14'sd 4643) * $signed(input_fmap_4[15:0]) +
	( 16'sd 23703) * $signed(input_fmap_5[15:0]) +
	( 16'sd 18416) * $signed(input_fmap_6[15:0]) +
	( 16'sd 16531) * $signed(input_fmap_7[15:0]) +
	( 16'sd 26028) * $signed(input_fmap_8[15:0]) +
	( 12'sd 1025) * $signed(input_fmap_9[15:0]) +
	( 16'sd 26045) * $signed(input_fmap_10[15:0]) +
	( 15'sd 10443) * $signed(input_fmap_11[15:0]) +
	( 16'sd 29841) * $signed(input_fmap_12[15:0]) +
	( 16'sd 19072) * $signed(input_fmap_13[15:0]) +
	( 15'sd 15696) * $signed(input_fmap_14[15:0]) +
	( 16'sd 23052) * $signed(input_fmap_15[15:0]) +
	( 16'sd 25750) * $signed(input_fmap_16[15:0]) +
	( 15'sd 9145) * $signed(input_fmap_17[15:0]) +
	( 16'sd 27845) * $signed(input_fmap_18[15:0]) +
	( 16'sd 24238) * $signed(input_fmap_19[15:0]) +
	( 16'sd 29089) * $signed(input_fmap_20[15:0]) +
	( 16'sd 19261) * $signed(input_fmap_21[15:0]) +
	( 15'sd 10688) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24272) * $signed(input_fmap_23[15:0]) +
	( 15'sd 12635) * $signed(input_fmap_24[15:0]) +
	( 16'sd 16697) * $signed(input_fmap_25[15:0]) +
	( 13'sd 2265) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2651) * $signed(input_fmap_27[15:0]) +
	( 16'sd 28718) * $signed(input_fmap_28[15:0]) +
	( 14'sd 4930) * $signed(input_fmap_29[15:0]) +
	( 13'sd 2831) * $signed(input_fmap_30[15:0]) +
	( 16'sd 24129) * $signed(input_fmap_31[15:0]) +
	( 16'sd 23554) * $signed(input_fmap_32[15:0]) +
	( 13'sd 2276) * $signed(input_fmap_33[15:0]) +
	( 15'sd 14087) * $signed(input_fmap_34[15:0]) +
	( 15'sd 10994) * $signed(input_fmap_35[15:0]) +
	( 16'sd 23851) * $signed(input_fmap_36[15:0]) +
	( 15'sd 16085) * $signed(input_fmap_37[15:0]) +
	( 16'sd 21734) * $signed(input_fmap_38[15:0]) +
	( 15'sd 9087) * $signed(input_fmap_39[15:0]) +
	( 15'sd 13637) * $signed(input_fmap_40[15:0]) +
	( 11'sd 625) * $signed(input_fmap_41[15:0]) +
	( 16'sd 27571) * $signed(input_fmap_42[15:0]) +
	( 12'sd 1940) * $signed(input_fmap_43[15:0]) +
	( 14'sd 7772) * $signed(input_fmap_44[15:0]) +
	( 8'sd 99) * $signed(input_fmap_45[15:0]) +
	( 16'sd 20221) * $signed(input_fmap_46[15:0]) +
	( 13'sd 3997) * $signed(input_fmap_47[15:0]) +
	( 13'sd 2902) * $signed(input_fmap_48[15:0]) +
	( 15'sd 16290) * $signed(input_fmap_49[15:0]) +
	( 14'sd 5439) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15881) * $signed(input_fmap_51[15:0]) +
	( 16'sd 17762) * $signed(input_fmap_52[15:0]) +
	( 16'sd 31788) * $signed(input_fmap_53[15:0]) +
	( 16'sd 20413) * $signed(input_fmap_54[15:0]) +
	( 16'sd 26751) * $signed(input_fmap_55[15:0]) +
	( 14'sd 7567) * $signed(input_fmap_56[15:0]) +
	( 16'sd 30832) * $signed(input_fmap_57[15:0]) +
	( 15'sd 11662) * $signed(input_fmap_58[15:0]) +
	( 14'sd 7840) * $signed(input_fmap_59[15:0]) +
	( 16'sd 26201) * $signed(input_fmap_60[15:0]) +
	( 14'sd 5557) * $signed(input_fmap_61[15:0]) +
	( 15'sd 11090) * $signed(input_fmap_62[15:0]) +
	( 14'sd 5843) * $signed(input_fmap_63[15:0]) +
	( 14'sd 4939) * $signed(input_fmap_64[15:0]) +
	( 15'sd 15005) * $signed(input_fmap_65[15:0]) +
	( 16'sd 23001) * $signed(input_fmap_66[15:0]) +
	( 14'sd 7064) * $signed(input_fmap_67[15:0]) +
	( 16'sd 24340) * $signed(input_fmap_68[15:0]) +
	( 15'sd 16295) * $signed(input_fmap_69[15:0]) +
	( 16'sd 30029) * $signed(input_fmap_70[15:0]) +
	( 15'sd 10892) * $signed(input_fmap_71[15:0]) +
	( 16'sd 26503) * $signed(input_fmap_72[15:0]) +
	( 15'sd 13846) * $signed(input_fmap_73[15:0]) +
	( 15'sd 9570) * $signed(input_fmap_74[15:0]) +
	( 15'sd 11124) * $signed(input_fmap_75[15:0]) +
	( 13'sd 3738) * $signed(input_fmap_76[15:0]) +
	( 16'sd 21022) * $signed(input_fmap_77[15:0]) +
	( 13'sd 2250) * $signed(input_fmap_78[15:0]) +
	( 15'sd 13188) * $signed(input_fmap_79[15:0]) +
	( 14'sd 5647) * $signed(input_fmap_80[15:0]) +
	( 13'sd 3788) * $signed(input_fmap_81[15:0]) +
	( 15'sd 8859) * $signed(input_fmap_82[15:0]) +
	( 13'sd 3023) * $signed(input_fmap_83[15:0]) +
	( 16'sd 18447) * $signed(input_fmap_84[15:0]) +
	( 16'sd 25652) * $signed(input_fmap_85[15:0]) +
	( 14'sd 6988) * $signed(input_fmap_86[15:0]) +
	( 12'sd 1074) * $signed(input_fmap_87[15:0]) +
	( 16'sd 27572) * $signed(input_fmap_88[15:0]) +
	( 16'sd 18344) * $signed(input_fmap_89[15:0]) +
	( 16'sd 25775) * $signed(input_fmap_90[15:0]) +
	( 12'sd 1983) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25483) * $signed(input_fmap_92[15:0]) +
	( 16'sd 29316) * $signed(input_fmap_93[15:0]) +
	( 16'sd 24069) * $signed(input_fmap_94[15:0]) +
	( 14'sd 7623) * $signed(input_fmap_95[15:0]) +
	( 12'sd 1659) * $signed(input_fmap_96[15:0]) +
	( 16'sd 18046) * $signed(input_fmap_97[15:0]) +
	( 15'sd 9503) * $signed(input_fmap_98[15:0]) +
	( 15'sd 15075) * $signed(input_fmap_99[15:0]) +
	( 16'sd 18824) * $signed(input_fmap_100[15:0]) +
	( 12'sd 1683) * $signed(input_fmap_101[15:0]) +
	( 16'sd 32603) * $signed(input_fmap_102[15:0]) +
	( 14'sd 7302) * $signed(input_fmap_103[15:0]) +
	( 9'sd 249) * $signed(input_fmap_104[15:0]) +
	( 15'sd 8272) * $signed(input_fmap_105[15:0]) +
	( 16'sd 20343) * $signed(input_fmap_106[15:0]) +
	( 15'sd 8816) * $signed(input_fmap_107[15:0]) +
	( 16'sd 26518) * $signed(input_fmap_108[15:0]) +
	( 15'sd 14912) * $signed(input_fmap_109[15:0]) +
	( 15'sd 13642) * $signed(input_fmap_110[15:0]) +
	( 16'sd 25376) * $signed(input_fmap_111[15:0]) +
	( 14'sd 7997) * $signed(input_fmap_112[15:0]) +
	( 16'sd 28312) * $signed(input_fmap_113[15:0]) +
	( 16'sd 17199) * $signed(input_fmap_114[15:0]) +
	( 16'sd 31730) * $signed(input_fmap_115[15:0]) +
	( 16'sd 24229) * $signed(input_fmap_116[15:0]) +
	( 14'sd 4594) * $signed(input_fmap_117[15:0]) +
	( 15'sd 9135) * $signed(input_fmap_118[15:0]) +
	( 16'sd 24949) * $signed(input_fmap_119[15:0]) +
	( 15'sd 15203) * $signed(input_fmap_120[15:0]) +
	( 14'sd 4718) * $signed(input_fmap_121[15:0]) +
	( 12'sd 1099) * $signed(input_fmap_122[15:0]) +
	( 15'sd 9248) * $signed(input_fmap_123[15:0]) +
	( 14'sd 7145) * $signed(input_fmap_124[15:0]) +
	( 15'sd 14949) * $signed(input_fmap_125[15:0]) +
	( 16'sd 24110) * $signed(input_fmap_126[15:0]) +
	( 16'sd 24137) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 15'sd 10662) * $signed(input_fmap_0[15:0]) +
	( 15'sd 14059) * $signed(input_fmap_1[15:0]) +
	( 16'sd 23676) * $signed(input_fmap_2[15:0]) +
	( 13'sd 2897) * $signed(input_fmap_3[15:0]) +
	( 15'sd 12524) * $signed(input_fmap_4[15:0]) +
	( 14'sd 8186) * $signed(input_fmap_5[15:0]) +
	( 16'sd 32204) * $signed(input_fmap_6[15:0]) +
	( 15'sd 14363) * $signed(input_fmap_7[15:0]) +
	( 16'sd 26686) * $signed(input_fmap_8[15:0]) +
	( 13'sd 3984) * $signed(input_fmap_9[15:0]) +
	( 15'sd 14744) * $signed(input_fmap_10[15:0]) +
	( 14'sd 7317) * $signed(input_fmap_11[15:0]) +
	( 16'sd 17789) * $signed(input_fmap_12[15:0]) +
	( 14'sd 6552) * $signed(input_fmap_13[15:0]) +
	( 12'sd 1238) * $signed(input_fmap_14[15:0]) +
	( 15'sd 10197) * $signed(input_fmap_15[15:0]) +
	( 16'sd 22520) * $signed(input_fmap_16[15:0]) +
	( 16'sd 20349) * $signed(input_fmap_17[15:0]) +
	( 16'sd 17442) * $signed(input_fmap_18[15:0]) +
	( 13'sd 3203) * $signed(input_fmap_19[15:0]) +
	( 14'sd 4860) * $signed(input_fmap_20[15:0]) +
	( 12'sd 1228) * $signed(input_fmap_21[15:0]) +
	( 13'sd 3223) * $signed(input_fmap_22[15:0]) +
	( 16'sd 19801) * $signed(input_fmap_23[15:0]) +
	( 16'sd 25778) * $signed(input_fmap_24[15:0]) +
	( 13'sd 3652) * $signed(input_fmap_25[15:0]) +
	( 16'sd 26783) * $signed(input_fmap_26[15:0]) +
	( 16'sd 28890) * $signed(input_fmap_27[15:0]) +
	( 11'sd 845) * $signed(input_fmap_28[15:0]) +
	( 14'sd 7040) * $signed(input_fmap_29[15:0]) +
	( 14'sd 5486) * $signed(input_fmap_30[15:0]) +
	( 16'sd 21424) * $signed(input_fmap_31[15:0]) +
	( 15'sd 12941) * $signed(input_fmap_32[15:0]) +
	( 15'sd 15049) * $signed(input_fmap_33[15:0]) +
	( 16'sd 32327) * $signed(input_fmap_34[15:0]) +
	( 16'sd 26748) * $signed(input_fmap_35[15:0]) +
	( 15'sd 13649) * $signed(input_fmap_36[15:0]) +
	( 16'sd 32632) * $signed(input_fmap_37[15:0]) +
	( 14'sd 6444) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24317) * $signed(input_fmap_39[15:0]) +
	( 16'sd 20682) * $signed(input_fmap_40[15:0]) +
	( 15'sd 15583) * $signed(input_fmap_41[15:0]) +
	( 16'sd 26430) * $signed(input_fmap_42[15:0]) +
	( 15'sd 15701) * $signed(input_fmap_43[15:0]) +
	( 16'sd 28121) * $signed(input_fmap_44[15:0]) +
	( 16'sd 24529) * $signed(input_fmap_45[15:0]) +
	( 12'sd 1466) * $signed(input_fmap_46[15:0]) +
	( 15'sd 8225) * $signed(input_fmap_47[15:0]) +
	( 16'sd 30376) * $signed(input_fmap_48[15:0]) +
	( 16'sd 28622) * $signed(input_fmap_49[15:0]) +
	( 15'sd 10230) * $signed(input_fmap_50[15:0]) +
	( 15'sd 10145) * $signed(input_fmap_51[15:0]) +
	( 16'sd 26476) * $signed(input_fmap_52[15:0]) +
	( 12'sd 1387) * $signed(input_fmap_53[15:0]) +
	( 16'sd 24206) * $signed(input_fmap_54[15:0]) +
	( 15'sd 15368) * $signed(input_fmap_55[15:0]) +
	( 16'sd 28459) * $signed(input_fmap_56[15:0]) +
	( 14'sd 4525) * $signed(input_fmap_57[15:0]) +
	( 14'sd 5662) * $signed(input_fmap_58[15:0]) +
	( 15'sd 10943) * $signed(input_fmap_59[15:0]) +
	( 16'sd 26122) * $signed(input_fmap_60[15:0]) +
	( 16'sd 17552) * $signed(input_fmap_61[15:0]) +
	( 16'sd 21824) * $signed(input_fmap_62[15:0]) +
	( 16'sd 30368) * $signed(input_fmap_63[15:0]) +
	( 10'sd 430) * $signed(input_fmap_64[15:0]) +
	( 14'sd 6448) * $signed(input_fmap_65[15:0]) +
	( 15'sd 8499) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28977) * $signed(input_fmap_67[15:0]) +
	( 16'sd 28831) * $signed(input_fmap_68[15:0]) +
	( 16'sd 22047) * $signed(input_fmap_69[15:0]) +
	( 15'sd 8902) * $signed(input_fmap_70[15:0]) +
	( 14'sd 4705) * $signed(input_fmap_71[15:0]) +
	( 16'sd 29709) * $signed(input_fmap_72[15:0]) +
	( 16'sd 28059) * $signed(input_fmap_73[15:0]) +
	( 16'sd 32129) * $signed(input_fmap_74[15:0]) +
	( 15'sd 12127) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19205) * $signed(input_fmap_76[15:0]) +
	( 16'sd 24243) * $signed(input_fmap_77[15:0]) +
	( 15'sd 12507) * $signed(input_fmap_78[15:0]) +
	( 11'sd 593) * $signed(input_fmap_79[15:0]) +
	( 16'sd 29923) * $signed(input_fmap_80[15:0]) +
	( 15'sd 13667) * $signed(input_fmap_81[15:0]) +
	( 16'sd 25071) * $signed(input_fmap_82[15:0]) +
	( 16'sd 21990) * $signed(input_fmap_83[15:0]) +
	( 14'sd 7224) * $signed(input_fmap_84[15:0]) +
	( 13'sd 2069) * $signed(input_fmap_85[15:0]) +
	( 15'sd 11890) * $signed(input_fmap_86[15:0]) +
	( 14'sd 6865) * $signed(input_fmap_87[15:0]) +
	( 14'sd 8064) * $signed(input_fmap_88[15:0]) +
	( 16'sd 26923) * $signed(input_fmap_89[15:0]) +
	( 16'sd 26479) * $signed(input_fmap_90[15:0]) +
	( 15'sd 12466) * $signed(input_fmap_91[15:0]) +
	( 14'sd 7412) * $signed(input_fmap_92[15:0]) +
	( 16'sd 24344) * $signed(input_fmap_93[15:0]) +
	( 16'sd 23356) * $signed(input_fmap_94[15:0]) +
	( 15'sd 14073) * $signed(input_fmap_95[15:0]) +
	( 15'sd 10839) * $signed(input_fmap_96[15:0]) +
	( 16'sd 29338) * $signed(input_fmap_97[15:0]) +
	( 15'sd 10502) * $signed(input_fmap_98[15:0]) +
	( 15'sd 16198) * $signed(input_fmap_99[15:0]) +
	( 15'sd 15878) * $signed(input_fmap_100[15:0]) +
	( 13'sd 3954) * $signed(input_fmap_101[15:0]) +
	( 15'sd 12710) * $signed(input_fmap_102[15:0]) +
	( 15'sd 11387) * $signed(input_fmap_103[15:0]) +
	( 16'sd 25336) * $signed(input_fmap_104[15:0]) +
	( 16'sd 27822) * $signed(input_fmap_105[15:0]) +
	( 10'sd 361) * $signed(input_fmap_106[15:0]) +
	( 14'sd 7736) * $signed(input_fmap_107[15:0]) +
	( 16'sd 30841) * $signed(input_fmap_108[15:0]) +
	( 15'sd 9704) * $signed(input_fmap_109[15:0]) +
	( 15'sd 13780) * $signed(input_fmap_110[15:0]) +
	( 14'sd 7272) * $signed(input_fmap_111[15:0]) +
	( 14'sd 6065) * $signed(input_fmap_112[15:0]) +
	( 16'sd 30997) * $signed(input_fmap_113[15:0]) +
	( 15'sd 9276) * $signed(input_fmap_114[15:0]) +
	( 15'sd 11199) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26517) * $signed(input_fmap_116[15:0]) +
	( 9'sd 164) * $signed(input_fmap_117[15:0]) +
	( 12'sd 1125) * $signed(input_fmap_118[15:0]) +
	( 16'sd 30683) * $signed(input_fmap_119[15:0]) +
	( 16'sd 30857) * $signed(input_fmap_120[15:0]) +
	( 16'sd 26976) * $signed(input_fmap_121[15:0]) +
	( 15'sd 14458) * $signed(input_fmap_122[15:0]) +
	( 16'sd 23112) * $signed(input_fmap_123[15:0]) +
	( 16'sd 17726) * $signed(input_fmap_124[15:0]) +
	( 14'sd 5290) * $signed(input_fmap_125[15:0]) +
	( 16'sd 32007) * $signed(input_fmap_126[15:0]) +
	( 16'sd 25404) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 16'sd 24435) * $signed(input_fmap_0[15:0]) +
	( 14'sd 8102) * $signed(input_fmap_1[15:0]) +
	( 16'sd 31678) * $signed(input_fmap_2[15:0]) +
	( 16'sd 16543) * $signed(input_fmap_3[15:0]) +
	( 12'sd 2025) * $signed(input_fmap_4[15:0]) +
	( 16'sd 28445) * $signed(input_fmap_5[15:0]) +
	( 16'sd 29749) * $signed(input_fmap_6[15:0]) +
	( 11'sd 684) * $signed(input_fmap_7[15:0]) +
	( 16'sd 28990) * $signed(input_fmap_8[15:0]) +
	( 16'sd 26758) * $signed(input_fmap_9[15:0]) +
	( 15'sd 15649) * $signed(input_fmap_10[15:0]) +
	( 15'sd 14201) * $signed(input_fmap_11[15:0]) +
	( 15'sd 8612) * $signed(input_fmap_12[15:0]) +
	( 16'sd 19694) * $signed(input_fmap_13[15:0]) +
	( 15'sd 11602) * $signed(input_fmap_14[15:0]) +
	( 14'sd 7548) * $signed(input_fmap_15[15:0]) +
	( 15'sd 13022) * $signed(input_fmap_16[15:0]) +
	( 16'sd 29151) * $signed(input_fmap_17[15:0]) +
	( 16'sd 24136) * $signed(input_fmap_18[15:0]) +
	( 14'sd 4358) * $signed(input_fmap_19[15:0]) +
	( 16'sd 27849) * $signed(input_fmap_20[15:0]) +
	( 13'sd 3223) * $signed(input_fmap_21[15:0]) +
	( 15'sd 8982) * $signed(input_fmap_22[15:0]) +
	( 16'sd 17954) * $signed(input_fmap_23[15:0]) +
	( 11'sd 885) * $signed(input_fmap_24[15:0]) +
	( 16'sd 31041) * $signed(input_fmap_25[15:0]) +
	( 16'sd 31925) * $signed(input_fmap_26[15:0]) +
	( 16'sd 22623) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24734) * $signed(input_fmap_28[15:0]) +
	( 16'sd 16469) * $signed(input_fmap_29[15:0]) +
	( 16'sd 29649) * $signed(input_fmap_30[15:0]) +
	( 16'sd 29185) * $signed(input_fmap_31[15:0]) +
	( 15'sd 10744) * $signed(input_fmap_32[15:0]) +
	( 16'sd 30928) * $signed(input_fmap_33[15:0]) +
	( 15'sd 15907) * $signed(input_fmap_34[15:0]) +
	( 16'sd 29013) * $signed(input_fmap_35[15:0]) +
	( 15'sd 14621) * $signed(input_fmap_36[15:0]) +
	( 16'sd 21873) * $signed(input_fmap_37[15:0]) +
	( 16'sd 24182) * $signed(input_fmap_38[15:0]) +
	( 16'sd 32118) * $signed(input_fmap_39[15:0]) +
	( 15'sd 11716) * $signed(input_fmap_40[15:0]) +
	( 16'sd 30418) * $signed(input_fmap_41[15:0]) +
	( 16'sd 28901) * $signed(input_fmap_42[15:0]) +
	( 15'sd 8459) * $signed(input_fmap_43[15:0]) +
	( 14'sd 6569) * $signed(input_fmap_44[15:0]) +
	( 15'sd 10854) * $signed(input_fmap_45[15:0]) +
	( 15'sd 15721) * $signed(input_fmap_46[15:0]) +
	( 14'sd 7189) * $signed(input_fmap_47[15:0]) +
	( 16'sd 25771) * $signed(input_fmap_48[15:0]) +
	( 15'sd 16212) * $signed(input_fmap_49[15:0]) +
	( 13'sd 3980) * $signed(input_fmap_50[15:0]) +
	( 14'sd 7154) * $signed(input_fmap_51[15:0]) +
	( 15'sd 16338) * $signed(input_fmap_52[15:0]) +
	( 15'sd 15848) * $signed(input_fmap_53[15:0]) +
	( 16'sd 25830) * $signed(input_fmap_54[15:0]) +
	( 16'sd 20843) * $signed(input_fmap_55[15:0]) +
	( 15'sd 12676) * $signed(input_fmap_56[15:0]) +
	( 15'sd 8356) * $signed(input_fmap_57[15:0]) +
	( 15'sd 14418) * $signed(input_fmap_58[15:0]) +
	( 16'sd 27236) * $signed(input_fmap_59[15:0]) +
	( 14'sd 7962) * $signed(input_fmap_60[15:0]) +
	( 16'sd 21036) * $signed(input_fmap_61[15:0]) +
	( 14'sd 5309) * $signed(input_fmap_62[15:0]) +
	( 14'sd 7127) * $signed(input_fmap_63[15:0]) +
	( 16'sd 30550) * $signed(input_fmap_64[15:0]) +
	( 15'sd 14388) * $signed(input_fmap_65[15:0]) +
	( 16'sd 32716) * $signed(input_fmap_66[15:0]) +
	( 16'sd 22764) * $signed(input_fmap_67[15:0]) +
	( 16'sd 31585) * $signed(input_fmap_68[15:0]) +
	( 12'sd 1353) * $signed(input_fmap_69[15:0]) +
	( 16'sd 25521) * $signed(input_fmap_70[15:0]) +
	( 16'sd 22384) * $signed(input_fmap_71[15:0]) +
	( 16'sd 21075) * $signed(input_fmap_72[15:0]) +
	( 15'sd 15096) * $signed(input_fmap_73[15:0]) +
	( 16'sd 17505) * $signed(input_fmap_74[15:0]) +
	( 14'sd 5637) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19986) * $signed(input_fmap_76[15:0]) +
	( 14'sd 7853) * $signed(input_fmap_77[15:0]) +
	( 16'sd 19065) * $signed(input_fmap_78[15:0]) +
	( 15'sd 14526) * $signed(input_fmap_79[15:0]) +
	( 16'sd 30607) * $signed(input_fmap_80[15:0]) +
	( 16'sd 26217) * $signed(input_fmap_81[15:0]) +
	( 16'sd 29214) * $signed(input_fmap_82[15:0]) +
	( 16'sd 30110) * $signed(input_fmap_83[15:0]) +
	( 16'sd 21428) * $signed(input_fmap_84[15:0]) +
	( 13'sd 3668) * $signed(input_fmap_85[15:0]) +
	( 14'sd 7452) * $signed(input_fmap_86[15:0]) +
	( 15'sd 9692) * $signed(input_fmap_87[15:0]) +
	( 15'sd 10284) * $signed(input_fmap_88[15:0]) +
	( 16'sd 25305) * $signed(input_fmap_89[15:0]) +
	( 15'sd 13882) * $signed(input_fmap_90[15:0]) +
	( 16'sd 22498) * $signed(input_fmap_91[15:0]) +
	( 16'sd 24654) * $signed(input_fmap_92[15:0]) +
	( 16'sd 29625) * $signed(input_fmap_93[15:0]) +
	( 12'sd 1071) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25428) * $signed(input_fmap_95[15:0]) +
	( 16'sd 19073) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27347) * $signed(input_fmap_97[15:0]) +
	( 15'sd 12151) * $signed(input_fmap_98[15:0]) +
	( 16'sd 26522) * $signed(input_fmap_99[15:0]) +
	( 15'sd 14181) * $signed(input_fmap_100[15:0]) +
	( 15'sd 14314) * $signed(input_fmap_101[15:0]) +
	( 16'sd 19887) * $signed(input_fmap_102[15:0]) +
	( 16'sd 17642) * $signed(input_fmap_103[15:0]) +
	( 16'sd 17641) * $signed(input_fmap_104[15:0]) +
	( 14'sd 7302) * $signed(input_fmap_105[15:0]) +
	( 16'sd 21342) * $signed(input_fmap_106[15:0]) +
	( 16'sd 16604) * $signed(input_fmap_107[15:0]) +
	( 16'sd 32050) * $signed(input_fmap_108[15:0]) +
	( 15'sd 10690) * $signed(input_fmap_109[15:0]) +
	( 16'sd 27265) * $signed(input_fmap_110[15:0]) +
	( 16'sd 16893) * $signed(input_fmap_111[15:0]) +
	( 14'sd 4267) * $signed(input_fmap_112[15:0]) +
	( 16'sd 29905) * $signed(input_fmap_113[15:0]) +
	( 13'sd 2467) * $signed(input_fmap_114[15:0]) +
	( 16'sd 28632) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15087) * $signed(input_fmap_116[15:0]) +
	( 16'sd 26452) * $signed(input_fmap_117[15:0]) +
	( 16'sd 22349) * $signed(input_fmap_118[15:0]) +
	( 16'sd 26350) * $signed(input_fmap_119[15:0]) +
	( 11'sd 564) * $signed(input_fmap_120[15:0]) +
	( 16'sd 28349) * $signed(input_fmap_121[15:0]) +
	( 14'sd 7890) * $signed(input_fmap_122[15:0]) +
	( 15'sd 14962) * $signed(input_fmap_123[15:0]) +
	( 15'sd 12653) * $signed(input_fmap_124[15:0]) +
	( 16'sd 28718) * $signed(input_fmap_125[15:0]) +
	( 16'sd 20587) * $signed(input_fmap_126[15:0]) +
	( 15'sd 8262) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 16'sd 18638) * $signed(input_fmap_0[15:0]) +
	( 16'sd 22224) * $signed(input_fmap_1[15:0]) +
	( 13'sd 2371) * $signed(input_fmap_2[15:0]) +
	( 13'sd 4005) * $signed(input_fmap_3[15:0]) +
	( 16'sd 17569) * $signed(input_fmap_4[15:0]) +
	( 11'sd 744) * $signed(input_fmap_5[15:0]) +
	( 16'sd 21191) * $signed(input_fmap_6[15:0]) +
	( 16'sd 29208) * $signed(input_fmap_7[15:0]) +
	( 13'sd 2257) * $signed(input_fmap_8[15:0]) +
	( 16'sd 25153) * $signed(input_fmap_9[15:0]) +
	( 16'sd 28690) * $signed(input_fmap_10[15:0]) +
	( 16'sd 28766) * $signed(input_fmap_11[15:0]) +
	( 16'sd 31377) * $signed(input_fmap_12[15:0]) +
	( 12'sd 1368) * $signed(input_fmap_13[15:0]) +
	( 16'sd 20935) * $signed(input_fmap_14[15:0]) +
	( 14'sd 7692) * $signed(input_fmap_15[15:0]) +
	( 15'sd 12683) * $signed(input_fmap_16[15:0]) +
	( 16'sd 26414) * $signed(input_fmap_17[15:0]) +
	( 14'sd 6349) * $signed(input_fmap_18[15:0]) +
	( 16'sd 21372) * $signed(input_fmap_19[15:0]) +
	( 13'sd 3381) * $signed(input_fmap_20[15:0]) +
	( 15'sd 12743) * $signed(input_fmap_21[15:0]) +
	( 16'sd 20756) * $signed(input_fmap_22[15:0]) +
	( 16'sd 31533) * $signed(input_fmap_23[15:0]) +
	( 16'sd 28826) * $signed(input_fmap_24[15:0]) +
	( 16'sd 29900) * $signed(input_fmap_25[15:0]) +
	( 13'sd 3567) * $signed(input_fmap_26[15:0]) +
	( 16'sd 32709) * $signed(input_fmap_27[15:0]) +
	( 16'sd 30373) * $signed(input_fmap_28[15:0]) +
	( 16'sd 25802) * $signed(input_fmap_29[15:0]) +
	( 16'sd 22261) * $signed(input_fmap_30[15:0]) +
	( 16'sd 28492) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28118) * $signed(input_fmap_32[15:0]) +
	( 15'sd 11805) * $signed(input_fmap_33[15:0]) +
	( 13'sd 3599) * $signed(input_fmap_34[15:0]) +
	( 15'sd 13164) * $signed(input_fmap_35[15:0]) +
	( 14'sd 4540) * $signed(input_fmap_36[15:0]) +
	( 16'sd 24180) * $signed(input_fmap_37[15:0]) +
	( 16'sd 32005) * $signed(input_fmap_38[15:0]) +
	( 16'sd 31094) * $signed(input_fmap_39[15:0]) +
	( 16'sd 26035) * $signed(input_fmap_40[15:0]) +
	( 15'sd 8743) * $signed(input_fmap_41[15:0]) +
	( 16'sd 24548) * $signed(input_fmap_42[15:0]) +
	( 15'sd 15383) * $signed(input_fmap_43[15:0]) +
	( 15'sd 9682) * $signed(input_fmap_44[15:0]) +
	( 15'sd 9233) * $signed(input_fmap_45[15:0]) +
	( 16'sd 25633) * $signed(input_fmap_46[15:0]) +
	( 16'sd 28230) * $signed(input_fmap_47[15:0]) +
	( 16'sd 21601) * $signed(input_fmap_48[15:0]) +
	( 16'sd 27216) * $signed(input_fmap_49[15:0]) +
	( 15'sd 13792) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15454) * $signed(input_fmap_51[15:0]) +
	( 15'sd 8306) * $signed(input_fmap_52[15:0]) +
	( 16'sd 23564) * $signed(input_fmap_53[15:0]) +
	( 13'sd 2630) * $signed(input_fmap_54[15:0]) +
	( 15'sd 9296) * $signed(input_fmap_55[15:0]) +
	( 16'sd 29414) * $signed(input_fmap_56[15:0]) +
	( 16'sd 18885) * $signed(input_fmap_57[15:0]) +
	( 16'sd 24371) * $signed(input_fmap_58[15:0]) +
	( 15'sd 11893) * $signed(input_fmap_59[15:0]) +
	( 14'sd 5341) * $signed(input_fmap_60[15:0]) +
	( 15'sd 9262) * $signed(input_fmap_61[15:0]) +
	( 16'sd 21704) * $signed(input_fmap_62[15:0]) +
	( 15'sd 8640) * $signed(input_fmap_63[15:0]) +
	( 14'sd 7249) * $signed(input_fmap_64[15:0]) +
	( 16'sd 22692) * $signed(input_fmap_65[15:0]) +
	( 16'sd 26123) * $signed(input_fmap_66[15:0]) +
	( 16'sd 30569) * $signed(input_fmap_67[15:0]) +
	( 15'sd 10582) * $signed(input_fmap_68[15:0]) +
	( 15'sd 12649) * $signed(input_fmap_69[15:0]) +
	( 16'sd 21595) * $signed(input_fmap_70[15:0]) +
	( 16'sd 24518) * $signed(input_fmap_71[15:0]) +
	( 15'sd 15219) * $signed(input_fmap_72[15:0]) +
	( 16'sd 19202) * $signed(input_fmap_73[15:0]) +
	( 15'sd 10996) * $signed(input_fmap_74[15:0]) +
	( 15'sd 12909) * $signed(input_fmap_75[15:0]) +
	( 16'sd 29534) * $signed(input_fmap_76[15:0]) +
	( 16'sd 16875) * $signed(input_fmap_77[15:0]) +
	( 13'sd 2688) * $signed(input_fmap_78[15:0]) +
	( 16'sd 30454) * $signed(input_fmap_79[15:0]) +
	( 11'sd 682) * $signed(input_fmap_80[15:0]) +
	( 15'sd 12049) * $signed(input_fmap_81[15:0]) +
	( 16'sd 27931) * $signed(input_fmap_82[15:0]) +
	( 16'sd 22803) * $signed(input_fmap_83[15:0]) +
	( 16'sd 16453) * $signed(input_fmap_84[15:0]) +
	( 14'sd 5304) * $signed(input_fmap_85[15:0]) +
	( 15'sd 14674) * $signed(input_fmap_86[15:0]) +
	( 16'sd 28694) * $signed(input_fmap_87[15:0]) +
	( 15'sd 16289) * $signed(input_fmap_88[15:0]) +
	( 16'sd 24529) * $signed(input_fmap_89[15:0]) +
	( 15'sd 15508) * $signed(input_fmap_90[15:0]) +
	( 15'sd 12066) * $signed(input_fmap_91[15:0]) +
	( 15'sd 8999) * $signed(input_fmap_92[15:0]) +
	( 16'sd 30791) * $signed(input_fmap_93[15:0]) +
	( 16'sd 23110) * $signed(input_fmap_94[15:0]) +
	( 15'sd 10928) * $signed(input_fmap_95[15:0]) +
	( 13'sd 3222) * $signed(input_fmap_96[15:0]) +
	( 15'sd 12334) * $signed(input_fmap_97[15:0]) +
	( 15'sd 12726) * $signed(input_fmap_98[15:0]) +
	( 11'sd 670) * $signed(input_fmap_99[15:0]) +
	( 15'sd 12533) * $signed(input_fmap_100[15:0]) +
	( 16'sd 22273) * $signed(input_fmap_101[15:0]) +
	( 14'sd 4727) * $signed(input_fmap_102[15:0]) +
	( 16'sd 27632) * $signed(input_fmap_103[15:0]) +
	( 16'sd 24444) * $signed(input_fmap_104[15:0]) +
	( 16'sd 28903) * $signed(input_fmap_105[15:0]) +
	( 16'sd 23211) * $signed(input_fmap_106[15:0]) +
	( 16'sd 17713) * $signed(input_fmap_107[15:0]) +
	( 15'sd 13419) * $signed(input_fmap_108[15:0]) +
	( 15'sd 14979) * $signed(input_fmap_109[15:0]) +
	( 16'sd 19373) * $signed(input_fmap_110[15:0]) +
	( 14'sd 5740) * $signed(input_fmap_111[15:0]) +
	( 14'sd 4807) * $signed(input_fmap_112[15:0]) +
	( 14'sd 8116) * $signed(input_fmap_113[15:0]) +
	( 16'sd 28360) * $signed(input_fmap_114[15:0]) +
	( 15'sd 9332) * $signed(input_fmap_115[15:0]) +
	( 16'sd 22419) * $signed(input_fmap_116[15:0]) +
	( 15'sd 10953) * $signed(input_fmap_117[15:0]) +
	( 15'sd 8729) * $signed(input_fmap_118[15:0]) +
	( 15'sd 12805) * $signed(input_fmap_119[15:0]) +
	( 12'sd 2016) * $signed(input_fmap_120[15:0]) +
	( 16'sd 22732) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9535) * $signed(input_fmap_122[15:0]) +
	( 14'sd 5840) * $signed(input_fmap_123[15:0]) +
	( 12'sd 1304) * $signed(input_fmap_124[15:0]) +
	( 15'sd 9487) * $signed(input_fmap_125[15:0]) +
	( 13'sd 3433) * $signed(input_fmap_126[15:0]) +
	( 15'sd 15412) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 14'sd 7498) * $signed(input_fmap_0[15:0]) +
	( 16'sd 28801) * $signed(input_fmap_1[15:0]) +
	( 12'sd 1187) * $signed(input_fmap_2[15:0]) +
	( 16'sd 22228) * $signed(input_fmap_3[15:0]) +
	( 16'sd 27607) * $signed(input_fmap_4[15:0]) +
	( 16'sd 21168) * $signed(input_fmap_5[15:0]) +
	( 14'sd 7671) * $signed(input_fmap_6[15:0]) +
	( 15'sd 9698) * $signed(input_fmap_7[15:0]) +
	( 14'sd 4793) * $signed(input_fmap_8[15:0]) +
	( 15'sd 16021) * $signed(input_fmap_9[15:0]) +
	( 13'sd 2171) * $signed(input_fmap_10[15:0]) +
	( 15'sd 10061) * $signed(input_fmap_11[15:0]) +
	( 16'sd 21627) * $signed(input_fmap_12[15:0]) +
	( 15'sd 8280) * $signed(input_fmap_13[15:0]) +
	( 16'sd 26285) * $signed(input_fmap_14[15:0]) +
	( 13'sd 4041) * $signed(input_fmap_15[15:0]) +
	( 16'sd 31481) * $signed(input_fmap_16[15:0]) +
	( 14'sd 6569) * $signed(input_fmap_17[15:0]) +
	( 16'sd 24371) * $signed(input_fmap_18[15:0]) +
	( 15'sd 10336) * $signed(input_fmap_19[15:0]) +
	( 13'sd 4060) * $signed(input_fmap_20[15:0]) +
	( 16'sd 30989) * $signed(input_fmap_21[15:0]) +
	( 16'sd 32099) * $signed(input_fmap_22[15:0]) +
	( 15'sd 15673) * $signed(input_fmap_23[15:0]) +
	( 14'sd 7761) * $signed(input_fmap_24[15:0]) +
	( 16'sd 19218) * $signed(input_fmap_25[15:0]) +
	( 11'sd 667) * $signed(input_fmap_26[15:0]) +
	( 16'sd 30513) * $signed(input_fmap_27[15:0]) +
	( 14'sd 5115) * $signed(input_fmap_28[15:0]) +
	( 15'sd 14359) * $signed(input_fmap_29[15:0]) +
	( 13'sd 2365) * $signed(input_fmap_30[15:0]) +
	( 16'sd 31270) * $signed(input_fmap_31[15:0]) +
	( 15'sd 11380) * $signed(input_fmap_32[15:0]) +
	( 15'sd 9237) * $signed(input_fmap_33[15:0]) +
	( 14'sd 7264) * $signed(input_fmap_34[15:0]) +
	( 16'sd 17898) * $signed(input_fmap_35[15:0]) +
	( 15'sd 12230) * $signed(input_fmap_36[15:0]) +
	( 16'sd 24514) * $signed(input_fmap_37[15:0]) +
	( 13'sd 3201) * $signed(input_fmap_38[15:0]) +
	( 16'sd 23392) * $signed(input_fmap_39[15:0]) +
	( 14'sd 7488) * $signed(input_fmap_40[15:0]) +
	( 16'sd 31044) * $signed(input_fmap_41[15:0]) +
	( 16'sd 24819) * $signed(input_fmap_42[15:0]) +
	( 16'sd 26114) * $signed(input_fmap_43[15:0]) +
	( 16'sd 17801) * $signed(input_fmap_44[15:0]) +
	( 16'sd 21882) * $signed(input_fmap_45[15:0]) +
	( 16'sd 29023) * $signed(input_fmap_46[15:0]) +
	( 16'sd 21428) * $signed(input_fmap_47[15:0]) +
	( 13'sd 3291) * $signed(input_fmap_48[15:0]) +
	( 15'sd 10084) * $signed(input_fmap_49[15:0]) +
	( 16'sd 28164) * $signed(input_fmap_50[15:0]) +
	( 16'sd 20974) * $signed(input_fmap_51[15:0]) +
	( 16'sd 20247) * $signed(input_fmap_52[15:0]) +
	( 16'sd 29108) * $signed(input_fmap_53[15:0]) +
	( 16'sd 29222) * $signed(input_fmap_54[15:0]) +
	( 15'sd 9284) * $signed(input_fmap_55[15:0]) +
	( 16'sd 27147) * $signed(input_fmap_56[15:0]) +
	( 15'sd 8886) * $signed(input_fmap_57[15:0]) +
	( 14'sd 7163) * $signed(input_fmap_58[15:0]) +
	( 14'sd 7194) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1730) * $signed(input_fmap_60[15:0]) +
	( 16'sd 28690) * $signed(input_fmap_61[15:0]) +
	( 16'sd 31924) * $signed(input_fmap_62[15:0]) +
	( 16'sd 19881) * $signed(input_fmap_63[15:0]) +
	( 15'sd 12807) * $signed(input_fmap_64[15:0]) +
	( 16'sd 16779) * $signed(input_fmap_65[15:0]) +
	( 16'sd 27087) * $signed(input_fmap_66[15:0]) +
	( 16'sd 23917) * $signed(input_fmap_67[15:0]) +
	( 15'sd 14627) * $signed(input_fmap_68[15:0]) +
	( 16'sd 27330) * $signed(input_fmap_69[15:0]) +
	( 16'sd 18627) * $signed(input_fmap_70[15:0]) +
	( 16'sd 20166) * $signed(input_fmap_71[15:0]) +
	( 14'sd 7807) * $signed(input_fmap_72[15:0]) +
	( 14'sd 6730) * $signed(input_fmap_73[15:0]) +
	( 16'sd 25469) * $signed(input_fmap_74[15:0]) +
	( 15'sd 11305) * $signed(input_fmap_75[15:0]) +
	( 15'sd 13272) * $signed(input_fmap_76[15:0]) +
	( 14'sd 4692) * $signed(input_fmap_77[15:0]) +
	( 16'sd 25204) * $signed(input_fmap_78[15:0]) +
	( 16'sd 25248) * $signed(input_fmap_79[15:0]) +
	( 16'sd 23327) * $signed(input_fmap_80[15:0]) +
	( 15'sd 8251) * $signed(input_fmap_81[15:0]) +
	( 16'sd 21439) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25241) * $signed(input_fmap_83[15:0]) +
	( 16'sd 31275) * $signed(input_fmap_84[15:0]) +
	( 16'sd 29973) * $signed(input_fmap_85[15:0]) +
	( 16'sd 21558) * $signed(input_fmap_86[15:0]) +
	( 16'sd 25227) * $signed(input_fmap_87[15:0]) +
	( 15'sd 13368) * $signed(input_fmap_88[15:0]) +
	( 14'sd 7742) * $signed(input_fmap_89[15:0]) +
	( 16'sd 31750) * $signed(input_fmap_90[15:0]) +
	( 16'sd 24382) * $signed(input_fmap_91[15:0]) +
	( 15'sd 11255) * $signed(input_fmap_92[15:0]) +
	( 16'sd 26722) * $signed(input_fmap_93[15:0]) +
	( 16'sd 25577) * $signed(input_fmap_94[15:0]) +
	( 16'sd 26956) * $signed(input_fmap_95[15:0]) +
	( 16'sd 26109) * $signed(input_fmap_96[15:0]) +
	( 16'sd 16618) * $signed(input_fmap_97[15:0]) +
	( 14'sd 7323) * $signed(input_fmap_98[15:0]) +
	( 15'sd 14759) * $signed(input_fmap_99[15:0]) +
	( 16'sd 27885) * $signed(input_fmap_100[15:0]) +
	( 15'sd 14896) * $signed(input_fmap_101[15:0]) +
	( 14'sd 8076) * $signed(input_fmap_102[15:0]) +
	( 16'sd 30817) * $signed(input_fmap_103[15:0]) +
	( 16'sd 27772) * $signed(input_fmap_104[15:0]) +
	( 14'sd 4604) * $signed(input_fmap_105[15:0]) +
	( 16'sd 17514) * $signed(input_fmap_106[15:0]) +
	( 15'sd 11657) * $signed(input_fmap_107[15:0]) +
	( 12'sd 1803) * $signed(input_fmap_108[15:0]) +
	( 16'sd 24906) * $signed(input_fmap_109[15:0]) +
	( 16'sd 27623) * $signed(input_fmap_110[15:0]) +
	( 13'sd 2654) * $signed(input_fmap_111[15:0]) +
	( 16'sd 23152) * $signed(input_fmap_112[15:0]) +
	( 16'sd 25233) * $signed(input_fmap_113[15:0]) +
	( 15'sd 8605) * $signed(input_fmap_114[15:0]) +
	( 15'sd 10155) * $signed(input_fmap_115[15:0]) +
	( 14'sd 7668) * $signed(input_fmap_116[15:0]) +
	( 16'sd 32268) * $signed(input_fmap_117[15:0]) +
	( 16'sd 31080) * $signed(input_fmap_118[15:0]) +
	( 15'sd 14613) * $signed(input_fmap_119[15:0]) +
	( 16'sd 28870) * $signed(input_fmap_120[15:0]) +
	( 16'sd 20185) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9780) * $signed(input_fmap_122[15:0]) +
	( 16'sd 28987) * $signed(input_fmap_123[15:0]) +
	( 16'sd 25898) * $signed(input_fmap_124[15:0]) +
	( 16'sd 30400) * $signed(input_fmap_125[15:0]) +
	( 15'sd 9103) * $signed(input_fmap_126[15:0]) +
	( 16'sd 24268) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 15'sd 12565) * $signed(input_fmap_0[15:0]) +
	( 16'sd 21652) * $signed(input_fmap_1[15:0]) +
	( 15'sd 9359) * $signed(input_fmap_2[15:0]) +
	( 15'sd 14462) * $signed(input_fmap_3[15:0]) +
	( 16'sd 24278) * $signed(input_fmap_4[15:0]) +
	( 15'sd 10720) * $signed(input_fmap_5[15:0]) +
	( 13'sd 3952) * $signed(input_fmap_6[15:0]) +
	( 16'sd 32513) * $signed(input_fmap_7[15:0]) +
	( 15'sd 14738) * $signed(input_fmap_8[15:0]) +
	( 16'sd 22242) * $signed(input_fmap_9[15:0]) +
	( 16'sd 22353) * $signed(input_fmap_10[15:0]) +
	( 14'sd 5439) * $signed(input_fmap_11[15:0]) +
	( 15'sd 13867) * $signed(input_fmap_12[15:0]) +
	( 15'sd 13103) * $signed(input_fmap_13[15:0]) +
	( 16'sd 27318) * $signed(input_fmap_14[15:0]) +
	( 16'sd 24188) * $signed(input_fmap_15[15:0]) +
	( 16'sd 23685) * $signed(input_fmap_16[15:0]) +
	( 15'sd 8696) * $signed(input_fmap_17[15:0]) +
	( 15'sd 14377) * $signed(input_fmap_18[15:0]) +
	( 16'sd 29001) * $signed(input_fmap_19[15:0]) +
	( 16'sd 31198) * $signed(input_fmap_20[15:0]) +
	( 14'sd 4524) * $signed(input_fmap_21[15:0]) +
	( 16'sd 28492) * $signed(input_fmap_22[15:0]) +
	( 14'sd 5577) * $signed(input_fmap_23[15:0]) +
	( 15'sd 12696) * $signed(input_fmap_24[15:0]) +
	( 16'sd 31283) * $signed(input_fmap_25[15:0]) +
	( 16'sd 18065) * $signed(input_fmap_26[15:0]) +
	( 16'sd 22932) * $signed(input_fmap_27[15:0]) +
	( 16'sd 20427) * $signed(input_fmap_28[15:0]) +
	( 16'sd 17599) * $signed(input_fmap_29[15:0]) +
	( 14'sd 6269) * $signed(input_fmap_30[15:0]) +
	( 16'sd 28290) * $signed(input_fmap_31[15:0]) +
	( 16'sd 29130) * $signed(input_fmap_32[15:0]) +
	( 12'sd 1677) * $signed(input_fmap_33[15:0]) +
	( 16'sd 29354) * $signed(input_fmap_34[15:0]) +
	( 16'sd 24976) * $signed(input_fmap_35[15:0]) +
	( 16'sd 24301) * $signed(input_fmap_36[15:0]) +
	( 16'sd 30499) * $signed(input_fmap_37[15:0]) +
	( 15'sd 11976) * $signed(input_fmap_38[15:0]) +
	( 16'sd 31112) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6343) * $signed(input_fmap_40[15:0]) +
	( 15'sd 9024) * $signed(input_fmap_41[15:0]) +
	( 14'sd 6116) * $signed(input_fmap_42[15:0]) +
	( 15'sd 12669) * $signed(input_fmap_43[15:0]) +
	( 15'sd 9234) * $signed(input_fmap_44[15:0]) +
	( 16'sd 25531) * $signed(input_fmap_45[15:0]) +
	( 15'sd 9167) * $signed(input_fmap_46[15:0]) +
	( 16'sd 31778) * $signed(input_fmap_47[15:0]) +
	( 10'sd 309) * $signed(input_fmap_48[15:0]) +
	( 15'sd 9673) * $signed(input_fmap_49[15:0]) +
	( 16'sd 24241) * $signed(input_fmap_50[15:0]) +
	( 15'sd 13993) * $signed(input_fmap_51[15:0]) +
	( 16'sd 21069) * $signed(input_fmap_52[15:0]) +
	( 16'sd 26913) * $signed(input_fmap_53[15:0]) +
	( 16'sd 31831) * $signed(input_fmap_54[15:0]) +
	( 14'sd 4479) * $signed(input_fmap_55[15:0]) +
	( 8'sd 117) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17713) * $signed(input_fmap_57[15:0]) +
	( 16'sd 19353) * $signed(input_fmap_58[15:0]) +
	( 16'sd 17670) * $signed(input_fmap_59[15:0]) +
	( 14'sd 5897) * $signed(input_fmap_60[15:0]) +
	( 16'sd 23443) * $signed(input_fmap_61[15:0]) +
	( 10'sd 358) * $signed(input_fmap_62[15:0]) +
	( 15'sd 15111) * $signed(input_fmap_63[15:0]) +
	( 14'sd 4464) * $signed(input_fmap_64[15:0]) +
	( 16'sd 25709) * $signed(input_fmap_65[15:0]) +
	( 16'sd 32257) * $signed(input_fmap_66[15:0]) +
	( 15'sd 12363) * $signed(input_fmap_67[15:0]) +
	( 15'sd 13286) * $signed(input_fmap_68[15:0]) +
	( 16'sd 23883) * $signed(input_fmap_69[15:0]) +
	( 13'sd 2665) * $signed(input_fmap_70[15:0]) +
	( 16'sd 18366) * $signed(input_fmap_71[15:0]) +
	( 16'sd 20721) * $signed(input_fmap_72[15:0]) +
	( 16'sd 24783) * $signed(input_fmap_73[15:0]) +
	( 16'sd 32142) * $signed(input_fmap_74[15:0]) +
	( 16'sd 29422) * $signed(input_fmap_75[15:0]) +
	( 16'sd 25360) * $signed(input_fmap_76[15:0]) +
	( 16'sd 31056) * $signed(input_fmap_77[15:0]) +
	( 15'sd 15334) * $signed(input_fmap_78[15:0]) +
	( 16'sd 29422) * $signed(input_fmap_79[15:0]) +
	( 16'sd 29080) * $signed(input_fmap_80[15:0]) +
	( 16'sd 23800) * $signed(input_fmap_81[15:0]) +
	( 16'sd 18222) * $signed(input_fmap_82[15:0]) +
	( 16'sd 31094) * $signed(input_fmap_83[15:0]) +
	( 16'sd 23991) * $signed(input_fmap_84[15:0]) +
	( 15'sd 15360) * $signed(input_fmap_85[15:0]) +
	( 16'sd 28269) * $signed(input_fmap_86[15:0]) +
	( 16'sd 31050) * $signed(input_fmap_87[15:0]) +
	( 14'sd 5644) * $signed(input_fmap_88[15:0]) +
	( 16'sd 19952) * $signed(input_fmap_89[15:0]) +
	( 14'sd 8087) * $signed(input_fmap_90[15:0]) +
	( 13'sd 3505) * $signed(input_fmap_91[15:0]) +
	( 16'sd 28982) * $signed(input_fmap_92[15:0]) +
	( 15'sd 10312) * $signed(input_fmap_93[15:0]) +
	( 16'sd 26025) * $signed(input_fmap_94[15:0]) +
	( 14'sd 4761) * $signed(input_fmap_95[15:0]) +
	( 16'sd 30499) * $signed(input_fmap_96[15:0]) +
	( 16'sd 28131) * $signed(input_fmap_97[15:0]) +
	( 16'sd 17313) * $signed(input_fmap_98[15:0]) +
	( 14'sd 7787) * $signed(input_fmap_99[15:0]) +
	( 15'sd 8303) * $signed(input_fmap_100[15:0]) +
	( 15'sd 9708) * $signed(input_fmap_101[15:0]) +
	( 15'sd 10446) * $signed(input_fmap_102[15:0]) +
	( 15'sd 15184) * $signed(input_fmap_103[15:0]) +
	( 16'sd 31598) * $signed(input_fmap_104[15:0]) +
	( 16'sd 32321) * $signed(input_fmap_105[15:0]) +
	( 16'sd 21810) * $signed(input_fmap_106[15:0]) +
	( 16'sd 24390) * $signed(input_fmap_107[15:0]) +
	( 16'sd 23535) * $signed(input_fmap_108[15:0]) +
	( 16'sd 20447) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22807) * $signed(input_fmap_110[15:0]) +
	( 14'sd 7623) * $signed(input_fmap_111[15:0]) +
	( 16'sd 24871) * $signed(input_fmap_112[15:0]) +
	( 14'sd 6804) * $signed(input_fmap_113[15:0]) +
	( 15'sd 15211) * $signed(input_fmap_114[15:0]) +
	( 14'sd 6647) * $signed(input_fmap_115[15:0]) +
	( 16'sd 32636) * $signed(input_fmap_116[15:0]) +
	( 16'sd 21094) * $signed(input_fmap_117[15:0]) +
	( 16'sd 26160) * $signed(input_fmap_118[15:0]) +
	( 16'sd 22766) * $signed(input_fmap_119[15:0]) +
	( 15'sd 10019) * $signed(input_fmap_120[15:0]) +
	( 16'sd 25320) * $signed(input_fmap_121[15:0]) +
	( 16'sd 22939) * $signed(input_fmap_122[15:0]) +
	( 14'sd 7484) * $signed(input_fmap_123[15:0]) +
	( 16'sd 16428) * $signed(input_fmap_124[15:0]) +
	( 16'sd 27882) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6288) * $signed(input_fmap_126[15:0]) +
	( 14'sd 6452) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 16'sd 19391) * $signed(input_fmap_0[15:0]) +
	( 14'sd 6131) * $signed(input_fmap_1[15:0]) +
	( 15'sd 8317) * $signed(input_fmap_2[15:0]) +
	( 16'sd 26494) * $signed(input_fmap_3[15:0]) +
	( 16'sd 28969) * $signed(input_fmap_4[15:0]) +
	( 15'sd 10448) * $signed(input_fmap_5[15:0]) +
	( 16'sd 22098) * $signed(input_fmap_6[15:0]) +
	( 12'sd 1237) * $signed(input_fmap_7[15:0]) +
	( 12'sd 1183) * $signed(input_fmap_8[15:0]) +
	( 15'sd 13037) * $signed(input_fmap_9[15:0]) +
	( 15'sd 9995) * $signed(input_fmap_10[15:0]) +
	( 16'sd 30794) * $signed(input_fmap_11[15:0]) +
	( 16'sd 31163) * $signed(input_fmap_12[15:0]) +
	( 15'sd 14775) * $signed(input_fmap_13[15:0]) +
	( 16'sd 21620) * $signed(input_fmap_14[15:0]) +
	( 14'sd 6690) * $signed(input_fmap_15[15:0]) +
	( 14'sd 5942) * $signed(input_fmap_16[15:0]) +
	( 14'sd 6789) * $signed(input_fmap_17[15:0]) +
	( 15'sd 15134) * $signed(input_fmap_18[15:0]) +
	( 16'sd 19022) * $signed(input_fmap_19[15:0]) +
	( 14'sd 4542) * $signed(input_fmap_20[15:0]) +
	( 14'sd 5718) * $signed(input_fmap_21[15:0]) +
	( 16'sd 21020) * $signed(input_fmap_22[15:0]) +
	( 16'sd 27148) * $signed(input_fmap_23[15:0]) +
	( 16'sd 20545) * $signed(input_fmap_24[15:0]) +
	( 15'sd 15129) * $signed(input_fmap_25[15:0]) +
	( 15'sd 15792) * $signed(input_fmap_26[15:0]) +
	( 14'sd 6002) * $signed(input_fmap_27[15:0]) +
	( 15'sd 10192) * $signed(input_fmap_28[15:0]) +
	( 14'sd 6135) * $signed(input_fmap_29[15:0]) +
	( 15'sd 13828) * $signed(input_fmap_30[15:0]) +
	( 10'sd 277) * $signed(input_fmap_31[15:0]) +
	( 15'sd 8693) * $signed(input_fmap_32[15:0]) +
	( 15'sd 14960) * $signed(input_fmap_33[15:0]) +
	( 16'sd 17915) * $signed(input_fmap_34[15:0]) +
	( 16'sd 27576) * $signed(input_fmap_35[15:0]) +
	( 16'sd 24459) * $signed(input_fmap_36[15:0]) +
	( 16'sd 18402) * $signed(input_fmap_37[15:0]) +
	( 15'sd 14775) * $signed(input_fmap_38[15:0]) +
	( 16'sd 18274) * $signed(input_fmap_39[15:0]) +
	( 14'sd 8101) * $signed(input_fmap_40[15:0]) +
	( 12'sd 1661) * $signed(input_fmap_41[15:0]) +
	( 14'sd 5166) * $signed(input_fmap_42[15:0]) +
	( 16'sd 19479) * $signed(input_fmap_43[15:0]) +
	( 14'sd 7765) * $signed(input_fmap_44[15:0]) +
	( 15'sd 8985) * $signed(input_fmap_45[15:0]) +
	( 16'sd 16845) * $signed(input_fmap_46[15:0]) +
	( 16'sd 26509) * $signed(input_fmap_47[15:0]) +
	( 16'sd 31786) * $signed(input_fmap_48[15:0]) +
	( 16'sd 21649) * $signed(input_fmap_49[15:0]) +
	( 16'sd 24676) * $signed(input_fmap_50[15:0]) +
	( 16'sd 28013) * $signed(input_fmap_51[15:0]) +
	( 14'sd 7698) * $signed(input_fmap_52[15:0]) +
	( 13'sd 2788) * $signed(input_fmap_53[15:0]) +
	( 14'sd 6874) * $signed(input_fmap_54[15:0]) +
	( 15'sd 8830) * $signed(input_fmap_55[15:0]) +
	( 16'sd 16901) * $signed(input_fmap_56[15:0]) +
	( 10'sd 485) * $signed(input_fmap_57[15:0]) +
	( 16'sd 21887) * $signed(input_fmap_58[15:0]) +
	( 15'sd 10851) * $signed(input_fmap_59[15:0]) +
	( 14'sd 5096) * $signed(input_fmap_60[15:0]) +
	( 16'sd 30675) * $signed(input_fmap_61[15:0]) +
	( 16'sd 18148) * $signed(input_fmap_62[15:0]) +
	( 16'sd 27030) * $signed(input_fmap_63[15:0]) +
	( 16'sd 16665) * $signed(input_fmap_64[15:0]) +
	( 16'sd 26976) * $signed(input_fmap_65[15:0]) +
	( 16'sd 20589) * $signed(input_fmap_66[15:0]) +
	( 16'sd 20868) * $signed(input_fmap_67[15:0]) +
	( 16'sd 22011) * $signed(input_fmap_68[15:0]) +
	( 16'sd 23687) * $signed(input_fmap_69[15:0]) +
	( 16'sd 22732) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11173) * $signed(input_fmap_71[15:0]) +
	( 16'sd 22888) * $signed(input_fmap_72[15:0]) +
	( 15'sd 9769) * $signed(input_fmap_73[15:0]) +
	( 16'sd 18264) * $signed(input_fmap_74[15:0]) +
	( 16'sd 25083) * $signed(input_fmap_75[15:0]) +
	( 16'sd 28960) * $signed(input_fmap_76[15:0]) +
	( 14'sd 8059) * $signed(input_fmap_77[15:0]) +
	( 15'sd 11978) * $signed(input_fmap_78[15:0]) +
	( 13'sd 3275) * $signed(input_fmap_79[15:0]) +
	( 16'sd 23294) * $signed(input_fmap_80[15:0]) +
	( 15'sd 11229) * $signed(input_fmap_81[15:0]) +
	( 16'sd 21958) * $signed(input_fmap_82[15:0]) +
	( 15'sd 10062) * $signed(input_fmap_83[15:0]) +
	( 16'sd 17937) * $signed(input_fmap_84[15:0]) +
	( 16'sd 21393) * $signed(input_fmap_85[15:0]) +
	( 16'sd 31226) * $signed(input_fmap_86[15:0]) +
	( 16'sd 18069) * $signed(input_fmap_87[15:0]) +
	( 16'sd 24460) * $signed(input_fmap_88[15:0]) +
	( 16'sd 25125) * $signed(input_fmap_89[15:0]) +
	( 13'sd 3703) * $signed(input_fmap_90[15:0]) +
	( 15'sd 14474) * $signed(input_fmap_91[15:0]) +
	( 16'sd 18371) * $signed(input_fmap_92[15:0]) +
	( 15'sd 10650) * $signed(input_fmap_93[15:0]) +
	( 16'sd 30069) * $signed(input_fmap_94[15:0]) +
	( 14'sd 4551) * $signed(input_fmap_95[15:0]) +
	( 14'sd 7944) * $signed(input_fmap_96[15:0]) +
	( 16'sd 16601) * $signed(input_fmap_97[15:0]) +
	( 16'sd 29321) * $signed(input_fmap_98[15:0]) +
	( 16'sd 31627) * $signed(input_fmap_99[15:0]) +
	( 15'sd 14684) * $signed(input_fmap_100[15:0]) +
	( 16'sd 29268) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5258) * $signed(input_fmap_102[15:0]) +
	( 15'sd 12179) * $signed(input_fmap_103[15:0]) +
	( 16'sd 30782) * $signed(input_fmap_104[15:0]) +
	( 13'sd 4072) * $signed(input_fmap_105[15:0]) +
	( 15'sd 14233) * $signed(input_fmap_106[15:0]) +
	( 16'sd 16710) * $signed(input_fmap_107[15:0]) +
	( 16'sd 27794) * $signed(input_fmap_108[15:0]) +
	( 14'sd 7385) * $signed(input_fmap_109[15:0]) +
	( 16'sd 27025) * $signed(input_fmap_110[15:0]) +
	( 14'sd 5860) * $signed(input_fmap_111[15:0]) +
	( 15'sd 10533) * $signed(input_fmap_112[15:0]) +
	( 13'sd 3192) * $signed(input_fmap_113[15:0]) +
	( 15'sd 15929) * $signed(input_fmap_114[15:0]) +
	( 16'sd 19622) * $signed(input_fmap_115[15:0]) +
	( 10'sd 486) * $signed(input_fmap_116[15:0]) +
	( 13'sd 3063) * $signed(input_fmap_117[15:0]) +
	( 15'sd 10235) * $signed(input_fmap_118[15:0]) +
	( 16'sd 30572) * $signed(input_fmap_119[15:0]) +
	( 15'sd 13404) * $signed(input_fmap_120[15:0]) +
	( 16'sd 29379) * $signed(input_fmap_121[15:0]) +
	( 16'sd 26127) * $signed(input_fmap_122[15:0]) +
	( 13'sd 2997) * $signed(input_fmap_123[15:0]) +
	( 16'sd 26475) * $signed(input_fmap_124[15:0]) +
	( 16'sd 31700) * $signed(input_fmap_125[15:0]) +
	( 16'sd 24269) * $signed(input_fmap_126[15:0]) +
	( 16'sd 17702) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 15'sd 13733) * $signed(input_fmap_0[15:0]) +
	( 16'sd 31029) * $signed(input_fmap_1[15:0]) +
	( 14'sd 4459) * $signed(input_fmap_2[15:0]) +
	( 15'sd 12506) * $signed(input_fmap_3[15:0]) +
	( 16'sd 18017) * $signed(input_fmap_4[15:0]) +
	( 13'sd 3949) * $signed(input_fmap_5[15:0]) +
	( 16'sd 27339) * $signed(input_fmap_6[15:0]) +
	( 14'sd 5769) * $signed(input_fmap_7[15:0]) +
	( 16'sd 22027) * $signed(input_fmap_8[15:0]) +
	( 16'sd 29850) * $signed(input_fmap_9[15:0]) +
	( 16'sd 22186) * $signed(input_fmap_10[15:0]) +
	( 16'sd 20093) * $signed(input_fmap_11[15:0]) +
	( 15'sd 9661) * $signed(input_fmap_12[15:0]) +
	( 15'sd 13247) * $signed(input_fmap_13[15:0]) +
	( 16'sd 25887) * $signed(input_fmap_14[15:0]) +
	( 15'sd 13547) * $signed(input_fmap_15[15:0]) +
	( 16'sd 26821) * $signed(input_fmap_16[15:0]) +
	( 16'sd 28556) * $signed(input_fmap_17[15:0]) +
	( 15'sd 8734) * $signed(input_fmap_18[15:0]) +
	( 15'sd 13646) * $signed(input_fmap_19[15:0]) +
	( 16'sd 25265) * $signed(input_fmap_20[15:0]) +
	( 16'sd 23839) * $signed(input_fmap_21[15:0]) +
	( 15'sd 8373) * $signed(input_fmap_22[15:0]) +
	( 15'sd 9811) * $signed(input_fmap_23[15:0]) +
	( 14'sd 5214) * $signed(input_fmap_24[15:0]) +
	( 16'sd 30982) * $signed(input_fmap_25[15:0]) +
	( 14'sd 7662) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1672) * $signed(input_fmap_27[15:0]) +
	( 16'sd 31308) * $signed(input_fmap_28[15:0]) +
	( 16'sd 24384) * $signed(input_fmap_29[15:0]) +
	( 15'sd 13907) * $signed(input_fmap_30[15:0]) +
	( 16'sd 25645) * $signed(input_fmap_31[15:0]) +
	( 16'sd 19535) * $signed(input_fmap_32[15:0]) +
	( 12'sd 1123) * $signed(input_fmap_33[15:0]) +
	( 15'sd 13738) * $signed(input_fmap_34[15:0]) +
	( 16'sd 25543) * $signed(input_fmap_35[15:0]) +
	( 16'sd 28211) * $signed(input_fmap_36[15:0]) +
	( 16'sd 32695) * $signed(input_fmap_37[15:0]) +
	( 16'sd 31887) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24975) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6585) * $signed(input_fmap_40[15:0]) +
	( 14'sd 5725) * $signed(input_fmap_41[15:0]) +
	( 16'sd 16852) * $signed(input_fmap_42[15:0]) +
	( 16'sd 30035) * $signed(input_fmap_43[15:0]) +
	( 16'sd 17329) * $signed(input_fmap_44[15:0]) +
	( 16'sd 16947) * $signed(input_fmap_45[15:0]) +
	( 12'sd 1846) * $signed(input_fmap_46[15:0]) +
	( 11'sd 700) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13799) * $signed(input_fmap_48[15:0]) +
	( 16'sd 31221) * $signed(input_fmap_49[15:0]) +
	( 15'sd 11218) * $signed(input_fmap_50[15:0]) +
	( 15'sd 8591) * $signed(input_fmap_51[15:0]) +
	( 15'sd 9396) * $signed(input_fmap_52[15:0]) +
	( 16'sd 18297) * $signed(input_fmap_53[15:0]) +
	( 16'sd 21616) * $signed(input_fmap_54[15:0]) +
	( 15'sd 15586) * $signed(input_fmap_55[15:0]) +
	( 16'sd 25381) * $signed(input_fmap_56[15:0]) +
	( 16'sd 27301) * $signed(input_fmap_57[15:0]) +
	( 16'sd 30030) * $signed(input_fmap_58[15:0]) +
	( 15'sd 12385) * $signed(input_fmap_59[15:0]) +
	( 16'sd 25562) * $signed(input_fmap_60[15:0]) +
	( 15'sd 8695) * $signed(input_fmap_61[15:0]) +
	( 15'sd 13299) * $signed(input_fmap_62[15:0]) +
	( 16'sd 29299) * $signed(input_fmap_63[15:0]) +
	( 15'sd 9555) * $signed(input_fmap_64[15:0]) +
	( 15'sd 15910) * $signed(input_fmap_65[15:0]) +
	( 16'sd 18889) * $signed(input_fmap_66[15:0]) +
	( 11'sd 573) * $signed(input_fmap_67[15:0]) +
	( 15'sd 13281) * $signed(input_fmap_68[15:0]) +
	( 15'sd 10598) * $signed(input_fmap_69[15:0]) +
	( 15'sd 13659) * $signed(input_fmap_70[15:0]) +
	( 16'sd 27730) * $signed(input_fmap_71[15:0]) +
	( 13'sd 3669) * $signed(input_fmap_72[15:0]) +
	( 15'sd 9638) * $signed(input_fmap_73[15:0]) +
	( 16'sd 32459) * $signed(input_fmap_74[15:0]) +
	( 16'sd 23361) * $signed(input_fmap_75[15:0]) +
	( 16'sd 18505) * $signed(input_fmap_76[15:0]) +
	( 14'sd 6500) * $signed(input_fmap_77[15:0]) +
	( 15'sd 13760) * $signed(input_fmap_78[15:0]) +
	( 14'sd 7538) * $signed(input_fmap_79[15:0]) +
	( 14'sd 6555) * $signed(input_fmap_80[15:0]) +
	( 15'sd 9512) * $signed(input_fmap_81[15:0]) +
	( 16'sd 18440) * $signed(input_fmap_82[15:0]) +
	( 16'sd 29851) * $signed(input_fmap_83[15:0]) +
	( 16'sd 27681) * $signed(input_fmap_84[15:0]) +
	( 15'sd 16142) * $signed(input_fmap_85[15:0]) +
	( 16'sd 25949) * $signed(input_fmap_86[15:0]) +
	( 16'sd 16878) * $signed(input_fmap_87[15:0]) +
	( 13'sd 3276) * $signed(input_fmap_88[15:0]) +
	( 16'sd 30267) * $signed(input_fmap_89[15:0]) +
	( 16'sd 23225) * $signed(input_fmap_90[15:0]) +
	( 16'sd 30716) * $signed(input_fmap_91[15:0]) +
	( 12'sd 1991) * $signed(input_fmap_92[15:0]) +
	( 14'sd 7243) * $signed(input_fmap_93[15:0]) +
	( 14'sd 4747) * $signed(input_fmap_94[15:0]) +
	( 16'sd 22107) * $signed(input_fmap_95[15:0]) +
	( 16'sd 19802) * $signed(input_fmap_96[15:0]) +
	( 16'sd 20913) * $signed(input_fmap_97[15:0]) +
	( 14'sd 7266) * $signed(input_fmap_98[15:0]) +
	( 16'sd 19581) * $signed(input_fmap_99[15:0]) +
	( 15'sd 15710) * $signed(input_fmap_100[15:0]) +
	( 16'sd 23924) * $signed(input_fmap_101[15:0]) +
	( 16'sd 21757) * $signed(input_fmap_102[15:0]) +
	( 16'sd 29307) * $signed(input_fmap_103[15:0]) +
	( 16'sd 25947) * $signed(input_fmap_104[15:0]) +
	( 16'sd 23275) * $signed(input_fmap_105[15:0]) +
	( 15'sd 10295) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27135) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15769) * $signed(input_fmap_108[15:0]) +
	( 16'sd 16449) * $signed(input_fmap_109[15:0]) +
	( 16'sd 17615) * $signed(input_fmap_110[15:0]) +
	( 15'sd 8657) * $signed(input_fmap_111[15:0]) +
	( 12'sd 1564) * $signed(input_fmap_112[15:0]) +
	( 16'sd 21247) * $signed(input_fmap_113[15:0]) +
	( 16'sd 18420) * $signed(input_fmap_114[15:0]) +
	( 15'sd 8875) * $signed(input_fmap_115[15:0]) +
	( 16'sd 17069) * $signed(input_fmap_116[15:0]) +
	( 16'sd 18725) * $signed(input_fmap_117[15:0]) +
	( 16'sd 26071) * $signed(input_fmap_118[15:0]) +
	( 16'sd 25479) * $signed(input_fmap_119[15:0]) +
	( 15'sd 15330) * $signed(input_fmap_120[15:0]) +
	( 14'sd 6191) * $signed(input_fmap_121[15:0]) +
	( 11'sd 602) * $signed(input_fmap_122[15:0]) +
	( 16'sd 26026) * $signed(input_fmap_123[15:0]) +
	( 16'sd 18834) * $signed(input_fmap_124[15:0]) +
	( 11'sd 605) * $signed(input_fmap_125[15:0]) +
	( 16'sd 26970) * $signed(input_fmap_126[15:0]) +
	( 14'sd 7037) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 15'sd 13664) * $signed(input_fmap_0[15:0]) +
	( 16'sd 28847) * $signed(input_fmap_1[15:0]) +
	( 16'sd 27434) * $signed(input_fmap_2[15:0]) +
	( 15'sd 15644) * $signed(input_fmap_3[15:0]) +
	( 16'sd 18376) * $signed(input_fmap_4[15:0]) +
	( 11'sd 513) * $signed(input_fmap_5[15:0]) +
	( 15'sd 14827) * $signed(input_fmap_6[15:0]) +
	( 15'sd 10987) * $signed(input_fmap_7[15:0]) +
	( 16'sd 26419) * $signed(input_fmap_8[15:0]) +
	( 15'sd 8961) * $signed(input_fmap_9[15:0]) +
	( 12'sd 1203) * $signed(input_fmap_10[15:0]) +
	( 16'sd 23056) * $signed(input_fmap_11[15:0]) +
	( 16'sd 25417) * $signed(input_fmap_12[15:0]) +
	( 15'sd 10636) * $signed(input_fmap_13[15:0]) +
	( 15'sd 12871) * $signed(input_fmap_14[15:0]) +
	( 12'sd 1904) * $signed(input_fmap_15[15:0]) +
	( 16'sd 24284) * $signed(input_fmap_16[15:0]) +
	( 15'sd 12765) * $signed(input_fmap_17[15:0]) +
	( 15'sd 12332) * $signed(input_fmap_18[15:0]) +
	( 15'sd 9520) * $signed(input_fmap_19[15:0]) +
	( 16'sd 25914) * $signed(input_fmap_20[15:0]) +
	( 16'sd 18867) * $signed(input_fmap_21[15:0]) +
	( 14'sd 5717) * $signed(input_fmap_22[15:0]) +
	( 13'sd 3031) * $signed(input_fmap_23[15:0]) +
	( 13'sd 3048) * $signed(input_fmap_24[15:0]) +
	( 13'sd 3344) * $signed(input_fmap_25[15:0]) +
	( 16'sd 25594) * $signed(input_fmap_26[15:0]) +
	( 15'sd 15228) * $signed(input_fmap_27[15:0]) +
	( 13'sd 3899) * $signed(input_fmap_28[15:0]) +
	( 16'sd 24247) * $signed(input_fmap_29[15:0]) +
	( 14'sd 5829) * $signed(input_fmap_30[15:0]) +
	( 15'sd 8657) * $signed(input_fmap_31[15:0]) +
	( 16'sd 27455) * $signed(input_fmap_32[15:0]) +
	( 16'sd 24838) * $signed(input_fmap_33[15:0]) +
	( 16'sd 30478) * $signed(input_fmap_34[15:0]) +
	( 16'sd 19243) * $signed(input_fmap_35[15:0]) +
	( 16'sd 16786) * $signed(input_fmap_36[15:0]) +
	( 16'sd 17839) * $signed(input_fmap_37[15:0]) +
	( 13'sd 2893) * $signed(input_fmap_38[15:0]) +
	( 15'sd 15570) * $signed(input_fmap_39[15:0]) +
	( 15'sd 15748) * $signed(input_fmap_40[15:0]) +
	( 12'sd 1120) * $signed(input_fmap_41[15:0]) +
	( 16'sd 25165) * $signed(input_fmap_42[15:0]) +
	( 16'sd 30439) * $signed(input_fmap_43[15:0]) +
	( 16'sd 27681) * $signed(input_fmap_44[15:0]) +
	( 16'sd 17604) * $signed(input_fmap_45[15:0]) +
	( 10'sd 463) * $signed(input_fmap_46[15:0]) +
	( 16'sd 18860) * $signed(input_fmap_47[15:0]) +
	( 16'sd 25292) * $signed(input_fmap_48[15:0]) +
	( 16'sd 20348) * $signed(input_fmap_49[15:0]) +
	( 16'sd 20326) * $signed(input_fmap_50[15:0]) +
	( 16'sd 28108) * $signed(input_fmap_51[15:0]) +
	( 15'sd 13882) * $signed(input_fmap_52[15:0]) +
	( 15'sd 15697) * $signed(input_fmap_53[15:0]) +
	( 16'sd 23577) * $signed(input_fmap_54[15:0]) +
	( 15'sd 8236) * $signed(input_fmap_55[15:0]) +
	( 16'sd 19571) * $signed(input_fmap_56[15:0]) +
	( 13'sd 2375) * $signed(input_fmap_57[15:0]) +
	( 16'sd 23687) * $signed(input_fmap_58[15:0]) +
	( 16'sd 26773) * $signed(input_fmap_59[15:0]) +
	( 16'sd 18747) * $signed(input_fmap_60[15:0]) +
	( 16'sd 32386) * $signed(input_fmap_61[15:0]) +
	( 15'sd 11388) * $signed(input_fmap_62[15:0]) +
	( 14'sd 4784) * $signed(input_fmap_63[15:0]) +
	( 16'sd 22185) * $signed(input_fmap_64[15:0]) +
	( 16'sd 16930) * $signed(input_fmap_65[15:0]) +
	( 16'sd 28286) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28219) * $signed(input_fmap_67[15:0]) +
	( 14'sd 6409) * $signed(input_fmap_68[15:0]) +
	( 16'sd 29634) * $signed(input_fmap_69[15:0]) +
	( 16'sd 23539) * $signed(input_fmap_70[15:0]) +
	( 16'sd 20947) * $signed(input_fmap_71[15:0]) +
	( 16'sd 22439) * $signed(input_fmap_72[15:0]) +
	( 15'sd 12658) * $signed(input_fmap_73[15:0]) +
	( 15'sd 14071) * $signed(input_fmap_74[15:0]) +
	( 14'sd 4104) * $signed(input_fmap_75[15:0]) +
	( 16'sd 18637) * $signed(input_fmap_76[15:0]) +
	( 16'sd 18242) * $signed(input_fmap_77[15:0]) +
	( 15'sd 13241) * $signed(input_fmap_78[15:0]) +
	( 15'sd 12675) * $signed(input_fmap_79[15:0]) +
	( 16'sd 21341) * $signed(input_fmap_80[15:0]) +
	( 13'sd 2777) * $signed(input_fmap_81[15:0]) +
	( 16'sd 31192) * $signed(input_fmap_82[15:0]) +
	( 15'sd 10296) * $signed(input_fmap_83[15:0]) +
	( 16'sd 21183) * $signed(input_fmap_84[15:0]) +
	( 16'sd 32089) * $signed(input_fmap_85[15:0]) +
	( 16'sd 19772) * $signed(input_fmap_86[15:0]) +
	( 9'sd 188) * $signed(input_fmap_87[15:0]) +
	( 16'sd 23479) * $signed(input_fmap_88[15:0]) +
	( 16'sd 23221) * $signed(input_fmap_89[15:0]) +
	( 16'sd 24353) * $signed(input_fmap_90[15:0]) +
	( 16'sd 18127) * $signed(input_fmap_91[15:0]) +
	( 16'sd 20233) * $signed(input_fmap_92[15:0]) +
	( 16'sd 27153) * $signed(input_fmap_93[15:0]) +
	( 16'sd 18345) * $signed(input_fmap_94[15:0]) +
	( 16'sd 19527) * $signed(input_fmap_95[15:0]) +
	( 16'sd 24662) * $signed(input_fmap_96[15:0]) +
	( 16'sd 32167) * $signed(input_fmap_97[15:0]) +
	( 15'sd 9685) * $signed(input_fmap_98[15:0]) +
	( 16'sd 29424) * $signed(input_fmap_99[15:0]) +
	( 16'sd 19842) * $signed(input_fmap_100[15:0]) +
	( 13'sd 4057) * $signed(input_fmap_101[15:0]) +
	( 16'sd 23899) * $signed(input_fmap_102[15:0]) +
	( 16'sd 32345) * $signed(input_fmap_103[15:0]) +
	( 14'sd 4917) * $signed(input_fmap_104[15:0]) +
	( 16'sd 20701) * $signed(input_fmap_105[15:0]) +
	( 14'sd 7705) * $signed(input_fmap_106[15:0]) +
	( 16'sd 29393) * $signed(input_fmap_107[15:0]) +
	( 16'sd 24935) * $signed(input_fmap_108[15:0]) +
	( 16'sd 31591) * $signed(input_fmap_109[15:0]) +
	( 16'sd 17771) * $signed(input_fmap_110[15:0]) +
	( 16'sd 23301) * $signed(input_fmap_111[15:0]) +
	( 16'sd 17547) * $signed(input_fmap_112[15:0]) +
	( 12'sd 1851) * $signed(input_fmap_113[15:0]) +
	( 16'sd 24296) * $signed(input_fmap_114[15:0]) +
	( 16'sd 25687) * $signed(input_fmap_115[15:0]) +
	( 16'sd 17037) * $signed(input_fmap_116[15:0]) +
	( 15'sd 15735) * $signed(input_fmap_117[15:0]) +
	( 14'sd 7109) * $signed(input_fmap_118[15:0]) +
	( 15'sd 15755) * $signed(input_fmap_119[15:0]) +
	( 16'sd 24542) * $signed(input_fmap_120[15:0]) +
	( 15'sd 10084) * $signed(input_fmap_121[15:0]) +
	( 10'sd 281) * $signed(input_fmap_122[15:0]) +
	( 16'sd 23668) * $signed(input_fmap_123[15:0]) +
	( 14'sd 5115) * $signed(input_fmap_124[15:0]) +
	( 15'sd 14222) * $signed(input_fmap_125[15:0]) +
	( 14'sd 5404) * $signed(input_fmap_126[15:0]) +
	( 13'sd 3897) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 16'sd 27132) * $signed(input_fmap_0[15:0]) +
	( 16'sd 27690) * $signed(input_fmap_1[15:0]) +
	( 15'sd 13596) * $signed(input_fmap_2[15:0]) +
	( 15'sd 12861) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30244) * $signed(input_fmap_4[15:0]) +
	( 15'sd 11609) * $signed(input_fmap_5[15:0]) +
	( 13'sd 3861) * $signed(input_fmap_6[15:0]) +
	( 15'sd 11278) * $signed(input_fmap_7[15:0]) +
	( 16'sd 27816) * $signed(input_fmap_8[15:0]) +
	( 16'sd 19698) * $signed(input_fmap_9[15:0]) +
	( 16'sd 31643) * $signed(input_fmap_10[15:0]) +
	( 16'sd 17977) * $signed(input_fmap_11[15:0]) +
	( 16'sd 21966) * $signed(input_fmap_12[15:0]) +
	( 16'sd 21951) * $signed(input_fmap_13[15:0]) +
	( 16'sd 22564) * $signed(input_fmap_14[15:0]) +
	( 15'sd 15563) * $signed(input_fmap_15[15:0]) +
	( 15'sd 16203) * $signed(input_fmap_16[15:0]) +
	( 15'sd 10712) * $signed(input_fmap_17[15:0]) +
	( 16'sd 27038) * $signed(input_fmap_18[15:0]) +
	( 16'sd 20851) * $signed(input_fmap_19[15:0]) +
	( 16'sd 23135) * $signed(input_fmap_20[15:0]) +
	( 15'sd 12034) * $signed(input_fmap_21[15:0]) +
	( 16'sd 24904) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28359) * $signed(input_fmap_23[15:0]) +
	( 15'sd 15070) * $signed(input_fmap_24[15:0]) +
	( 14'sd 7979) * $signed(input_fmap_25[15:0]) +
	( 14'sd 6053) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1142) * $signed(input_fmap_27[15:0]) +
	( 16'sd 19837) * $signed(input_fmap_28[15:0]) +
	( 16'sd 32653) * $signed(input_fmap_29[15:0]) +
	( 16'sd 17253) * $signed(input_fmap_30[15:0]) +
	( 15'sd 8933) * $signed(input_fmap_31[15:0]) +
	( 16'sd 19321) * $signed(input_fmap_32[15:0]) +
	( 16'sd 32175) * $signed(input_fmap_33[15:0]) +
	( 16'sd 22784) * $signed(input_fmap_34[15:0]) +
	( 13'sd 3464) * $signed(input_fmap_35[15:0]) +
	( 16'sd 27158) * $signed(input_fmap_36[15:0]) +
	( 16'sd 29764) * $signed(input_fmap_37[15:0]) +
	( 16'sd 18888) * $signed(input_fmap_38[15:0]) +
	( 14'sd 6423) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6795) * $signed(input_fmap_40[15:0]) +
	( 15'sd 14557) * $signed(input_fmap_41[15:0]) +
	( 15'sd 8759) * $signed(input_fmap_42[15:0]) +
	( 13'sd 4067) * $signed(input_fmap_43[15:0]) +
	( 16'sd 32286) * $signed(input_fmap_44[15:0]) +
	( 16'sd 20690) * $signed(input_fmap_45[15:0]) +
	( 14'sd 6723) * $signed(input_fmap_46[15:0]) +
	( 16'sd 16567) * $signed(input_fmap_47[15:0]) +
	( 16'sd 24147) * $signed(input_fmap_48[15:0]) +
	( 16'sd 20955) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22289) * $signed(input_fmap_50[15:0]) +
	( 11'sd 661) * $signed(input_fmap_51[15:0]) +
	( 16'sd 25407) * $signed(input_fmap_52[15:0]) +
	( 16'sd 26266) * $signed(input_fmap_53[15:0]) +
	( 10'sd 316) * $signed(input_fmap_54[15:0]) +
	( 16'sd 22905) * $signed(input_fmap_55[15:0]) +
	( 16'sd 31850) * $signed(input_fmap_56[15:0]) +
	( 12'sd 1487) * $signed(input_fmap_57[15:0]) +
	( 14'sd 4400) * $signed(input_fmap_58[15:0]) +
	( 16'sd 23508) * $signed(input_fmap_59[15:0]) +
	( 14'sd 5834) * $signed(input_fmap_60[15:0]) +
	( 16'sd 26331) * $signed(input_fmap_61[15:0]) +
	( 16'sd 17884) * $signed(input_fmap_62[15:0]) +
	( 14'sd 7799) * $signed(input_fmap_63[15:0]) +
	( 15'sd 10513) * $signed(input_fmap_64[15:0]) +
	( 16'sd 23365) * $signed(input_fmap_65[15:0]) +
	( 16'sd 20488) * $signed(input_fmap_66[15:0]) +
	( 14'sd 5964) * $signed(input_fmap_67[15:0]) +
	( 16'sd 21370) * $signed(input_fmap_68[15:0]) +
	( 15'sd 13575) * $signed(input_fmap_69[15:0]) +
	( 14'sd 6843) * $signed(input_fmap_70[15:0]) +
	( 15'sd 9333) * $signed(input_fmap_71[15:0]) +
	( 15'sd 15739) * $signed(input_fmap_72[15:0]) +
	( 15'sd 11590) * $signed(input_fmap_73[15:0]) +
	( 16'sd 19880) * $signed(input_fmap_74[15:0]) +
	( 16'sd 24260) * $signed(input_fmap_75[15:0]) +
	( 16'sd 25028) * $signed(input_fmap_76[15:0]) +
	( 14'sd 4324) * $signed(input_fmap_77[15:0]) +
	( 15'sd 15363) * $signed(input_fmap_78[15:0]) +
	( 16'sd 18441) * $signed(input_fmap_79[15:0]) +
	( 16'sd 31847) * $signed(input_fmap_80[15:0]) +
	( 14'sd 4238) * $signed(input_fmap_81[15:0]) +
	( 13'sd 3275) * $signed(input_fmap_82[15:0]) +
	( 15'sd 13720) * $signed(input_fmap_83[15:0]) +
	( 15'sd 9127) * $signed(input_fmap_84[15:0]) +
	( 16'sd 22551) * $signed(input_fmap_85[15:0]) +
	( 16'sd 30998) * $signed(input_fmap_86[15:0]) +
	( 15'sd 11060) * $signed(input_fmap_87[15:0]) +
	( 15'sd 9823) * $signed(input_fmap_88[15:0]) +
	( 15'sd 10180) * $signed(input_fmap_89[15:0]) +
	( 16'sd 22689) * $signed(input_fmap_90[15:0]) +
	( 16'sd 22871) * $signed(input_fmap_91[15:0]) +
	( 16'sd 19639) * $signed(input_fmap_92[15:0]) +
	( 16'sd 30595) * $signed(input_fmap_93[15:0]) +
	( 16'sd 27004) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25945) * $signed(input_fmap_95[15:0]) +
	( 15'sd 14225) * $signed(input_fmap_96[15:0]) +
	( 16'sd 19099) * $signed(input_fmap_97[15:0]) +
	( 14'sd 4295) * $signed(input_fmap_98[15:0]) +
	( 16'sd 22221) * $signed(input_fmap_99[15:0]) +
	( 16'sd 18516) * $signed(input_fmap_100[15:0]) +
	( 16'sd 27101) * $signed(input_fmap_101[15:0]) +
	( 16'sd 26949) * $signed(input_fmap_102[15:0]) +
	( 16'sd 20802) * $signed(input_fmap_103[15:0]) +
	( 14'sd 4732) * $signed(input_fmap_104[15:0]) +
	( 15'sd 14154) * $signed(input_fmap_105[15:0]) +
	( 16'sd 27220) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27767) * $signed(input_fmap_107[15:0]) +
	( 15'sd 14467) * $signed(input_fmap_108[15:0]) +
	( 15'sd 9929) * $signed(input_fmap_109[15:0]) +
	( 16'sd 30822) * $signed(input_fmap_110[15:0]) +
	( 15'sd 12262) * $signed(input_fmap_111[15:0]) +
	( 13'sd 3910) * $signed(input_fmap_112[15:0]) +
	( 13'sd 3476) * $signed(input_fmap_113[15:0]) +
	( 15'sd 11532) * $signed(input_fmap_114[15:0]) +
	( 16'sd 22307) * $signed(input_fmap_115[15:0]) +
	( 16'sd 24460) * $signed(input_fmap_116[15:0]) +
	( 15'sd 14393) * $signed(input_fmap_117[15:0]) +
	( 15'sd 10554) * $signed(input_fmap_118[15:0]) +
	( 16'sd 28240) * $signed(input_fmap_119[15:0]) +
	( 15'sd 10961) * $signed(input_fmap_120[15:0]) +
	( 16'sd 27115) * $signed(input_fmap_121[15:0]) +
	( 16'sd 32176) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21293) * $signed(input_fmap_123[15:0]) +
	( 15'sd 16356) * $signed(input_fmap_124[15:0]) +
	( 16'sd 26403) * $signed(input_fmap_125[15:0]) +
	( 16'sd 19497) * $signed(input_fmap_126[15:0]) +
	( 15'sd 15635) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 16'sd 20568) * $signed(input_fmap_0[15:0]) +
	( 15'sd 12009) * $signed(input_fmap_1[15:0]) +
	( 15'sd 8983) * $signed(input_fmap_2[15:0]) +
	( 15'sd 10876) * $signed(input_fmap_3[15:0]) +
	( 15'sd 8268) * $signed(input_fmap_4[15:0]) +
	( 16'sd 28248) * $signed(input_fmap_5[15:0]) +
	( 16'sd 30808) * $signed(input_fmap_6[15:0]) +
	( 15'sd 11813) * $signed(input_fmap_7[15:0]) +
	( 12'sd 1065) * $signed(input_fmap_8[15:0]) +
	( 13'sd 2192) * $signed(input_fmap_9[15:0]) +
	( 14'sd 5900) * $signed(input_fmap_10[15:0]) +
	( 15'sd 13669) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20773) * $signed(input_fmap_12[15:0]) +
	( 16'sd 29287) * $signed(input_fmap_13[15:0]) +
	( 14'sd 4965) * $signed(input_fmap_14[15:0]) +
	( 16'sd 21179) * $signed(input_fmap_15[15:0]) +
	( 15'sd 9935) * $signed(input_fmap_16[15:0]) +
	( 15'sd 9832) * $signed(input_fmap_17[15:0]) +
	( 14'sd 7147) * $signed(input_fmap_18[15:0]) +
	( 15'sd 11959) * $signed(input_fmap_19[15:0]) +
	( 16'sd 32580) * $signed(input_fmap_20[15:0]) +
	( 14'sd 8162) * $signed(input_fmap_21[15:0]) +
	( 16'sd 31292) * $signed(input_fmap_22[15:0]) +
	( 16'sd 31430) * $signed(input_fmap_23[15:0]) +
	( 11'sd 867) * $signed(input_fmap_24[15:0]) +
	( 16'sd 21858) * $signed(input_fmap_25[15:0]) +
	( 16'sd 32307) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2657) * $signed(input_fmap_27[15:0]) +
	( 16'sd 23730) * $signed(input_fmap_28[15:0]) +
	( 12'sd 1607) * $signed(input_fmap_29[15:0]) +
	( 16'sd 18374) * $signed(input_fmap_30[15:0]) +
	( 16'sd 17898) * $signed(input_fmap_31[15:0]) +
	( 15'sd 8715) * $signed(input_fmap_32[15:0]) +
	( 16'sd 18175) * $signed(input_fmap_33[15:0]) +
	( 16'sd 26684) * $signed(input_fmap_34[15:0]) +
	( 16'sd 17624) * $signed(input_fmap_35[15:0]) +
	( 16'sd 18895) * $signed(input_fmap_36[15:0]) +
	( 14'sd 6003) * $signed(input_fmap_37[15:0]) +
	( 16'sd 28575) * $signed(input_fmap_38[15:0]) +
	( 14'sd 7306) * $signed(input_fmap_39[15:0]) +
	( 10'sd 356) * $signed(input_fmap_40[15:0]) +
	( 13'sd 3185) * $signed(input_fmap_41[15:0]) +
	( 16'sd 21650) * $signed(input_fmap_42[15:0]) +
	( 14'sd 7187) * $signed(input_fmap_43[15:0]) +
	( 12'sd 1548) * $signed(input_fmap_44[15:0]) +
	( 16'sd 32498) * $signed(input_fmap_45[15:0]) +
	( 16'sd 24412) * $signed(input_fmap_46[15:0]) +
	( 16'sd 17251) * $signed(input_fmap_47[15:0]) +
	( 16'sd 28095) * $signed(input_fmap_48[15:0]) +
	( 16'sd 20885) * $signed(input_fmap_49[15:0]) +
	( 16'sd 28573) * $signed(input_fmap_50[15:0]) +
	( 16'sd 21398) * $signed(input_fmap_51[15:0]) +
	( 11'sd 954) * $signed(input_fmap_52[15:0]) +
	( 16'sd 21045) * $signed(input_fmap_53[15:0]) +
	( 15'sd 15042) * $signed(input_fmap_54[15:0]) +
	( 16'sd 18185) * $signed(input_fmap_55[15:0]) +
	( 15'sd 13720) * $signed(input_fmap_56[15:0]) +
	( 16'sd 16713) * $signed(input_fmap_57[15:0]) +
	( 16'sd 21514) * $signed(input_fmap_58[15:0]) +
	( 16'sd 27719) * $signed(input_fmap_59[15:0]) +
	( 16'sd 18845) * $signed(input_fmap_60[15:0]) +
	( 16'sd 22715) * $signed(input_fmap_61[15:0]) +
	( 15'sd 15870) * $signed(input_fmap_62[15:0]) +
	( 15'sd 10799) * $signed(input_fmap_63[15:0]) +
	( 14'sd 7755) * $signed(input_fmap_64[15:0]) +
	( 16'sd 20041) * $signed(input_fmap_65[15:0]) +
	( 13'sd 3534) * $signed(input_fmap_66[15:0]) +
	( 16'sd 29136) * $signed(input_fmap_67[15:0]) +
	( 13'sd 2195) * $signed(input_fmap_68[15:0]) +
	( 16'sd 23997) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31634) * $signed(input_fmap_70[15:0]) +
	( 15'sd 10231) * $signed(input_fmap_71[15:0]) +
	( 13'sd 2792) * $signed(input_fmap_72[15:0]) +
	( 16'sd 29208) * $signed(input_fmap_73[15:0]) +
	( 15'sd 13947) * $signed(input_fmap_74[15:0]) +
	( 15'sd 12156) * $signed(input_fmap_75[15:0]) +
	( 14'sd 7100) * $signed(input_fmap_76[15:0]) +
	( 16'sd 18129) * $signed(input_fmap_77[15:0]) +
	( 15'sd 12206) * $signed(input_fmap_78[15:0]) +
	( 16'sd 23324) * $signed(input_fmap_79[15:0]) +
	( 16'sd 17611) * $signed(input_fmap_80[15:0]) +
	( 16'sd 20000) * $signed(input_fmap_81[15:0]) +
	( 16'sd 28583) * $signed(input_fmap_82[15:0]) +
	( 16'sd 26741) * $signed(input_fmap_83[15:0]) +
	( 15'sd 11622) * $signed(input_fmap_84[15:0]) +
	( 14'sd 6179) * $signed(input_fmap_85[15:0]) +
	( 15'sd 13961) * $signed(input_fmap_86[15:0]) +
	( 16'sd 19750) * $signed(input_fmap_87[15:0]) +
	( 16'sd 22796) * $signed(input_fmap_88[15:0]) +
	( 15'sd 15189) * $signed(input_fmap_89[15:0]) +
	( 15'sd 12853) * $signed(input_fmap_90[15:0]) +
	( 10'sd 335) * $signed(input_fmap_91[15:0]) +
	( 16'sd 21720) * $signed(input_fmap_92[15:0]) +
	( 13'sd 2891) * $signed(input_fmap_93[15:0]) +
	( 15'sd 13023) * $signed(input_fmap_94[15:0]) +
	( 16'sd 16505) * $signed(input_fmap_95[15:0]) +
	( 15'sd 13093) * $signed(input_fmap_96[15:0]) +
	( 15'sd 8592) * $signed(input_fmap_97[15:0]) +
	( 16'sd 23877) * $signed(input_fmap_98[15:0]) +
	( 15'sd 11027) * $signed(input_fmap_99[15:0]) +
	( 16'sd 27058) * $signed(input_fmap_100[15:0]) +
	( 14'sd 5265) * $signed(input_fmap_101[15:0]) +
	( 14'sd 4901) * $signed(input_fmap_102[15:0]) +
	( 16'sd 30411) * $signed(input_fmap_103[15:0]) +
	( 15'sd 10159) * $signed(input_fmap_104[15:0]) +
	( 15'sd 11429) * $signed(input_fmap_105[15:0]) +
	( 15'sd 9484) * $signed(input_fmap_106[15:0]) +
	( 7'sd 38) * $signed(input_fmap_107[15:0]) +
	( 16'sd 26369) * $signed(input_fmap_108[15:0]) +
	( 13'sd 2877) * $signed(input_fmap_109[15:0]) +
	( 16'sd 21828) * $signed(input_fmap_110[15:0]) +
	( 14'sd 4733) * $signed(input_fmap_111[15:0]) +
	( 16'sd 16952) * $signed(input_fmap_112[15:0]) +
	( 16'sd 26852) * $signed(input_fmap_113[15:0]) +
	( 16'sd 29542) * $signed(input_fmap_114[15:0]) +
	( 7'sd 46) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26553) * $signed(input_fmap_116[15:0]) +
	( 14'sd 4723) * $signed(input_fmap_117[15:0]) +
	( 13'sd 2617) * $signed(input_fmap_118[15:0]) +
	( 9'sd 212) * $signed(input_fmap_119[15:0]) +
	( 15'sd 9197) * $signed(input_fmap_120[15:0]) +
	( 16'sd 27081) * $signed(input_fmap_121[15:0]) +
	( 16'sd 22706) * $signed(input_fmap_122[15:0]) +
	( 14'sd 6376) * $signed(input_fmap_123[15:0]) +
	( 13'sd 3781) * $signed(input_fmap_124[15:0]) +
	( 13'sd 3914) * $signed(input_fmap_125[15:0]) +
	( 15'sd 11640) * $signed(input_fmap_126[15:0]) +
	( 16'sd 25690) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 14'sd 7149) * $signed(input_fmap_0[15:0]) +
	( 15'sd 12578) * $signed(input_fmap_1[15:0]) +
	( 16'sd 25061) * $signed(input_fmap_2[15:0]) +
	( 12'sd 1870) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30536) * $signed(input_fmap_4[15:0]) +
	( 16'sd 23823) * $signed(input_fmap_5[15:0]) +
	( 16'sd 23965) * $signed(input_fmap_6[15:0]) +
	( 16'sd 22420) * $signed(input_fmap_7[15:0]) +
	( 16'sd 29759) * $signed(input_fmap_8[15:0]) +
	( 15'sd 12195) * $signed(input_fmap_9[15:0]) +
	( 14'sd 6499) * $signed(input_fmap_10[15:0]) +
	( 15'sd 12658) * $signed(input_fmap_11[15:0]) +
	( 15'sd 13956) * $signed(input_fmap_12[15:0]) +
	( 12'sd 1705) * $signed(input_fmap_13[15:0]) +
	( 14'sd 6666) * $signed(input_fmap_14[15:0]) +
	( 16'sd 18383) * $signed(input_fmap_15[15:0]) +
	( 16'sd 31121) * $signed(input_fmap_16[15:0]) +
	( 12'sd 1158) * $signed(input_fmap_17[15:0]) +
	( 15'sd 15948) * $signed(input_fmap_18[15:0]) +
	( 12'sd 1657) * $signed(input_fmap_19[15:0]) +
	( 14'sd 5880) * $signed(input_fmap_20[15:0]) +
	( 14'sd 7779) * $signed(input_fmap_21[15:0]) +
	( 14'sd 4553) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28386) * $signed(input_fmap_23[15:0]) +
	( 16'sd 18582) * $signed(input_fmap_24[15:0]) +
	( 15'sd 9400) * $signed(input_fmap_25[15:0]) +
	( 16'sd 23387) * $signed(input_fmap_26[15:0]) +
	( 15'sd 15955) * $signed(input_fmap_27[15:0]) +
	( 15'sd 10654) * $signed(input_fmap_28[15:0]) +
	( 12'sd 1331) * $signed(input_fmap_29[15:0]) +
	( 16'sd 28520) * $signed(input_fmap_30[15:0]) +
	( 10'sd 508) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28323) * $signed(input_fmap_32[15:0]) +
	( 16'sd 23475) * $signed(input_fmap_33[15:0]) +
	( 15'sd 9542) * $signed(input_fmap_34[15:0]) +
	( 16'sd 31142) * $signed(input_fmap_35[15:0]) +
	( 14'sd 5086) * $signed(input_fmap_36[15:0]) +
	( 15'sd 8525) * $signed(input_fmap_37[15:0]) +
	( 11'sd 603) * $signed(input_fmap_38[15:0]) +
	( 12'sd 1570) * $signed(input_fmap_39[15:0]) +
	( 16'sd 19175) * $signed(input_fmap_40[15:0]) +
	( 16'sd 22502) * $signed(input_fmap_41[15:0]) +
	( 15'sd 16159) * $signed(input_fmap_42[15:0]) +
	( 16'sd 19062) * $signed(input_fmap_43[15:0]) +
	( 16'sd 17844) * $signed(input_fmap_44[15:0]) +
	( 16'sd 25901) * $signed(input_fmap_45[15:0]) +
	( 15'sd 10863) * $signed(input_fmap_46[15:0]) +
	( 16'sd 24456) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13721) * $signed(input_fmap_48[15:0]) +
	( 16'sd 18323) * $signed(input_fmap_49[15:0]) +
	( 14'sd 4652) * $signed(input_fmap_50[15:0]) +
	( 16'sd 25081) * $signed(input_fmap_51[15:0]) +
	( 16'sd 30036) * $signed(input_fmap_52[15:0]) +
	( 14'sd 5206) * $signed(input_fmap_53[15:0]) +
	( 15'sd 14736) * $signed(input_fmap_54[15:0]) +
	( 13'sd 2741) * $signed(input_fmap_55[15:0]) +
	( 16'sd 18685) * $signed(input_fmap_56[15:0]) +
	( 15'sd 11509) * $signed(input_fmap_57[15:0]) +
	( 11'sd 933) * $signed(input_fmap_58[15:0]) +
	( 11'sd 984) * $signed(input_fmap_59[15:0]) +
	( 16'sd 24262) * $signed(input_fmap_60[15:0]) +
	( 13'sd 4062) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29995) * $signed(input_fmap_62[15:0]) +
	( 14'sd 7484) * $signed(input_fmap_63[15:0]) +
	( 16'sd 27829) * $signed(input_fmap_64[15:0]) +
	( 16'sd 26960) * $signed(input_fmap_65[15:0]) +
	( 15'sd 10560) * $signed(input_fmap_66[15:0]) +
	( 14'sd 8047) * $signed(input_fmap_67[15:0]) +
	( 16'sd 16849) * $signed(input_fmap_68[15:0]) +
	( 14'sd 5339) * $signed(input_fmap_69[15:0]) +
	( 16'sd 20970) * $signed(input_fmap_70[15:0]) +
	( 16'sd 22270) * $signed(input_fmap_71[15:0]) +
	( 14'sd 4937) * $signed(input_fmap_72[15:0]) +
	( 10'sd 367) * $signed(input_fmap_73[15:0]) +
	( 16'sd 22728) * $signed(input_fmap_74[15:0]) +
	( 14'sd 7339) * $signed(input_fmap_75[15:0]) +
	( 16'sd 26339) * $signed(input_fmap_76[15:0]) +
	( 16'sd 17268) * $signed(input_fmap_77[15:0]) +
	( 16'sd 30549) * $signed(input_fmap_78[15:0]) +
	( 16'sd 27895) * $signed(input_fmap_79[15:0]) +
	( 14'sd 5153) * $signed(input_fmap_80[15:0]) +
	( 16'sd 31462) * $signed(input_fmap_81[15:0]) +
	( 16'sd 27787) * $signed(input_fmap_82[15:0]) +
	( 16'sd 26826) * $signed(input_fmap_83[15:0]) +
	( 16'sd 23528) * $signed(input_fmap_84[15:0]) +
	( 15'sd 12742) * $signed(input_fmap_85[15:0]) +
	( 14'sd 5743) * $signed(input_fmap_86[15:0]) +
	( 16'sd 20874) * $signed(input_fmap_87[15:0]) +
	( 16'sd 18117) * $signed(input_fmap_88[15:0]) +
	( 16'sd 17982) * $signed(input_fmap_89[15:0]) +
	( 16'sd 24132) * $signed(input_fmap_90[15:0]) +
	( 15'sd 12687) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25860) * $signed(input_fmap_92[15:0]) +
	( 16'sd 19860) * $signed(input_fmap_93[15:0]) +
	( 12'sd 1938) * $signed(input_fmap_94[15:0]) +
	( 16'sd 16779) * $signed(input_fmap_95[15:0]) +
	( 16'sd 25153) * $signed(input_fmap_96[15:0]) +
	( 15'sd 13772) * $signed(input_fmap_97[15:0]) +
	( 15'sd 15886) * $signed(input_fmap_98[15:0]) +
	( 16'sd 17840) * $signed(input_fmap_99[15:0]) +
	( 10'sd 452) * $signed(input_fmap_100[15:0]) +
	( 16'sd 26793) * $signed(input_fmap_101[15:0]) +
	( 16'sd 20778) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28847) * $signed(input_fmap_103[15:0]) +
	( 16'sd 23533) * $signed(input_fmap_104[15:0]) +
	( 16'sd 22178) * $signed(input_fmap_105[15:0]) +
	( 15'sd 12933) * $signed(input_fmap_106[15:0]) +
	( 16'sd 28342) * $signed(input_fmap_107[15:0]) +
	( 14'sd 6861) * $signed(input_fmap_108[15:0]) +
	( 14'sd 5099) * $signed(input_fmap_109[15:0]) +
	( 16'sd 17165) * $signed(input_fmap_110[15:0]) +
	( 16'sd 20420) * $signed(input_fmap_111[15:0]) +
	( 16'sd 28549) * $signed(input_fmap_112[15:0]) +
	( 15'sd 15028) * $signed(input_fmap_113[15:0]) +
	( 16'sd 30467) * $signed(input_fmap_114[15:0]) +
	( 16'sd 17133) * $signed(input_fmap_115[15:0]) +
	( 14'sd 4864) * $signed(input_fmap_116[15:0]) +
	( 13'sd 2969) * $signed(input_fmap_117[15:0]) +
	( 13'sd 2529) * $signed(input_fmap_118[15:0]) +
	( 15'sd 10705) * $signed(input_fmap_119[15:0]) +
	( 16'sd 25248) * $signed(input_fmap_120[15:0]) +
	( 16'sd 30414) * $signed(input_fmap_121[15:0]) +
	( 11'sd 557) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21654) * $signed(input_fmap_123[15:0]) +
	( 16'sd 30502) * $signed(input_fmap_124[15:0]) +
	( 14'sd 6162) * $signed(input_fmap_125[15:0]) +
	( 13'sd 3679) * $signed(input_fmap_126[15:0]) +
	( 15'sd 8765) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 13'sd 2853) * $signed(input_fmap_0[15:0]) +
	( 16'sd 32662) * $signed(input_fmap_1[15:0]) +
	( 16'sd 17624) * $signed(input_fmap_2[15:0]) +
	( 14'sd 5850) * $signed(input_fmap_3[15:0]) +
	( 14'sd 4881) * $signed(input_fmap_4[15:0]) +
	( 15'sd 13481) * $signed(input_fmap_5[15:0]) +
	( 12'sd 1224) * $signed(input_fmap_6[15:0]) +
	( 15'sd 10309) * $signed(input_fmap_7[15:0]) +
	( 16'sd 18532) * $signed(input_fmap_8[15:0]) +
	( 15'sd 15911) * $signed(input_fmap_9[15:0]) +
	( 15'sd 10000) * $signed(input_fmap_10[15:0]) +
	( 15'sd 9640) * $signed(input_fmap_11[15:0]) +
	( 16'sd 28919) * $signed(input_fmap_12[15:0]) +
	( 16'sd 19097) * $signed(input_fmap_13[15:0]) +
	( 14'sd 6185) * $signed(input_fmap_14[15:0]) +
	( 16'sd 24280) * $signed(input_fmap_15[15:0]) +
	( 16'sd 30402) * $signed(input_fmap_16[15:0]) +
	( 13'sd 2499) * $signed(input_fmap_17[15:0]) +
	( 16'sd 18498) * $signed(input_fmap_18[15:0]) +
	( 15'sd 13295) * $signed(input_fmap_19[15:0]) +
	( 14'sd 6093) * $signed(input_fmap_20[15:0]) +
	( 16'sd 20968) * $signed(input_fmap_21[15:0]) +
	( 16'sd 30053) * $signed(input_fmap_22[15:0]) +
	( 15'sd 15985) * $signed(input_fmap_23[15:0]) +
	( 16'sd 18966) * $signed(input_fmap_24[15:0]) +
	( 16'sd 31329) * $signed(input_fmap_25[15:0]) +
	( 14'sd 6919) * $signed(input_fmap_26[15:0]) +
	( 16'sd 21079) * $signed(input_fmap_27[15:0]) +
	( 16'sd 23887) * $signed(input_fmap_28[15:0]) +
	( 16'sd 21999) * $signed(input_fmap_29[15:0]) +
	( 16'sd 20555) * $signed(input_fmap_30[15:0]) +
	( 14'sd 7230) * $signed(input_fmap_31[15:0]) +
	( 16'sd 23930) * $signed(input_fmap_32[15:0]) +
	( 14'sd 7100) * $signed(input_fmap_33[15:0]) +
	( 13'sd 2322) * $signed(input_fmap_34[15:0]) +
	( 15'sd 12849) * $signed(input_fmap_35[15:0]) +
	( 14'sd 4824) * $signed(input_fmap_36[15:0]) +
	( 15'sd 16230) * $signed(input_fmap_37[15:0]) +
	( 16'sd 17393) * $signed(input_fmap_38[15:0]) +
	( 15'sd 14730) * $signed(input_fmap_39[15:0]) +
	( 15'sd 10167) * $signed(input_fmap_40[15:0]) +
	( 14'sd 4800) * $signed(input_fmap_41[15:0]) +
	( 15'sd 14931) * $signed(input_fmap_42[15:0]) +
	( 16'sd 25023) * $signed(input_fmap_43[15:0]) +
	( 16'sd 27301) * $signed(input_fmap_44[15:0]) +
	( 16'sd 32413) * $signed(input_fmap_45[15:0]) +
	( 16'sd 21926) * $signed(input_fmap_46[15:0]) +
	( 16'sd 16605) * $signed(input_fmap_47[15:0]) +
	( 16'sd 18721) * $signed(input_fmap_48[15:0]) +
	( 15'sd 13234) * $signed(input_fmap_49[15:0]) +
	( 16'sd 24673) * $signed(input_fmap_50[15:0]) +
	( 15'sd 11390) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3842) * $signed(input_fmap_52[15:0]) +
	( 16'sd 27128) * $signed(input_fmap_53[15:0]) +
	( 15'sd 11052) * $signed(input_fmap_54[15:0]) +
	( 15'sd 10383) * $signed(input_fmap_55[15:0]) +
	( 13'sd 3668) * $signed(input_fmap_56[15:0]) +
	( 16'sd 27177) * $signed(input_fmap_57[15:0]) +
	( 16'sd 24314) * $signed(input_fmap_58[15:0]) +
	( 15'sd 13510) * $signed(input_fmap_59[15:0]) +
	( 15'sd 15950) * $signed(input_fmap_60[15:0]) +
	( 14'sd 7560) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29151) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20670) * $signed(input_fmap_63[15:0]) +
	( 16'sd 30307) * $signed(input_fmap_64[15:0]) +
	( 16'sd 31695) * $signed(input_fmap_65[15:0]) +
	( 15'sd 9929) * $signed(input_fmap_66[15:0]) +
	( 16'sd 27884) * $signed(input_fmap_67[15:0]) +
	( 16'sd 20480) * $signed(input_fmap_68[15:0]) +
	( 13'sd 3640) * $signed(input_fmap_69[15:0]) +
	( 14'sd 7275) * $signed(input_fmap_70[15:0]) +
	( 16'sd 28728) * $signed(input_fmap_71[15:0]) +
	( 15'sd 10261) * $signed(input_fmap_72[15:0]) +
	( 14'sd 5908) * $signed(input_fmap_73[15:0]) +
	( 16'sd 17032) * $signed(input_fmap_74[15:0]) +
	( 10'sd 420) * $signed(input_fmap_75[15:0]) +
	( 16'sd 28343) * $signed(input_fmap_76[15:0]) +
	( 16'sd 32262) * $signed(input_fmap_77[15:0]) +
	( 11'sd 798) * $signed(input_fmap_78[15:0]) +
	( 16'sd 16825) * $signed(input_fmap_79[15:0]) +
	( 16'sd 32405) * $signed(input_fmap_80[15:0]) +
	( 15'sd 11295) * $signed(input_fmap_81[15:0]) +
	( 16'sd 18197) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25662) * $signed(input_fmap_83[15:0]) +
	( 16'sd 18376) * $signed(input_fmap_84[15:0]) +
	( 14'sd 5072) * $signed(input_fmap_85[15:0]) +
	( 15'sd 12775) * $signed(input_fmap_86[15:0]) +
	( 14'sd 4184) * $signed(input_fmap_87[15:0]) +
	( 16'sd 16796) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5297) * $signed(input_fmap_89[15:0]) +
	( 14'sd 4147) * $signed(input_fmap_90[15:0]) +
	( 16'sd 23297) * $signed(input_fmap_91[15:0]) +
	( 16'sd 26333) * $signed(input_fmap_92[15:0]) +
	( 14'sd 4659) * $signed(input_fmap_93[15:0]) +
	( 16'sd 19381) * $signed(input_fmap_94[15:0]) +
	( 16'sd 30322) * $signed(input_fmap_95[15:0]) +
	( 14'sd 4559) * $signed(input_fmap_96[15:0]) +
	( 14'sd 7833) * $signed(input_fmap_97[15:0]) +
	( 16'sd 22146) * $signed(input_fmap_98[15:0]) +
	( 15'sd 12280) * $signed(input_fmap_99[15:0]) +
	( 14'sd 8152) * $signed(input_fmap_100[15:0]) +
	( 15'sd 14723) * $signed(input_fmap_101[15:0]) +
	( 15'sd 9076) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28496) * $signed(input_fmap_103[15:0]) +
	( 16'sd 19343) * $signed(input_fmap_104[15:0]) +
	( 16'sd 26884) * $signed(input_fmap_105[15:0]) +
	( 13'sd 3560) * $signed(input_fmap_106[15:0]) +
	( 16'sd 19818) * $signed(input_fmap_107[15:0]) +
	( 14'sd 6210) * $signed(input_fmap_108[15:0]) +
	( 16'sd 29969) * $signed(input_fmap_109[15:0]) +
	( 16'sd 27140) * $signed(input_fmap_110[15:0]) +
	( 16'sd 22789) * $signed(input_fmap_111[15:0]) +
	( 14'sd 6589) * $signed(input_fmap_112[15:0]) +
	( 15'sd 10682) * $signed(input_fmap_113[15:0]) +
	( 13'sd 3775) * $signed(input_fmap_114[15:0]) +
	( 16'sd 20562) * $signed(input_fmap_115[15:0]) +
	( 16'sd 30241) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27233) * $signed(input_fmap_117[15:0]) +
	( 15'sd 13244) * $signed(input_fmap_118[15:0]) +
	( 16'sd 23081) * $signed(input_fmap_119[15:0]) +
	( 16'sd 23760) * $signed(input_fmap_120[15:0]) +
	( 16'sd 21136) * $signed(input_fmap_121[15:0]) +
	( 12'sd 1725) * $signed(input_fmap_122[15:0]) +
	( 16'sd 31735) * $signed(input_fmap_123[15:0]) +
	( 16'sd 28106) * $signed(input_fmap_124[15:0]) +
	( 16'sd 25349) * $signed(input_fmap_125[15:0]) +
	( 16'sd 23436) * $signed(input_fmap_126[15:0]) +
	( 16'sd 16630) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 16'sd 20779) * $signed(input_fmap_0[15:0]) +
	( 16'sd 30345) * $signed(input_fmap_1[15:0]) +
	( 15'sd 12086) * $signed(input_fmap_2[15:0]) +
	( 16'sd 26460) * $signed(input_fmap_3[15:0]) +
	( 16'sd 27255) * $signed(input_fmap_4[15:0]) +
	( 14'sd 7050) * $signed(input_fmap_5[15:0]) +
	( 15'sd 12167) * $signed(input_fmap_6[15:0]) +
	( 16'sd 18852) * $signed(input_fmap_7[15:0]) +
	( 13'sd 2155) * $signed(input_fmap_8[15:0]) +
	( 16'sd 22719) * $signed(input_fmap_9[15:0]) +
	( 16'sd 22478) * $signed(input_fmap_10[15:0]) +
	( 15'sd 10410) * $signed(input_fmap_11[15:0]) +
	( 14'sd 5426) * $signed(input_fmap_12[15:0]) +
	( 15'sd 16093) * $signed(input_fmap_13[15:0]) +
	( 16'sd 29719) * $signed(input_fmap_14[15:0]) +
	( 15'sd 11913) * $signed(input_fmap_15[15:0]) +
	( 16'sd 31272) * $signed(input_fmap_16[15:0]) +
	( 16'sd 30127) * $signed(input_fmap_17[15:0]) +
	( 16'sd 20898) * $signed(input_fmap_18[15:0]) +
	( 14'sd 4652) * $signed(input_fmap_19[15:0]) +
	( 16'sd 26922) * $signed(input_fmap_20[15:0]) +
	( 16'sd 18511) * $signed(input_fmap_21[15:0]) +
	( 16'sd 19001) * $signed(input_fmap_22[15:0]) +
	( 16'sd 19155) * $signed(input_fmap_23[15:0]) +
	( 12'sd 1398) * $signed(input_fmap_24[15:0]) +
	( 16'sd 22345) * $signed(input_fmap_25[15:0]) +
	( 16'sd 17864) * $signed(input_fmap_26[15:0]) +
	( 16'sd 18365) * $signed(input_fmap_27[15:0]) +
	( 15'sd 8738) * $signed(input_fmap_28[15:0]) +
	( 8'sd 84) * $signed(input_fmap_29[15:0]) +
	( 16'sd 26497) * $signed(input_fmap_30[15:0]) +
	( 15'sd 13340) * $signed(input_fmap_31[15:0]) +
	( 16'sd 17476) * $signed(input_fmap_32[15:0]) +
	( 14'sd 8099) * $signed(input_fmap_33[15:0]) +
	( 14'sd 5567) * $signed(input_fmap_34[15:0]) +
	( 15'sd 12792) * $signed(input_fmap_35[15:0]) +
	( 16'sd 26080) * $signed(input_fmap_36[15:0]) +
	( 11'sd 991) * $signed(input_fmap_37[15:0]) +
	( 16'sd 25930) * $signed(input_fmap_38[15:0]) +
	( 16'sd 18209) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6601) * $signed(input_fmap_40[15:0]) +
	( 13'sd 3127) * $signed(input_fmap_41[15:0]) +
	( 16'sd 18814) * $signed(input_fmap_42[15:0]) +
	( 13'sd 2593) * $signed(input_fmap_43[15:0]) +
	( 13'sd 3310) * $signed(input_fmap_44[15:0]) +
	( 16'sd 32431) * $signed(input_fmap_45[15:0]) +
	( 14'sd 4569) * $signed(input_fmap_46[15:0]) +
	( 12'sd 1601) * $signed(input_fmap_47[15:0]) +
	( 14'sd 6830) * $signed(input_fmap_48[15:0]) +
	( 16'sd 28836) * $signed(input_fmap_49[15:0]) +
	( 14'sd 4574) * $signed(input_fmap_50[15:0]) +
	( 16'sd 29067) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3791) * $signed(input_fmap_52[15:0]) +
	( 16'sd 18156) * $signed(input_fmap_53[15:0]) +
	( 12'sd 1113) * $signed(input_fmap_54[15:0]) +
	( 16'sd 22515) * $signed(input_fmap_55[15:0]) +
	( 16'sd 30640) * $signed(input_fmap_56[15:0]) +
	( 16'sd 27185) * $signed(input_fmap_57[15:0]) +
	( 16'sd 32038) * $signed(input_fmap_58[15:0]) +
	( 15'sd 12812) * $signed(input_fmap_59[15:0]) +
	( 15'sd 11262) * $signed(input_fmap_60[15:0]) +
	( 16'sd 26035) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3328) * $signed(input_fmap_62[15:0]) +
	( 14'sd 5150) * $signed(input_fmap_63[15:0]) +
	( 16'sd 26748) * $signed(input_fmap_64[15:0]) +
	( 12'sd 1646) * $signed(input_fmap_65[15:0]) +
	( 15'sd 13818) * $signed(input_fmap_66[15:0]) +
	( 15'sd 11838) * $signed(input_fmap_67[15:0]) +
	( 15'sd 10983) * $signed(input_fmap_68[15:0]) +
	( 14'sd 4618) * $signed(input_fmap_69[15:0]) +
	( 15'sd 11078) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31240) * $signed(input_fmap_71[15:0]) +
	( 15'sd 9194) * $signed(input_fmap_72[15:0]) +
	( 13'sd 2693) * $signed(input_fmap_73[15:0]) +
	( 11'sd 786) * $signed(input_fmap_74[15:0]) +
	( 15'sd 12167) * $signed(input_fmap_75[15:0]) +
	( 15'sd 10357) * $signed(input_fmap_76[15:0]) +
	( 16'sd 18557) * $signed(input_fmap_77[15:0]) +
	( 16'sd 27974) * $signed(input_fmap_78[15:0]) +
	( 16'sd 21889) * $signed(input_fmap_79[15:0]) +
	( 13'sd 3125) * $signed(input_fmap_80[15:0]) +
	( 16'sd 23691) * $signed(input_fmap_81[15:0]) +
	( 16'sd 17058) * $signed(input_fmap_82[15:0]) +
	( 15'sd 14792) * $signed(input_fmap_83[15:0]) +
	( 15'sd 13380) * $signed(input_fmap_84[15:0]) +
	( 15'sd 16135) * $signed(input_fmap_85[15:0]) +
	( 13'sd 2085) * $signed(input_fmap_86[15:0]) +
	( 14'sd 6645) * $signed(input_fmap_87[15:0]) +
	( 16'sd 24637) * $signed(input_fmap_88[15:0]) +
	( 15'sd 11262) * $signed(input_fmap_89[15:0]) +
	( 15'sd 10062) * $signed(input_fmap_90[15:0]) +
	( 16'sd 23024) * $signed(input_fmap_91[15:0]) +
	( 15'sd 13219) * $signed(input_fmap_92[15:0]) +
	( 16'sd 21780) * $signed(input_fmap_93[15:0]) +
	( 16'sd 30115) * $signed(input_fmap_94[15:0]) +
	( 16'sd 17960) * $signed(input_fmap_95[15:0]) +
	( 16'sd 21019) * $signed(input_fmap_96[15:0]) +
	( 14'sd 6853) * $signed(input_fmap_97[15:0]) +
	( 16'sd 30719) * $signed(input_fmap_98[15:0]) +
	( 16'sd 29667) * $signed(input_fmap_99[15:0]) +
	( 16'sd 21436) * $signed(input_fmap_100[15:0]) +
	( 12'sd 1548) * $signed(input_fmap_101[15:0]) +
	( 16'sd 17796) * $signed(input_fmap_102[15:0]) +
	( 13'sd 3372) * $signed(input_fmap_103[15:0]) +
	( 16'sd 19253) * $signed(input_fmap_104[15:0]) +
	( 16'sd 19194) * $signed(input_fmap_105[15:0]) +
	( 16'sd 29654) * $signed(input_fmap_106[15:0]) +
	( 16'sd 28942) * $signed(input_fmap_107[15:0]) +
	( 13'sd 3078) * $signed(input_fmap_108[15:0]) +
	( 16'sd 19875) * $signed(input_fmap_109[15:0]) +
	( 15'sd 10723) * $signed(input_fmap_110[15:0]) +
	( 14'sd 4894) * $signed(input_fmap_111[15:0]) +
	( 16'sd 30934) * $signed(input_fmap_112[15:0]) +
	( 16'sd 28990) * $signed(input_fmap_113[15:0]) +
	( 16'sd 18650) * $signed(input_fmap_114[15:0]) +
	( 14'sd 4801) * $signed(input_fmap_115[15:0]) +
	( 14'sd 7849) * $signed(input_fmap_116[15:0]) +
	( 13'sd 2053) * $signed(input_fmap_117[15:0]) +
	( 16'sd 28152) * $signed(input_fmap_118[15:0]) +
	( 15'sd 12942) * $signed(input_fmap_119[15:0]) +
	( 16'sd 21206) * $signed(input_fmap_120[15:0]) +
	( 15'sd 9656) * $signed(input_fmap_121[15:0]) +
	( 16'sd 22799) * $signed(input_fmap_122[15:0]) +
	( 16'sd 19669) * $signed(input_fmap_123[15:0]) +
	( 16'sd 29062) * $signed(input_fmap_124[15:0]) +
	( 16'sd 20174) * $signed(input_fmap_125[15:0]) +
	( 14'sd 7450) * $signed(input_fmap_126[15:0]) +
	( 15'sd 9237) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 15'sd 11902) * $signed(input_fmap_0[15:0]) +
	( 14'sd 4167) * $signed(input_fmap_1[15:0]) +
	( 16'sd 19798) * $signed(input_fmap_2[15:0]) +
	( 16'sd 26951) * $signed(input_fmap_3[15:0]) +
	( 14'sd 4434) * $signed(input_fmap_4[15:0]) +
	( 15'sd 12395) * $signed(input_fmap_5[15:0]) +
	( 16'sd 28780) * $signed(input_fmap_6[15:0]) +
	( 14'sd 6015) * $signed(input_fmap_7[15:0]) +
	( 14'sd 6460) * $signed(input_fmap_8[15:0]) +
	( 16'sd 21938) * $signed(input_fmap_9[15:0]) +
	( 16'sd 31626) * $signed(input_fmap_10[15:0]) +
	( 16'sd 23725) * $signed(input_fmap_11[15:0]) +
	( 16'sd 19245) * $signed(input_fmap_12[15:0]) +
	( 15'sd 11937) * $signed(input_fmap_13[15:0]) +
	( 16'sd 30661) * $signed(input_fmap_14[15:0]) +
	( 16'sd 17936) * $signed(input_fmap_15[15:0]) +
	( 16'sd 30594) * $signed(input_fmap_16[15:0]) +
	( 15'sd 11676) * $signed(input_fmap_17[15:0]) +
	( 15'sd 15784) * $signed(input_fmap_18[15:0]) +
	( 16'sd 24502) * $signed(input_fmap_19[15:0]) +
	( 14'sd 4250) * $signed(input_fmap_20[15:0]) +
	( 15'sd 14304) * $signed(input_fmap_21[15:0]) +
	( 16'sd 23019) * $signed(input_fmap_22[15:0]) +
	( 16'sd 26819) * $signed(input_fmap_23[15:0]) +
	( 15'sd 12103) * $signed(input_fmap_24[15:0]) +
	( 15'sd 11584) * $signed(input_fmap_25[15:0]) +
	( 16'sd 26533) * $signed(input_fmap_26[15:0]) +
	( 15'sd 12571) * $signed(input_fmap_27[15:0]) +
	( 15'sd 13192) * $signed(input_fmap_28[15:0]) +
	( 13'sd 2253) * $signed(input_fmap_29[15:0]) +
	( 16'sd 18451) * $signed(input_fmap_30[15:0]) +
	( 16'sd 22898) * $signed(input_fmap_31[15:0]) +
	( 15'sd 9836) * $signed(input_fmap_32[15:0]) +
	( 13'sd 3969) * $signed(input_fmap_33[15:0]) +
	( 14'sd 4301) * $signed(input_fmap_34[15:0]) +
	( 16'sd 26530) * $signed(input_fmap_35[15:0]) +
	( 15'sd 15397) * $signed(input_fmap_36[15:0]) +
	( 16'sd 19615) * $signed(input_fmap_37[15:0]) +
	( 16'sd 16463) * $signed(input_fmap_38[15:0]) +
	( 16'sd 17547) * $signed(input_fmap_39[15:0]) +
	( 14'sd 4331) * $signed(input_fmap_40[15:0]) +
	( 15'sd 14794) * $signed(input_fmap_41[15:0]) +
	( 16'sd 20787) * $signed(input_fmap_42[15:0]) +
	( 15'sd 14619) * $signed(input_fmap_43[15:0]) +
	( 14'sd 4134) * $signed(input_fmap_44[15:0]) +
	( 15'sd 10448) * $signed(input_fmap_45[15:0]) +
	( 16'sd 30062) * $signed(input_fmap_46[15:0]) +
	( 15'sd 15952) * $signed(input_fmap_47[15:0]) +
	( 14'sd 4165) * $signed(input_fmap_48[15:0]) +
	( 16'sd 25667) * $signed(input_fmap_49[15:0]) +
	( 15'sd 9269) * $signed(input_fmap_50[15:0]) +
	( 15'sd 13782) * $signed(input_fmap_51[15:0]) +
	( 15'sd 14184) * $signed(input_fmap_52[15:0]) +
	( 14'sd 7515) * $signed(input_fmap_53[15:0]) +
	( 15'sd 8493) * $signed(input_fmap_54[15:0]) +
	( 16'sd 31490) * $signed(input_fmap_55[15:0]) +
	( 16'sd 31400) * $signed(input_fmap_56[15:0]) +
	( 14'sd 4259) * $signed(input_fmap_57[15:0]) +
	( 12'sd 1557) * $signed(input_fmap_58[15:0]) +
	( 15'sd 9082) * $signed(input_fmap_59[15:0]) +
	( 13'sd 2976) * $signed(input_fmap_60[15:0]) +
	( 15'sd 15851) * $signed(input_fmap_61[15:0]) +
	( 16'sd 31800) * $signed(input_fmap_62[15:0]) +
	( 16'sd 25207) * $signed(input_fmap_63[15:0]) +
	( 15'sd 15308) * $signed(input_fmap_64[15:0]) +
	( 14'sd 5150) * $signed(input_fmap_65[15:0]) +
	( 15'sd 12473) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28481) * $signed(input_fmap_67[15:0]) +
	( 14'sd 5428) * $signed(input_fmap_68[15:0]) +
	( 13'sd 2696) * $signed(input_fmap_69[15:0]) +
	( 16'sd 30915) * $signed(input_fmap_70[15:0]) +
	( 13'sd 2560) * $signed(input_fmap_71[15:0]) +
	( 16'sd 29536) * $signed(input_fmap_72[15:0]) +
	( 15'sd 9647) * $signed(input_fmap_73[15:0]) +
	( 14'sd 7884) * $signed(input_fmap_74[15:0]) +
	( 16'sd 27163) * $signed(input_fmap_75[15:0]) +
	( 14'sd 7246) * $signed(input_fmap_76[15:0]) +
	( 16'sd 24415) * $signed(input_fmap_77[15:0]) +
	( 14'sd 5071) * $signed(input_fmap_78[15:0]) +
	( 13'sd 3442) * $signed(input_fmap_79[15:0]) +
	( 15'sd 13126) * $signed(input_fmap_80[15:0]) +
	( 16'sd 24745) * $signed(input_fmap_81[15:0]) +
	( 16'sd 26699) * $signed(input_fmap_82[15:0]) +
	( 15'sd 13596) * $signed(input_fmap_83[15:0]) +
	( 15'sd 12839) * $signed(input_fmap_84[15:0]) +
	( 16'sd 23647) * $signed(input_fmap_85[15:0]) +
	( 15'sd 9497) * $signed(input_fmap_86[15:0]) +
	( 16'sd 20402) * $signed(input_fmap_87[15:0]) +
	( 16'sd 16629) * $signed(input_fmap_88[15:0]) +
	( 15'sd 15793) * $signed(input_fmap_89[15:0]) +
	( 15'sd 8827) * $signed(input_fmap_90[15:0]) +
	( 12'sd 1139) * $signed(input_fmap_91[15:0]) +
	( 16'sd 29860) * $signed(input_fmap_92[15:0]) +
	( 16'sd 30699) * $signed(input_fmap_93[15:0]) +
	( 15'sd 14005) * $signed(input_fmap_94[15:0]) +
	( 16'sd 28215) * $signed(input_fmap_95[15:0]) +
	( 16'sd 31775) * $signed(input_fmap_96[15:0]) +
	( 15'sd 9387) * $signed(input_fmap_97[15:0]) +
	( 16'sd 27858) * $signed(input_fmap_98[15:0]) +
	( 16'sd 17326) * $signed(input_fmap_99[15:0]) +
	( 15'sd 13180) * $signed(input_fmap_100[15:0]) +
	( 14'sd 6854) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5938) * $signed(input_fmap_102[15:0]) +
	( 10'sd 469) * $signed(input_fmap_103[15:0]) +
	( 16'sd 21358) * $signed(input_fmap_104[15:0]) +
	( 16'sd 21416) * $signed(input_fmap_105[15:0]) +
	( 16'sd 20874) * $signed(input_fmap_106[15:0]) +
	( 16'sd 16410) * $signed(input_fmap_107[15:0]) +
	( 16'sd 24355) * $signed(input_fmap_108[15:0]) +
	( 14'sd 5753) * $signed(input_fmap_109[15:0]) +
	( 16'sd 26163) * $signed(input_fmap_110[15:0]) +
	( 16'sd 20864) * $signed(input_fmap_111[15:0]) +
	( 15'sd 15145) * $signed(input_fmap_112[15:0]) +
	( 16'sd 28749) * $signed(input_fmap_113[15:0]) +
	( 16'sd 30820) * $signed(input_fmap_114[15:0]) +
	( 15'sd 16177) * $signed(input_fmap_115[15:0]) +
	( 16'sd 18374) * $signed(input_fmap_116[15:0]) +
	( 14'sd 6385) * $signed(input_fmap_117[15:0]) +
	( 16'sd 16753) * $signed(input_fmap_118[15:0]) +
	( 15'sd 14075) * $signed(input_fmap_119[15:0]) +
	( 15'sd 8880) * $signed(input_fmap_120[15:0]) +
	( 13'sd 3147) * $signed(input_fmap_121[15:0]) +
	( 16'sd 17224) * $signed(input_fmap_122[15:0]) +
	( 15'sd 11377) * $signed(input_fmap_123[15:0]) +
	( 14'sd 4931) * $signed(input_fmap_124[15:0]) +
	( 15'sd 14387) * $signed(input_fmap_125[15:0]) +
	( 16'sd 27665) * $signed(input_fmap_126[15:0]) +
	( 16'sd 27359) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 13'sd 2770) * $signed(input_fmap_0[15:0]) +
	( 16'sd 26257) * $signed(input_fmap_1[15:0]) +
	( 15'sd 10713) * $signed(input_fmap_2[15:0]) +
	( 16'sd 24587) * $signed(input_fmap_3[15:0]) +
	( 13'sd 3078) * $signed(input_fmap_4[15:0]) +
	( 16'sd 23946) * $signed(input_fmap_5[15:0]) +
	( 16'sd 25793) * $signed(input_fmap_6[15:0]) +
	( 16'sd 18676) * $signed(input_fmap_7[15:0]) +
	( 16'sd 32353) * $signed(input_fmap_8[15:0]) +
	( 14'sd 6227) * $signed(input_fmap_9[15:0]) +
	( 16'sd 21657) * $signed(input_fmap_10[15:0]) +
	( 16'sd 17860) * $signed(input_fmap_11[15:0]) +
	( 13'sd 4031) * $signed(input_fmap_12[15:0]) +
	( 14'sd 7467) * $signed(input_fmap_13[15:0]) +
	( 16'sd 25028) * $signed(input_fmap_14[15:0]) +
	( 10'sd 494) * $signed(input_fmap_15[15:0]) +
	( 16'sd 17128) * $signed(input_fmap_16[15:0]) +
	( 15'sd 16013) * $signed(input_fmap_17[15:0]) +
	( 15'sd 16309) * $signed(input_fmap_18[15:0]) +
	( 16'sd 31514) * $signed(input_fmap_19[15:0]) +
	( 16'sd 21493) * $signed(input_fmap_20[15:0]) +
	( 16'sd 28332) * $signed(input_fmap_21[15:0]) +
	( 15'sd 12628) * $signed(input_fmap_22[15:0]) +
	( 16'sd 18235) * $signed(input_fmap_23[15:0]) +
	( 16'sd 31049) * $signed(input_fmap_24[15:0]) +
	( 15'sd 13849) * $signed(input_fmap_25[15:0]) +
	( 16'sd 29476) * $signed(input_fmap_26[15:0]) +
	( 15'sd 16302) * $signed(input_fmap_27[15:0]) +
	( 13'sd 2949) * $signed(input_fmap_28[15:0]) +
	( 16'sd 25416) * $signed(input_fmap_29[15:0]) +
	( 16'sd 23458) * $signed(input_fmap_30[15:0]) +
	( 16'sd 28930) * $signed(input_fmap_31[15:0]) +
	( 14'sd 6995) * $signed(input_fmap_32[15:0]) +
	( 15'sd 16180) * $signed(input_fmap_33[15:0]) +
	( 15'sd 13237) * $signed(input_fmap_34[15:0]) +
	( 15'sd 10907) * $signed(input_fmap_35[15:0]) +
	( 15'sd 14529) * $signed(input_fmap_36[15:0]) +
	( 13'sd 3311) * $signed(input_fmap_37[15:0]) +
	( 16'sd 29496) * $signed(input_fmap_38[15:0]) +
	( 16'sd 22807) * $signed(input_fmap_39[15:0]) +
	( 16'sd 16665) * $signed(input_fmap_40[15:0]) +
	( 15'sd 9842) * $signed(input_fmap_41[15:0]) +
	( 14'sd 6453) * $signed(input_fmap_42[15:0]) +
	( 16'sd 20894) * $signed(input_fmap_43[15:0]) +
	( 15'sd 8715) * $signed(input_fmap_44[15:0]) +
	( 16'sd 23855) * $signed(input_fmap_45[15:0]) +
	( 16'sd 28509) * $signed(input_fmap_46[15:0]) +
	( 15'sd 12525) * $signed(input_fmap_47[15:0]) +
	( 16'sd 29042) * $signed(input_fmap_48[15:0]) +
	( 16'sd 28880) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26833) * $signed(input_fmap_50[15:0]) +
	( 15'sd 16128) * $signed(input_fmap_51[15:0]) +
	( 16'sd 17222) * $signed(input_fmap_52[15:0]) +
	( 16'sd 32616) * $signed(input_fmap_53[15:0]) +
	( 15'sd 8502) * $signed(input_fmap_54[15:0]) +
	( 15'sd 15760) * $signed(input_fmap_55[15:0]) +
	( 16'sd 18634) * $signed(input_fmap_56[15:0]) +
	( 15'sd 16368) * $signed(input_fmap_57[15:0]) +
	( 13'sd 2605) * $signed(input_fmap_58[15:0]) +
	( 10'sd 443) * $signed(input_fmap_59[15:0]) +
	( 14'sd 5596) * $signed(input_fmap_60[15:0]) +
	( 15'sd 15382) * $signed(input_fmap_61[15:0]) +
	( 15'sd 13298) * $signed(input_fmap_62[15:0]) +
	( 15'sd 12143) * $signed(input_fmap_63[15:0]) +
	( 15'sd 13266) * $signed(input_fmap_64[15:0]) +
	( 14'sd 6228) * $signed(input_fmap_65[15:0]) +
	( 10'sd 410) * $signed(input_fmap_66[15:0]) +
	( 16'sd 29925) * $signed(input_fmap_67[15:0]) +
	( 16'sd 31870) * $signed(input_fmap_68[15:0]) +
	( 15'sd 9531) * $signed(input_fmap_69[15:0]) +
	( 12'sd 1209) * $signed(input_fmap_70[15:0]) +
	( 16'sd 28813) * $signed(input_fmap_71[15:0]) +
	( 16'sd 32197) * $signed(input_fmap_72[15:0]) +
	( 16'sd 28554) * $signed(input_fmap_73[15:0]) +
	( 16'sd 28508) * $signed(input_fmap_74[15:0]) +
	( 12'sd 1589) * $signed(input_fmap_75[15:0]) +
	( 16'sd 22396) * $signed(input_fmap_76[15:0]) +
	( 16'sd 25441) * $signed(input_fmap_77[15:0]) +
	( 16'sd 22084) * $signed(input_fmap_78[15:0]) +
	( 16'sd 23162) * $signed(input_fmap_79[15:0]) +
	( 15'sd 11084) * $signed(input_fmap_80[15:0]) +
	( 13'sd 3043) * $signed(input_fmap_81[15:0]) +
	( 15'sd 10182) * $signed(input_fmap_82[15:0]) +
	( 15'sd 15520) * $signed(input_fmap_83[15:0]) +
	( 16'sd 19263) * $signed(input_fmap_84[15:0]) +
	( 14'sd 5032) * $signed(input_fmap_85[15:0]) +
	( 16'sd 18782) * $signed(input_fmap_86[15:0]) +
	( 16'sd 16827) * $signed(input_fmap_87[15:0]) +
	( 13'sd 3775) * $signed(input_fmap_88[15:0]) +
	( 15'sd 13703) * $signed(input_fmap_89[15:0]) +
	( 16'sd 25272) * $signed(input_fmap_90[15:0]) +
	( 16'sd 29193) * $signed(input_fmap_91[15:0]) +
	( 16'sd 26333) * $signed(input_fmap_92[15:0]) +
	( 16'sd 23029) * $signed(input_fmap_93[15:0]) +
	( 11'sd 851) * $signed(input_fmap_94[15:0]) +
	( 15'sd 14065) * $signed(input_fmap_95[15:0]) +
	( 15'sd 13435) * $signed(input_fmap_96[15:0]) +
	( 15'sd 9030) * $signed(input_fmap_97[15:0]) +
	( 11'sd 880) * $signed(input_fmap_98[15:0]) +
	( 16'sd 26618) * $signed(input_fmap_99[15:0]) +
	( 14'sd 5350) * $signed(input_fmap_100[15:0]) +
	( 15'sd 12963) * $signed(input_fmap_101[15:0]) +
	( 16'sd 18407) * $signed(input_fmap_102[15:0]) +
	( 15'sd 9963) * $signed(input_fmap_103[15:0]) +
	( 16'sd 20329) * $signed(input_fmap_104[15:0]) +
	( 16'sd 17241) * $signed(input_fmap_105[15:0]) +
	( 16'sd 22664) * $signed(input_fmap_106[15:0]) +
	( 16'sd 25388) * $signed(input_fmap_107[15:0]) +
	( 16'sd 16519) * $signed(input_fmap_108[15:0]) +
	( 16'sd 21371) * $signed(input_fmap_109[15:0]) +
	( 16'sd 17613) * $signed(input_fmap_110[15:0]) +
	( 16'sd 26142) * $signed(input_fmap_111[15:0]) +
	( 15'sd 10626) * $signed(input_fmap_112[15:0]) +
	( 14'sd 5529) * $signed(input_fmap_113[15:0]) +
	( 16'sd 22234) * $signed(input_fmap_114[15:0]) +
	( 16'sd 24890) * $signed(input_fmap_115[15:0]) +
	( 16'sd 18469) * $signed(input_fmap_116[15:0]) +
	( 15'sd 9922) * $signed(input_fmap_117[15:0]) +
	( 15'sd 9984) * $signed(input_fmap_118[15:0]) +
	( 12'sd 1824) * $signed(input_fmap_119[15:0]) +
	( 16'sd 32717) * $signed(input_fmap_120[15:0]) +
	( 16'sd 18670) * $signed(input_fmap_121[15:0]) +
	( 16'sd 20935) * $signed(input_fmap_122[15:0]) +
	( 16'sd 30544) * $signed(input_fmap_123[15:0]) +
	( 15'sd 13603) * $signed(input_fmap_124[15:0]) +
	( 15'sd 13588) * $signed(input_fmap_125[15:0]) +
	( 16'sd 18608) * $signed(input_fmap_126[15:0]) +
	( 15'sd 12651) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 16'sd 22721) * $signed(input_fmap_0[15:0]) +
	( 13'sd 3336) * $signed(input_fmap_1[15:0]) +
	( 16'sd 28833) * $signed(input_fmap_2[15:0]) +
	( 14'sd 6610) * $signed(input_fmap_3[15:0]) +
	( 16'sd 20768) * $signed(input_fmap_4[15:0]) +
	( 16'sd 21456) * $signed(input_fmap_5[15:0]) +
	( 16'sd 21108) * $signed(input_fmap_6[15:0]) +
	( 13'sd 2050) * $signed(input_fmap_7[15:0]) +
	( 16'sd 16913) * $signed(input_fmap_8[15:0]) +
	( 14'sd 6646) * $signed(input_fmap_9[15:0]) +
	( 10'sd 401) * $signed(input_fmap_10[15:0]) +
	( 16'sd 26966) * $signed(input_fmap_11[15:0]) +
	( 15'sd 12088) * $signed(input_fmap_12[15:0]) +
	( 16'sd 23126) * $signed(input_fmap_13[15:0]) +
	( 14'sd 6687) * $signed(input_fmap_14[15:0]) +
	( 14'sd 7178) * $signed(input_fmap_15[15:0]) +
	( 13'sd 3767) * $signed(input_fmap_16[15:0]) +
	( 11'sd 684) * $signed(input_fmap_17[15:0]) +
	( 16'sd 32427) * $signed(input_fmap_18[15:0]) +
	( 16'sd 22127) * $signed(input_fmap_19[15:0]) +
	( 14'sd 5225) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17306) * $signed(input_fmap_21[15:0]) +
	( 16'sd 27450) * $signed(input_fmap_22[15:0]) +
	( 14'sd 6120) * $signed(input_fmap_23[15:0]) +
	( 15'sd 16274) * $signed(input_fmap_24[15:0]) +
	( 16'sd 32704) * $signed(input_fmap_25[15:0]) +
	( 16'sd 21170) * $signed(input_fmap_26[15:0]) +
	( 15'sd 10876) * $signed(input_fmap_27[15:0]) +
	( 16'sd 28627) * $signed(input_fmap_28[15:0]) +
	( 16'sd 27658) * $signed(input_fmap_29[15:0]) +
	( 10'sd 426) * $signed(input_fmap_30[15:0]) +
	( 14'sd 8128) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28613) * $signed(input_fmap_32[15:0]) +
	( 16'sd 22340) * $signed(input_fmap_33[15:0]) +
	( 13'sd 2806) * $signed(input_fmap_34[15:0]) +
	( 16'sd 19072) * $signed(input_fmap_35[15:0]) +
	( 16'sd 26591) * $signed(input_fmap_36[15:0]) +
	( 15'sd 8942) * $signed(input_fmap_37[15:0]) +
	( 16'sd 29463) * $signed(input_fmap_38[15:0]) +
	( 15'sd 10358) * $signed(input_fmap_39[15:0]) +
	( 15'sd 13014) * $signed(input_fmap_40[15:0]) +
	( 14'sd 6909) * $signed(input_fmap_41[15:0]) +
	( 16'sd 17251) * $signed(input_fmap_42[15:0]) +
	( 16'sd 19599) * $signed(input_fmap_43[15:0]) +
	( 16'sd 30399) * $signed(input_fmap_44[15:0]) +
	( 13'sd 3600) * $signed(input_fmap_45[15:0]) +
	( 14'sd 4488) * $signed(input_fmap_46[15:0]) +
	( 16'sd 25614) * $signed(input_fmap_47[15:0]) +
	( 16'sd 28588) * $signed(input_fmap_48[15:0]) +
	( 16'sd 16924) * $signed(input_fmap_49[15:0]) +
	( 16'sd 20703) * $signed(input_fmap_50[15:0]) +
	( 15'sd 13177) * $signed(input_fmap_51[15:0]) +
	( 15'sd 14863) * $signed(input_fmap_52[15:0]) +
	( 16'sd 17852) * $signed(input_fmap_53[15:0]) +
	( 15'sd 11666) * $signed(input_fmap_54[15:0]) +
	( 15'sd 9086) * $signed(input_fmap_55[15:0]) +
	( 13'sd 2777) * $signed(input_fmap_56[15:0]) +
	( 16'sd 25179) * $signed(input_fmap_57[15:0]) +
	( 14'sd 5030) * $signed(input_fmap_58[15:0]) +
	( 16'sd 18863) * $signed(input_fmap_59[15:0]) +
	( 15'sd 14629) * $signed(input_fmap_60[15:0]) +
	( 16'sd 30988) * $signed(input_fmap_61[15:0]) +
	( 16'sd 17781) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20215) * $signed(input_fmap_63[15:0]) +
	( 16'sd 31462) * $signed(input_fmap_64[15:0]) +
	( 15'sd 9780) * $signed(input_fmap_65[15:0]) +
	( 15'sd 12730) * $signed(input_fmap_66[15:0]) +
	( 16'sd 20148) * $signed(input_fmap_67[15:0]) +
	( 16'sd 21947) * $signed(input_fmap_68[15:0]) +
	( 15'sd 14960) * $signed(input_fmap_69[15:0]) +
	( 15'sd 15504) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31867) * $signed(input_fmap_71[15:0]) +
	( 16'sd 17068) * $signed(input_fmap_72[15:0]) +
	( 15'sd 14111) * $signed(input_fmap_73[15:0]) +
	( 14'sd 7357) * $signed(input_fmap_74[15:0]) +
	( 16'sd 16964) * $signed(input_fmap_75[15:0]) +
	( 16'sd 20848) * $signed(input_fmap_76[15:0]) +
	( 16'sd 20706) * $signed(input_fmap_77[15:0]) +
	( 16'sd 24168) * $signed(input_fmap_78[15:0]) +
	( 13'sd 2628) * $signed(input_fmap_79[15:0]) +
	( 15'sd 12243) * $signed(input_fmap_80[15:0]) +
	( 15'sd 13918) * $signed(input_fmap_81[15:0]) +
	( 16'sd 22232) * $signed(input_fmap_82[15:0]) +
	( 15'sd 13673) * $signed(input_fmap_83[15:0]) +
	( 12'sd 1835) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24098) * $signed(input_fmap_85[15:0]) +
	( 16'sd 28754) * $signed(input_fmap_86[15:0]) +
	( 16'sd 22384) * $signed(input_fmap_87[15:0]) +
	( 8'sd 81) * $signed(input_fmap_88[15:0]) +
	( 13'sd 2665) * $signed(input_fmap_89[15:0]) +
	( 15'sd 13431) * $signed(input_fmap_90[15:0]) +
	( 14'sd 7242) * $signed(input_fmap_91[15:0]) +
	( 16'sd 23247) * $signed(input_fmap_92[15:0]) +
	( 15'sd 10486) * $signed(input_fmap_93[15:0]) +
	( 16'sd 21847) * $signed(input_fmap_94[15:0]) +
	( 15'sd 15126) * $signed(input_fmap_95[15:0]) +
	( 16'sd 31796) * $signed(input_fmap_96[15:0]) +
	( 15'sd 16078) * $signed(input_fmap_97[15:0]) +
	( 16'sd 27654) * $signed(input_fmap_98[15:0]) +
	( 13'sd 2103) * $signed(input_fmap_99[15:0]) +
	( 14'sd 4835) * $signed(input_fmap_100[15:0]) +
	( 13'sd 2353) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5771) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28948) * $signed(input_fmap_103[15:0]) +
	( 15'sd 9995) * $signed(input_fmap_104[15:0]) +
	( 16'sd 32045) * $signed(input_fmap_105[15:0]) +
	( 14'sd 5589) * $signed(input_fmap_106[15:0]) +
	( 14'sd 5766) * $signed(input_fmap_107[15:0]) +
	( 14'sd 4681) * $signed(input_fmap_108[15:0]) +
	( 16'sd 22446) * $signed(input_fmap_109[15:0]) +
	( 16'sd 30180) * $signed(input_fmap_110[15:0]) +
	( 16'sd 25824) * $signed(input_fmap_111[15:0]) +
	( 14'sd 4135) * $signed(input_fmap_112[15:0]) +
	( 15'sd 13827) * $signed(input_fmap_113[15:0]) +
	( 15'sd 14639) * $signed(input_fmap_114[15:0]) +
	( 13'sd 2488) * $signed(input_fmap_115[15:0]) +
	( 16'sd 18638) * $signed(input_fmap_116[15:0]) +
	( 15'sd 15586) * $signed(input_fmap_117[15:0]) +
	( 16'sd 31158) * $signed(input_fmap_118[15:0]) +
	( 16'sd 19618) * $signed(input_fmap_119[15:0]) +
	( 14'sd 5248) * $signed(input_fmap_120[15:0]) +
	( 16'sd 20013) * $signed(input_fmap_121[15:0]) +
	( 14'sd 5547) * $signed(input_fmap_122[15:0]) +
	( 16'sd 32331) * $signed(input_fmap_123[15:0]) +
	( 16'sd 24462) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24438) * $signed(input_fmap_125[15:0]) +
	( 16'sd 28907) * $signed(input_fmap_126[15:0]) +
	( 15'sd 14697) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 15'sd 15678) * $signed(input_fmap_0[15:0]) +
	( 12'sd 1254) * $signed(input_fmap_1[15:0]) +
	( 16'sd 25596) * $signed(input_fmap_2[15:0]) +
	( 15'sd 10551) * $signed(input_fmap_3[15:0]) +
	( 15'sd 11372) * $signed(input_fmap_4[15:0]) +
	( 16'sd 30480) * $signed(input_fmap_5[15:0]) +
	( 15'sd 11174) * $signed(input_fmap_6[15:0]) +
	( 15'sd 9361) * $signed(input_fmap_7[15:0]) +
	( 16'sd 30723) * $signed(input_fmap_8[15:0]) +
	( 7'sd 39) * $signed(input_fmap_9[15:0]) +
	( 16'sd 28785) * $signed(input_fmap_10[15:0]) +
	( 16'sd 26970) * $signed(input_fmap_11[15:0]) +
	( 15'sd 11045) * $signed(input_fmap_12[15:0]) +
	( 16'sd 18185) * $signed(input_fmap_13[15:0]) +
	( 16'sd 30615) * $signed(input_fmap_14[15:0]) +
	( 15'sd 11025) * $signed(input_fmap_15[15:0]) +
	( 14'sd 7016) * $signed(input_fmap_16[15:0]) +
	( 11'sd 700) * $signed(input_fmap_17[15:0]) +
	( 14'sd 4860) * $signed(input_fmap_18[15:0]) +
	( 16'sd 21165) * $signed(input_fmap_19[15:0]) +
	( 15'sd 10280) * $signed(input_fmap_20[15:0]) +
	( 15'sd 8916) * $signed(input_fmap_21[15:0]) +
	( 16'sd 23442) * $signed(input_fmap_22[15:0]) +
	( 14'sd 6882) * $signed(input_fmap_23[15:0]) +
	( 16'sd 21910) * $signed(input_fmap_24[15:0]) +
	( 16'sd 31561) * $signed(input_fmap_25[15:0]) +
	( 15'sd 13898) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9372) * $signed(input_fmap_27[15:0]) +
	( 15'sd 9496) * $signed(input_fmap_28[15:0]) +
	( 15'sd 12517) * $signed(input_fmap_29[15:0]) +
	( 12'sd 1239) * $signed(input_fmap_30[15:0]) +
	( 15'sd 14913) * $signed(input_fmap_31[15:0]) +
	( 15'sd 12851) * $signed(input_fmap_32[15:0]) +
	( 16'sd 31607) * $signed(input_fmap_33[15:0]) +
	( 8'sd 73) * $signed(input_fmap_34[15:0]) +
	( 11'sd 796) * $signed(input_fmap_35[15:0]) +
	( 14'sd 5066) * $signed(input_fmap_36[15:0]) +
	( 16'sd 22921) * $signed(input_fmap_37[15:0]) +
	( 13'sd 3973) * $signed(input_fmap_38[15:0]) +
	( 9'sd 202) * $signed(input_fmap_39[15:0]) +
	( 11'sd 592) * $signed(input_fmap_40[15:0]) +
	( 16'sd 25456) * $signed(input_fmap_41[15:0]) +
	( 16'sd 30895) * $signed(input_fmap_42[15:0]) +
	( 16'sd 24456) * $signed(input_fmap_43[15:0]) +
	( 15'sd 9878) * $signed(input_fmap_44[15:0]) +
	( 14'sd 4577) * $signed(input_fmap_45[15:0]) +
	( 16'sd 17812) * $signed(input_fmap_46[15:0]) +
	( 15'sd 8667) * $signed(input_fmap_47[15:0]) +
	( 15'sd 10797) * $signed(input_fmap_48[15:0]) +
	( 16'sd 18685) * $signed(input_fmap_49[15:0]) +
	( 15'sd 12094) * $signed(input_fmap_50[15:0]) +
	( 16'sd 16678) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3487) * $signed(input_fmap_52[15:0]) +
	( 15'sd 9913) * $signed(input_fmap_53[15:0]) +
	( 16'sd 20665) * $signed(input_fmap_54[15:0]) +
	( 15'sd 16271) * $signed(input_fmap_55[15:0]) +
	( 15'sd 8792) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17737) * $signed(input_fmap_57[15:0]) +
	( 16'sd 17070) * $signed(input_fmap_58[15:0]) +
	( 16'sd 24179) * $signed(input_fmap_59[15:0]) +
	( 16'sd 20928) * $signed(input_fmap_60[15:0]) +
	( 13'sd 3486) * $signed(input_fmap_61[15:0]) +
	( 16'sd 21961) * $signed(input_fmap_62[15:0]) +
	( 6'sd 26) * $signed(input_fmap_63[15:0]) +
	( 16'sd 22720) * $signed(input_fmap_64[15:0]) +
	( 14'sd 7601) * $signed(input_fmap_65[15:0]) +
	( 13'sd 2820) * $signed(input_fmap_66[15:0]) +
	( 16'sd 23735) * $signed(input_fmap_67[15:0]) +
	( 15'sd 13522) * $signed(input_fmap_68[15:0]) +
	( 16'sd 23183) * $signed(input_fmap_69[15:0]) +
	( 14'sd 8187) * $signed(input_fmap_70[15:0]) +
	( 13'sd 2637) * $signed(input_fmap_71[15:0]) +
	( 15'sd 16372) * $signed(input_fmap_72[15:0]) +
	( 16'sd 27188) * $signed(input_fmap_73[15:0]) +
	( 16'sd 20603) * $signed(input_fmap_74[15:0]) +
	( 14'sd 7704) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19815) * $signed(input_fmap_76[15:0]) +
	( 16'sd 29833) * $signed(input_fmap_77[15:0]) +
	( 14'sd 6365) * $signed(input_fmap_78[15:0]) +
	( 16'sd 26716) * $signed(input_fmap_79[15:0]) +
	( 15'sd 14528) * $signed(input_fmap_80[15:0]) +
	( 15'sd 8211) * $signed(input_fmap_81[15:0]) +
	( 16'sd 23243) * $signed(input_fmap_82[15:0]) +
	( 16'sd 17543) * $signed(input_fmap_83[15:0]) +
	( 13'sd 3157) * $signed(input_fmap_84[15:0]) +
	( 16'sd 22071) * $signed(input_fmap_85[15:0]) +
	( 15'sd 13655) * $signed(input_fmap_86[15:0]) +
	( 15'sd 10002) * $signed(input_fmap_87[15:0]) +
	( 15'sd 9489) * $signed(input_fmap_88[15:0]) +
	( 15'sd 14386) * $signed(input_fmap_89[15:0]) +
	( 15'sd 14547) * $signed(input_fmap_90[15:0]) +
	( 14'sd 5848) * $signed(input_fmap_91[15:0]) +
	( 13'sd 3337) * $signed(input_fmap_92[15:0]) +
	( 15'sd 8650) * $signed(input_fmap_93[15:0]) +
	( 14'sd 8122) * $signed(input_fmap_94[15:0]) +
	( 16'sd 29959) * $signed(input_fmap_95[15:0]) +
	( 15'sd 13938) * $signed(input_fmap_96[15:0]) +
	( 16'sd 18789) * $signed(input_fmap_97[15:0]) +
	( 16'sd 27904) * $signed(input_fmap_98[15:0]) +
	( 15'sd 11242) * $signed(input_fmap_99[15:0]) +
	( 14'sd 7165) * $signed(input_fmap_100[15:0]) +
	( 10'sd 359) * $signed(input_fmap_101[15:0]) +
	( 16'sd 28979) * $signed(input_fmap_102[15:0]) +
	( 16'sd 30847) * $signed(input_fmap_103[15:0]) +
	( 15'sd 11921) * $signed(input_fmap_104[15:0]) +
	( 16'sd 24133) * $signed(input_fmap_105[15:0]) +
	( 14'sd 7680) * $signed(input_fmap_106[15:0]) +
	( 13'sd 3110) * $signed(input_fmap_107[15:0]) +
	( 16'sd 24362) * $signed(input_fmap_108[15:0]) +
	( 14'sd 7200) * $signed(input_fmap_109[15:0]) +
	( 16'sd 20897) * $signed(input_fmap_110[15:0]) +
	( 12'sd 1643) * $signed(input_fmap_111[15:0]) +
	( 15'sd 10775) * $signed(input_fmap_112[15:0]) +
	( 16'sd 24383) * $signed(input_fmap_113[15:0]) +
	( 16'sd 28855) * $signed(input_fmap_114[15:0]) +
	( 16'sd 25372) * $signed(input_fmap_115[15:0]) +
	( 16'sd 25924) * $signed(input_fmap_116[15:0]) +
	( 10'sd 403) * $signed(input_fmap_117[15:0]) +
	( 15'sd 15724) * $signed(input_fmap_118[15:0]) +
	( 13'sd 3695) * $signed(input_fmap_119[15:0]) +
	( 15'sd 16106) * $signed(input_fmap_120[15:0]) +
	( 16'sd 28856) * $signed(input_fmap_121[15:0]) +
	( 13'sd 2622) * $signed(input_fmap_122[15:0]) +
	( 16'sd 29550) * $signed(input_fmap_123[15:0]) +
	( 15'sd 15194) * $signed(input_fmap_124[15:0]) +
	( 14'sd 5700) * $signed(input_fmap_125[15:0]) +
	( 16'sd 26754) * $signed(input_fmap_126[15:0]) +
	( 16'sd 23513) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 12'sd 1424) * $signed(input_fmap_0[15:0]) +
	( 15'sd 14658) * $signed(input_fmap_1[15:0]) +
	( 14'sd 7935) * $signed(input_fmap_2[15:0]) +
	( 16'sd 27878) * $signed(input_fmap_3[15:0]) +
	( 16'sd 22876) * $signed(input_fmap_4[15:0]) +
	( 16'sd 19059) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2118) * $signed(input_fmap_6[15:0]) +
	( 16'sd 31202) * $signed(input_fmap_7[15:0]) +
	( 14'sd 6396) * $signed(input_fmap_8[15:0]) +
	( 15'sd 10712) * $signed(input_fmap_9[15:0]) +
	( 16'sd 19116) * $signed(input_fmap_10[15:0]) +
	( 15'sd 16217) * $signed(input_fmap_11[15:0]) +
	( 14'sd 5304) * $signed(input_fmap_12[15:0]) +
	( 16'sd 21781) * $signed(input_fmap_13[15:0]) +
	( 13'sd 3095) * $signed(input_fmap_14[15:0]) +
	( 16'sd 24807) * $signed(input_fmap_15[15:0]) +
	( 16'sd 17467) * $signed(input_fmap_16[15:0]) +
	( 16'sd 21033) * $signed(input_fmap_17[15:0]) +
	( 13'sd 2199) * $signed(input_fmap_18[15:0]) +
	( 16'sd 21675) * $signed(input_fmap_19[15:0]) +
	( 15'sd 16101) * $signed(input_fmap_20[15:0]) +
	( 14'sd 4686) * $signed(input_fmap_21[15:0]) +
	( 13'sd 4055) * $signed(input_fmap_22[15:0]) +
	( 15'sd 9115) * $signed(input_fmap_23[15:0]) +
	( 12'sd 1830) * $signed(input_fmap_24[15:0]) +
	( 15'sd 13312) * $signed(input_fmap_25[15:0]) +
	( 14'sd 7994) * $signed(input_fmap_26[15:0]) +
	( 11'sd 894) * $signed(input_fmap_27[15:0]) +
	( 16'sd 20637) * $signed(input_fmap_28[15:0]) +
	( 16'sd 19967) * $signed(input_fmap_29[15:0]) +
	( 16'sd 21647) * $signed(input_fmap_30[15:0]) +
	( 16'sd 30268) * $signed(input_fmap_31[15:0]) +
	( 12'sd 1890) * $signed(input_fmap_32[15:0]) +
	( 16'sd 17037) * $signed(input_fmap_33[15:0]) +
	( 16'sd 31734) * $signed(input_fmap_34[15:0]) +
	( 16'sd 22364) * $signed(input_fmap_35[15:0]) +
	( 16'sd 27176) * $signed(input_fmap_36[15:0]) +
	( 13'sd 2781) * $signed(input_fmap_37[15:0]) +
	( 13'sd 2364) * $signed(input_fmap_38[15:0]) +
	( 16'sd 28359) * $signed(input_fmap_39[15:0]) +
	( 16'sd 19220) * $signed(input_fmap_40[15:0]) +
	( 16'sd 16727) * $signed(input_fmap_41[15:0]) +
	( 16'sd 22426) * $signed(input_fmap_42[15:0]) +
	( 16'sd 21388) * $signed(input_fmap_43[15:0]) +
	( 15'sd 10252) * $signed(input_fmap_44[15:0]) +
	( 15'sd 10509) * $signed(input_fmap_45[15:0]) +
	( 15'sd 15061) * $signed(input_fmap_46[15:0]) +
	( 12'sd 2035) * $signed(input_fmap_47[15:0]) +
	( 15'sd 15005) * $signed(input_fmap_48[15:0]) +
	( 15'sd 15404) * $signed(input_fmap_49[15:0]) +
	( 15'sd 14148) * $signed(input_fmap_50[15:0]) +
	( 16'sd 17853) * $signed(input_fmap_51[15:0]) +
	( 16'sd 16523) * $signed(input_fmap_52[15:0]) +
	( 16'sd 19499) * $signed(input_fmap_53[15:0]) +
	( 16'sd 20031) * $signed(input_fmap_54[15:0]) +
	( 16'sd 29497) * $signed(input_fmap_55[15:0]) +
	( 16'sd 26424) * $signed(input_fmap_56[15:0]) +
	( 16'sd 24277) * $signed(input_fmap_57[15:0]) +
	( 16'sd 29643) * $signed(input_fmap_58[15:0]) +
	( 16'sd 29514) * $signed(input_fmap_59[15:0]) +
	( 13'sd 3580) * $signed(input_fmap_60[15:0]) +
	( 15'sd 15030) * $signed(input_fmap_61[15:0]) +
	( 14'sd 6640) * $signed(input_fmap_62[15:0]) +
	( 16'sd 24117) * $signed(input_fmap_63[15:0]) +
	( 15'sd 10534) * $signed(input_fmap_64[15:0]) +
	( 13'sd 3414) * $signed(input_fmap_65[15:0]) +
	( 14'sd 7216) * $signed(input_fmap_66[15:0]) +
	( 16'sd 31066) * $signed(input_fmap_67[15:0]) +
	( 16'sd 18733) * $signed(input_fmap_68[15:0]) +
	( 15'sd 13012) * $signed(input_fmap_69[15:0]) +
	( 16'sd 22621) * $signed(input_fmap_70[15:0]) +
	( 16'sd 17127) * $signed(input_fmap_71[15:0]) +
	( 16'sd 28507) * $signed(input_fmap_72[15:0]) +
	( 15'sd 11785) * $signed(input_fmap_73[15:0]) +
	( 16'sd 19855) * $signed(input_fmap_74[15:0]) +
	( 13'sd 3574) * $signed(input_fmap_75[15:0]) +
	( 16'sd 20577) * $signed(input_fmap_76[15:0]) +
	( 16'sd 25587) * $signed(input_fmap_77[15:0]) +
	( 16'sd 28735) * $signed(input_fmap_78[15:0]) +
	( 16'sd 31603) * $signed(input_fmap_79[15:0]) +
	( 16'sd 17151) * $signed(input_fmap_80[15:0]) +
	( 15'sd 15554) * $signed(input_fmap_81[15:0]) +
	( 16'sd 24894) * $signed(input_fmap_82[15:0]) +
	( 16'sd 17184) * $signed(input_fmap_83[15:0]) +
	( 15'sd 13323) * $signed(input_fmap_84[15:0]) +
	( 15'sd 8823) * $signed(input_fmap_85[15:0]) +
	( 15'sd 12303) * $signed(input_fmap_86[15:0]) +
	( 15'sd 16211) * $signed(input_fmap_87[15:0]) +
	( 15'sd 13789) * $signed(input_fmap_88[15:0]) +
	( 16'sd 27324) * $signed(input_fmap_89[15:0]) +
	( 14'sd 5371) * $signed(input_fmap_90[15:0]) +
	( 15'sd 12615) * $signed(input_fmap_91[15:0]) +
	( 13'sd 2237) * $signed(input_fmap_92[15:0]) +
	( 16'sd 20518) * $signed(input_fmap_93[15:0]) +
	( 16'sd 28649) * $signed(input_fmap_94[15:0]) +
	( 13'sd 2633) * $signed(input_fmap_95[15:0]) +
	( 13'sd 2529) * $signed(input_fmap_96[15:0]) +
	( 15'sd 15161) * $signed(input_fmap_97[15:0]) +
	( 8'sd 85) * $signed(input_fmap_98[15:0]) +
	( 16'sd 20961) * $signed(input_fmap_99[15:0]) +
	( 16'sd 18196) * $signed(input_fmap_100[15:0]) +
	( 16'sd 16745) * $signed(input_fmap_101[15:0]) +
	( 15'sd 10691) * $signed(input_fmap_102[15:0]) +
	( 14'sd 5019) * $signed(input_fmap_103[15:0]) +
	( 15'sd 8914) * $signed(input_fmap_104[15:0]) +
	( 16'sd 23610) * $signed(input_fmap_105[15:0]) +
	( 16'sd 24895) * $signed(input_fmap_106[15:0]) +
	( 16'sd 16812) * $signed(input_fmap_107[15:0]) +
	( 16'sd 22453) * $signed(input_fmap_108[15:0]) +
	( 15'sd 8824) * $signed(input_fmap_109[15:0]) +
	( 14'sd 4280) * $signed(input_fmap_110[15:0]) +
	( 14'sd 4863) * $signed(input_fmap_111[15:0]) +
	( 16'sd 32101) * $signed(input_fmap_112[15:0]) +
	( 15'sd 15541) * $signed(input_fmap_113[15:0]) +
	( 15'sd 15693) * $signed(input_fmap_114[15:0]) +
	( 16'sd 21287) * $signed(input_fmap_115[15:0]) +
	( 16'sd 23376) * $signed(input_fmap_116[15:0]) +
	( 16'sd 17574) * $signed(input_fmap_117[15:0]) +
	( 14'sd 7235) * $signed(input_fmap_118[15:0]) +
	( 15'sd 11261) * $signed(input_fmap_119[15:0]) +
	( 16'sd 24209) * $signed(input_fmap_120[15:0]) +
	( 14'sd 7893) * $signed(input_fmap_121[15:0]) +
	( 14'sd 6442) * $signed(input_fmap_122[15:0]) +
	( 16'sd 25375) * $signed(input_fmap_123[15:0]) +
	( 16'sd 20323) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24482) * $signed(input_fmap_125[15:0]) +
	( 16'sd 23360) * $signed(input_fmap_126[15:0]) +
	( 15'sd 12490) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 14'sd 7608) * $signed(input_fmap_0[15:0]) +
	( 14'sd 4458) * $signed(input_fmap_1[15:0]) +
	( 16'sd 31855) * $signed(input_fmap_2[15:0]) +
	( 16'sd 29964) * $signed(input_fmap_3[15:0]) +
	( 14'sd 4805) * $signed(input_fmap_4[15:0]) +
	( 16'sd 24262) * $signed(input_fmap_5[15:0]) +
	( 16'sd 24220) * $signed(input_fmap_6[15:0]) +
	( 16'sd 18479) * $signed(input_fmap_7[15:0]) +
	( 16'sd 16619) * $signed(input_fmap_8[15:0]) +
	( 16'sd 28849) * $signed(input_fmap_9[15:0]) +
	( 13'sd 3974) * $signed(input_fmap_10[15:0]) +
	( 16'sd 27582) * $signed(input_fmap_11[15:0]) +
	( 16'sd 30362) * $signed(input_fmap_12[15:0]) +
	( 16'sd 19098) * $signed(input_fmap_13[15:0]) +
	( 16'sd 21901) * $signed(input_fmap_14[15:0]) +
	( 15'sd 15515) * $signed(input_fmap_15[15:0]) +
	( 14'sd 7893) * $signed(input_fmap_16[15:0]) +
	( 16'sd 24673) * $signed(input_fmap_17[15:0]) +
	( 16'sd 18757) * $signed(input_fmap_18[15:0]) +
	( 11'sd 838) * $signed(input_fmap_19[15:0]) +
	( 16'sd 25749) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17345) * $signed(input_fmap_21[15:0]) +
	( 15'sd 13052) * $signed(input_fmap_22[15:0]) +
	( 15'sd 10714) * $signed(input_fmap_23[15:0]) +
	( 16'sd 23536) * $signed(input_fmap_24[15:0]) +
	( 15'sd 14217) * $signed(input_fmap_25[15:0]) +
	( 14'sd 7384) * $signed(input_fmap_26[15:0]) +
	( 16'sd 19949) * $signed(input_fmap_27[15:0]) +
	( 13'sd 2928) * $signed(input_fmap_28[15:0]) +
	( 15'sd 15237) * $signed(input_fmap_29[15:0]) +
	( 15'sd 8575) * $signed(input_fmap_30[15:0]) +
	( 16'sd 21653) * $signed(input_fmap_31[15:0]) +
	( 16'sd 22247) * $signed(input_fmap_32[15:0]) +
	( 14'sd 5220) * $signed(input_fmap_33[15:0]) +
	( 15'sd 9953) * $signed(input_fmap_34[15:0]) +
	( 10'sd 314) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2132) * $signed(input_fmap_36[15:0]) +
	( 13'sd 3202) * $signed(input_fmap_37[15:0]) +
	( 14'sd 5021) * $signed(input_fmap_38[15:0]) +
	( 15'sd 10571) * $signed(input_fmap_39[15:0]) +
	( 16'sd 20528) * $signed(input_fmap_40[15:0]) +
	( 16'sd 20956) * $signed(input_fmap_41[15:0]) +
	( 14'sd 6334) * $signed(input_fmap_42[15:0]) +
	( 15'sd 8597) * $signed(input_fmap_43[15:0]) +
	( 13'sd 3933) * $signed(input_fmap_44[15:0]) +
	( 16'sd 26112) * $signed(input_fmap_45[15:0]) +
	( 13'sd 2949) * $signed(input_fmap_46[15:0]) +
	( 12'sd 1358) * $signed(input_fmap_47[15:0]) +
	( 16'sd 22315) * $signed(input_fmap_48[15:0]) +
	( 13'sd 3727) * $signed(input_fmap_49[15:0]) +
	( 11'sd 692) * $signed(input_fmap_50[15:0]) +
	( 15'sd 13181) * $signed(input_fmap_51[15:0]) +
	( 16'sd 22240) * $signed(input_fmap_52[15:0]) +
	( 15'sd 11022) * $signed(input_fmap_53[15:0]) +
	( 10'sd 412) * $signed(input_fmap_54[15:0]) +
	( 15'sd 12944) * $signed(input_fmap_55[15:0]) +
	( 15'sd 10034) * $signed(input_fmap_56[15:0]) +
	( 14'sd 5252) * $signed(input_fmap_57[15:0]) +
	( 14'sd 6564) * $signed(input_fmap_58[15:0]) +
	( 15'sd 15856) * $signed(input_fmap_59[15:0]) +
	( 15'sd 14826) * $signed(input_fmap_60[15:0]) +
	( 16'sd 32374) * $signed(input_fmap_61[15:0]) +
	( 15'sd 12813) * $signed(input_fmap_62[15:0]) +
	( 16'sd 31500) * $signed(input_fmap_63[15:0]) +
	( 14'sd 7770) * $signed(input_fmap_64[15:0]) +
	( 15'sd 14096) * $signed(input_fmap_65[15:0]) +
	( 15'sd 11832) * $signed(input_fmap_66[15:0]) +
	( 15'sd 8323) * $signed(input_fmap_67[15:0]) +
	( 15'sd 11236) * $signed(input_fmap_68[15:0]) +
	( 16'sd 22505) * $signed(input_fmap_69[15:0]) +
	( 15'sd 13373) * $signed(input_fmap_70[15:0]) +
	( 16'sd 19646) * $signed(input_fmap_71[15:0]) +
	( 16'sd 24731) * $signed(input_fmap_72[15:0]) +
	( 15'sd 11478) * $signed(input_fmap_73[15:0]) +
	( 16'sd 29625) * $signed(input_fmap_74[15:0]) +
	( 15'sd 9832) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19279) * $signed(input_fmap_76[15:0]) +
	( 15'sd 13226) * $signed(input_fmap_77[15:0]) +
	( 15'sd 9248) * $signed(input_fmap_78[15:0]) +
	( 16'sd 29971) * $signed(input_fmap_79[15:0]) +
	( 16'sd 16736) * $signed(input_fmap_80[15:0]) +
	( 16'sd 27766) * $signed(input_fmap_81[15:0]) +
	( 16'sd 31804) * $signed(input_fmap_82[15:0]) +
	( 11'sd 735) * $signed(input_fmap_83[15:0]) +
	( 16'sd 23031) * $signed(input_fmap_84[15:0]) +
	( 16'sd 27784) * $signed(input_fmap_85[15:0]) +
	( 16'sd 18826) * $signed(input_fmap_86[15:0]) +
	( 16'sd 31633) * $signed(input_fmap_87[15:0]) +
	( 16'sd 19193) * $signed(input_fmap_88[15:0]) +
	( 14'sd 7762) * $signed(input_fmap_89[15:0]) +
	( 14'sd 6271) * $signed(input_fmap_90[15:0]) +
	( 16'sd 31480) * $signed(input_fmap_91[15:0]) +
	( 14'sd 5816) * $signed(input_fmap_92[15:0]) +
	( 14'sd 5436) * $signed(input_fmap_93[15:0]) +
	( 16'sd 20469) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25622) * $signed(input_fmap_95[15:0]) +
	( 14'sd 6346) * $signed(input_fmap_96[15:0]) +
	( 16'sd 28685) * $signed(input_fmap_97[15:0]) +
	( 15'sd 12859) * $signed(input_fmap_98[15:0]) +
	( 13'sd 2424) * $signed(input_fmap_99[15:0]) +
	( 15'sd 9237) * $signed(input_fmap_100[15:0]) +
	( 16'sd 23361) * $signed(input_fmap_101[15:0]) +
	( 15'sd 11320) * $signed(input_fmap_102[15:0]) +
	( 15'sd 10635) * $signed(input_fmap_103[15:0]) +
	( 16'sd 29983) * $signed(input_fmap_104[15:0]) +
	( 15'sd 13466) * $signed(input_fmap_105[15:0]) +
	( 16'sd 32395) * $signed(input_fmap_106[15:0]) +
	( 16'sd 22718) * $signed(input_fmap_107[15:0]) +
	( 16'sd 20859) * $signed(input_fmap_108[15:0]) +
	( 13'sd 3206) * $signed(input_fmap_109[15:0]) +
	( 15'sd 15717) * $signed(input_fmap_110[15:0]) +
	( 15'sd 10795) * $signed(input_fmap_111[15:0]) +
	( 12'sd 1395) * $signed(input_fmap_112[15:0]) +
	( 16'sd 22152) * $signed(input_fmap_113[15:0]) +
	( 16'sd 19007) * $signed(input_fmap_114[15:0]) +
	( 15'sd 8448) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26916) * $signed(input_fmap_116[15:0]) +
	( 15'sd 11421) * $signed(input_fmap_117[15:0]) +
	( 16'sd 29075) * $signed(input_fmap_118[15:0]) +
	( 16'sd 28453) * $signed(input_fmap_119[15:0]) +
	( 16'sd 28687) * $signed(input_fmap_120[15:0]) +
	( 15'sd 13104) * $signed(input_fmap_121[15:0]) +
	( 14'sd 6517) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21286) * $signed(input_fmap_123[15:0]) +
	( 15'sd 8776) * $signed(input_fmap_124[15:0]) +
	( 16'sd 26098) * $signed(input_fmap_125[15:0]) +
	( 16'sd 31896) * $signed(input_fmap_126[15:0]) +
	( 15'sd 15789) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 12'sd 1607) * $signed(input_fmap_0[15:0]) +
	( 16'sd 21298) * $signed(input_fmap_1[15:0]) +
	( 15'sd 13451) * $signed(input_fmap_2[15:0]) +
	( 16'sd 24375) * $signed(input_fmap_3[15:0]) +
	( 16'sd 25118) * $signed(input_fmap_4[15:0]) +
	( 16'sd 16926) * $signed(input_fmap_5[15:0]) +
	( 16'sd 25208) * $signed(input_fmap_6[15:0]) +
	( 13'sd 3006) * $signed(input_fmap_7[15:0]) +
	( 15'sd 9282) * $signed(input_fmap_8[15:0]) +
	( 14'sd 4206) * $signed(input_fmap_9[15:0]) +
	( 16'sd 20585) * $signed(input_fmap_10[15:0]) +
	( 16'sd 31628) * $signed(input_fmap_11[15:0]) +
	( 15'sd 12304) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24171) * $signed(input_fmap_13[15:0]) +
	( 16'sd 25085) * $signed(input_fmap_14[15:0]) +
	( 12'sd 1814) * $signed(input_fmap_15[15:0]) +
	( 12'sd 1131) * $signed(input_fmap_16[15:0]) +
	( 15'sd 11397) * $signed(input_fmap_17[15:0]) +
	( 15'sd 10821) * $signed(input_fmap_18[15:0]) +
	( 16'sd 18998) * $signed(input_fmap_19[15:0]) +
	( 15'sd 14333) * $signed(input_fmap_20[15:0]) +
	( 15'sd 12040) * $signed(input_fmap_21[15:0]) +
	( 15'sd 16269) * $signed(input_fmap_22[15:0]) +
	( 14'sd 4784) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17751) * $signed(input_fmap_24[15:0]) +
	( 15'sd 9059) * $signed(input_fmap_25[15:0]) +
	( 12'sd 1096) * $signed(input_fmap_26[15:0]) +
	( 14'sd 5398) * $signed(input_fmap_27[15:0]) +
	( 16'sd 19198) * $signed(input_fmap_28[15:0]) +
	( 15'sd 9315) * $signed(input_fmap_29[15:0]) +
	( 15'sd 9410) * $signed(input_fmap_30[15:0]) +
	( 15'sd 13456) * $signed(input_fmap_31[15:0]) +
	( 15'sd 12074) * $signed(input_fmap_32[15:0]) +
	( 16'sd 32191) * $signed(input_fmap_33[15:0]) +
	( 16'sd 30431) * $signed(input_fmap_34[15:0]) +
	( 15'sd 14592) * $signed(input_fmap_35[15:0]) +
	( 15'sd 13267) * $signed(input_fmap_36[15:0]) +
	( 16'sd 32710) * $signed(input_fmap_37[15:0]) +
	( 15'sd 15400) * $signed(input_fmap_38[15:0]) +
	( 12'sd 1052) * $signed(input_fmap_39[15:0]) +
	( 16'sd 26028) * $signed(input_fmap_40[15:0]) +
	( 16'sd 23450) * $signed(input_fmap_41[15:0]) +
	( 16'sd 29632) * $signed(input_fmap_42[15:0]) +
	( 15'sd 8353) * $signed(input_fmap_43[15:0]) +
	( 16'sd 20319) * $signed(input_fmap_44[15:0]) +
	( 16'sd 20100) * $signed(input_fmap_45[15:0]) +
	( 15'sd 12624) * $signed(input_fmap_46[15:0]) +
	( 16'sd 25219) * $signed(input_fmap_47[15:0]) +
	( 16'sd 23118) * $signed(input_fmap_48[15:0]) +
	( 15'sd 12424) * $signed(input_fmap_49[15:0]) +
	( 16'sd 30570) * $signed(input_fmap_50[15:0]) +
	( 15'sd 9788) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3649) * $signed(input_fmap_52[15:0]) +
	( 15'sd 8213) * $signed(input_fmap_53[15:0]) +
	( 16'sd 26304) * $signed(input_fmap_54[15:0]) +
	( 15'sd 9790) * $signed(input_fmap_55[15:0]) +
	( 15'sd 8767) * $signed(input_fmap_56[15:0]) +
	( 12'sd 1676) * $signed(input_fmap_57[15:0]) +
	( 15'sd 8945) * $signed(input_fmap_58[15:0]) +
	( 15'sd 13573) * $signed(input_fmap_59[15:0]) +
	( 16'sd 18325) * $signed(input_fmap_60[15:0]) +
	( 13'sd 3981) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3882) * $signed(input_fmap_62[15:0]) +
	( 14'sd 5717) * $signed(input_fmap_63[15:0]) +
	( 16'sd 27805) * $signed(input_fmap_64[15:0]) +
	( 15'sd 10000) * $signed(input_fmap_65[15:0]) +
	( 16'sd 23058) * $signed(input_fmap_66[15:0]) +
	( 13'sd 3989) * $signed(input_fmap_67[15:0]) +
	( 16'sd 24329) * $signed(input_fmap_68[15:0]) +
	( 16'sd 28601) * $signed(input_fmap_69[15:0]) +
	( 16'sd 30586) * $signed(input_fmap_70[15:0]) +
	( 16'sd 25117) * $signed(input_fmap_71[15:0]) +
	( 15'sd 8228) * $signed(input_fmap_72[15:0]) +
	( 15'sd 15851) * $signed(input_fmap_73[15:0]) +
	( 13'sd 2578) * $signed(input_fmap_74[15:0]) +
	( 16'sd 16942) * $signed(input_fmap_75[15:0]) +
	( 16'sd 22472) * $signed(input_fmap_76[15:0]) +
	( 15'sd 9525) * $signed(input_fmap_77[15:0]) +
	( 14'sd 4832) * $signed(input_fmap_78[15:0]) +
	( 16'sd 29931) * $signed(input_fmap_79[15:0]) +
	( 12'sd 1025) * $signed(input_fmap_80[15:0]) +
	( 16'sd 25426) * $signed(input_fmap_81[15:0]) +
	( 15'sd 9364) * $signed(input_fmap_82[15:0]) +
	( 15'sd 15814) * $signed(input_fmap_83[15:0]) +
	( 15'sd 11643) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24996) * $signed(input_fmap_85[15:0]) +
	( 16'sd 19265) * $signed(input_fmap_86[15:0]) +
	( 16'sd 24799) * $signed(input_fmap_87[15:0]) +
	( 15'sd 15919) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5116) * $signed(input_fmap_89[15:0]) +
	( 16'sd 22344) * $signed(input_fmap_90[15:0]) +
	( 15'sd 10930) * $signed(input_fmap_91[15:0]) +
	( 16'sd 21779) * $signed(input_fmap_92[15:0]) +
	( 16'sd 24932) * $signed(input_fmap_93[15:0]) +
	( 16'sd 32112) * $signed(input_fmap_94[15:0]) +
	( 16'sd 17760) * $signed(input_fmap_95[15:0]) +
	( 15'sd 8670) * $signed(input_fmap_96[15:0]) +
	( 16'sd 28507) * $signed(input_fmap_97[15:0]) +
	( 15'sd 13250) * $signed(input_fmap_98[15:0]) +
	( 15'sd 9596) * $signed(input_fmap_99[15:0]) +
	( 15'sd 15759) * $signed(input_fmap_100[15:0]) +
	( 16'sd 19470) * $signed(input_fmap_101[15:0]) +
	( 15'sd 11682) * $signed(input_fmap_102[15:0]) +
	( 16'sd 27598) * $signed(input_fmap_103[15:0]) +
	( 12'sd 1852) * $signed(input_fmap_104[15:0]) +
	( 15'sd 15632) * $signed(input_fmap_105[15:0]) +
	( 15'sd 11926) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27765) * $signed(input_fmap_107[15:0]) +
	( 16'sd 21108) * $signed(input_fmap_108[15:0]) +
	( 15'sd 13295) * $signed(input_fmap_109[15:0]) +
	( 16'sd 29316) * $signed(input_fmap_110[15:0]) +
	( 16'sd 31837) * $signed(input_fmap_111[15:0]) +
	( 15'sd 14047) * $signed(input_fmap_112[15:0]) +
	( 16'sd 27365) * $signed(input_fmap_113[15:0]) +
	( 15'sd 10469) * $signed(input_fmap_114[15:0]) +
	( 14'sd 6590) * $signed(input_fmap_115[15:0]) +
	( 16'sd 21985) * $signed(input_fmap_116[15:0]) +
	( 15'sd 15252) * $signed(input_fmap_117[15:0]) +
	( 15'sd 14638) * $signed(input_fmap_118[15:0]) +
	( 16'sd 18223) * $signed(input_fmap_119[15:0]) +
	( 13'sd 3956) * $signed(input_fmap_120[15:0]) +
	( 16'sd 20946) * $signed(input_fmap_121[15:0]) +
	( 16'sd 30885) * $signed(input_fmap_122[15:0]) +
	( 15'sd 11899) * $signed(input_fmap_123[15:0]) +
	( 11'sd 968) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24306) * $signed(input_fmap_125[15:0]) +
	( 16'sd 17501) * $signed(input_fmap_126[15:0]) +
	( 16'sd 26238) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 16'sd 26531) * $signed(input_fmap_0[15:0]) +
	( 15'sd 15823) * $signed(input_fmap_1[15:0]) +
	( 16'sd 26688) * $signed(input_fmap_2[15:0]) +
	( 15'sd 9524) * $signed(input_fmap_3[15:0]) +
	( 13'sd 4028) * $signed(input_fmap_4[15:0]) +
	( 16'sd 16926) * $signed(input_fmap_5[15:0]) +
	( 16'sd 28095) * $signed(input_fmap_6[15:0]) +
	( 16'sd 17341) * $signed(input_fmap_7[15:0]) +
	( 15'sd 8500) * $signed(input_fmap_8[15:0]) +
	( 15'sd 14326) * $signed(input_fmap_9[15:0]) +
	( 16'sd 21722) * $signed(input_fmap_10[15:0]) +
	( 13'sd 2751) * $signed(input_fmap_11[15:0]) +
	( 14'sd 7157) * $signed(input_fmap_12[15:0]) +
	( 15'sd 13656) * $signed(input_fmap_13[15:0]) +
	( 16'sd 22354) * $signed(input_fmap_14[15:0]) +
	( 16'sd 29427) * $signed(input_fmap_15[15:0]) +
	( 15'sd 16148) * $signed(input_fmap_16[15:0]) +
	( 16'sd 19064) * $signed(input_fmap_17[15:0]) +
	( 16'sd 16466) * $signed(input_fmap_18[15:0]) +
	( 16'sd 25499) * $signed(input_fmap_19[15:0]) +
	( 9'sd 211) * $signed(input_fmap_20[15:0]) +
	( 14'sd 4621) * $signed(input_fmap_21[15:0]) +
	( 16'sd 22710) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28753) * $signed(input_fmap_23[15:0]) +
	( 16'sd 31721) * $signed(input_fmap_24[15:0]) +
	( 16'sd 32399) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22894) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9089) * $signed(input_fmap_27[15:0]) +
	( 15'sd 14125) * $signed(input_fmap_28[15:0]) +
	( 16'sd 25447) * $signed(input_fmap_29[15:0]) +
	( 12'sd 1781) * $signed(input_fmap_30[15:0]) +
	( 16'sd 22948) * $signed(input_fmap_31[15:0]) +
	( 16'sd 21976) * $signed(input_fmap_32[15:0]) +
	( 16'sd 25447) * $signed(input_fmap_33[15:0]) +
	( 14'sd 6520) * $signed(input_fmap_34[15:0]) +
	( 13'sd 3346) * $signed(input_fmap_35[15:0]) +
	( 15'sd 13796) * $signed(input_fmap_36[15:0]) +
	( 13'sd 3945) * $signed(input_fmap_37[15:0]) +
	( 16'sd 32077) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24859) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6324) * $signed(input_fmap_40[15:0]) +
	( 16'sd 25528) * $signed(input_fmap_41[15:0]) +
	( 16'sd 29863) * $signed(input_fmap_42[15:0]) +
	( 16'sd 31947) * $signed(input_fmap_43[15:0]) +
	( 16'sd 17579) * $signed(input_fmap_44[15:0]) +
	( 15'sd 9136) * $signed(input_fmap_45[15:0]) +
	( 15'sd 14851) * $signed(input_fmap_46[15:0]) +
	( 12'sd 1242) * $signed(input_fmap_47[15:0]) +
	( 16'sd 17276) * $signed(input_fmap_48[15:0]) +
	( 16'sd 17234) * $signed(input_fmap_49[15:0]) +
	( 15'sd 14531) * $signed(input_fmap_50[15:0]) +
	( 16'sd 23905) * $signed(input_fmap_51[15:0]) +
	( 15'sd 9084) * $signed(input_fmap_52[15:0]) +
	( 10'sd 325) * $signed(input_fmap_53[15:0]) +
	( 13'sd 2310) * $signed(input_fmap_54[15:0]) +
	( 16'sd 25186) * $signed(input_fmap_55[15:0]) +
	( 15'sd 15347) * $signed(input_fmap_56[15:0]) +
	( 14'sd 6840) * $signed(input_fmap_57[15:0]) +
	( 15'sd 8918) * $signed(input_fmap_58[15:0]) +
	( 16'sd 21084) * $signed(input_fmap_59[15:0]) +
	( 15'sd 8303) * $signed(input_fmap_60[15:0]) +
	( 15'sd 8508) * $signed(input_fmap_61[15:0]) +
	( 15'sd 11934) * $signed(input_fmap_62[15:0]) +
	( 13'sd 3867) * $signed(input_fmap_63[15:0]) +
	( 14'sd 5014) * $signed(input_fmap_64[15:0]) +
	( 16'sd 19261) * $signed(input_fmap_65[15:0]) +
	( 15'sd 11846) * $signed(input_fmap_66[15:0]) +
	( 14'sd 5945) * $signed(input_fmap_67[15:0]) +
	( 16'sd 28627) * $signed(input_fmap_68[15:0]) +
	( 16'sd 21046) * $signed(input_fmap_69[15:0]) +
	( 16'sd 28277) * $signed(input_fmap_70[15:0]) +
	( 13'sd 3140) * $signed(input_fmap_71[15:0]) +
	( 12'sd 2018) * $signed(input_fmap_72[15:0]) +
	( 15'sd 10036) * $signed(input_fmap_73[15:0]) +
	( 16'sd 23117) * $signed(input_fmap_74[15:0]) +
	( 14'sd 4117) * $signed(input_fmap_75[15:0]) +
	( 16'sd 22646) * $signed(input_fmap_76[15:0]) +
	( 14'sd 7182) * $signed(input_fmap_77[15:0]) +
	( 15'sd 10078) * $signed(input_fmap_78[15:0]) +
	( 16'sd 17930) * $signed(input_fmap_79[15:0]) +
	( 15'sd 9166) * $signed(input_fmap_80[15:0]) +
	( 16'sd 29718) * $signed(input_fmap_81[15:0]) +
	( 15'sd 13917) * $signed(input_fmap_82[15:0]) +
	( 15'sd 14858) * $signed(input_fmap_83[15:0]) +
	( 14'sd 6163) * $signed(input_fmap_84[15:0]) +
	( 14'sd 4921) * $signed(input_fmap_85[15:0]) +
	( 14'sd 7063) * $signed(input_fmap_86[15:0]) +
	( 14'sd 6792) * $signed(input_fmap_87[15:0]) +
	( 16'sd 22758) * $signed(input_fmap_88[15:0]) +
	( 13'sd 3733) * $signed(input_fmap_89[15:0]) +
	( 16'sd 20515) * $signed(input_fmap_90[15:0]) +
	( 15'sd 15121) * $signed(input_fmap_91[15:0]) +
	( 10'sd 347) * $signed(input_fmap_92[15:0]) +
	( 15'sd 15779) * $signed(input_fmap_93[15:0]) +
	( 15'sd 14551) * $signed(input_fmap_94[15:0]) +
	( 14'sd 8016) * $signed(input_fmap_95[15:0]) +
	( 16'sd 26052) * $signed(input_fmap_96[15:0]) +
	( 16'sd 19309) * $signed(input_fmap_97[15:0]) +
	( 16'sd 17335) * $signed(input_fmap_98[15:0]) +
	( 16'sd 31085) * $signed(input_fmap_99[15:0]) +
	( 14'sd 6704) * $signed(input_fmap_100[15:0]) +
	( 15'sd 9582) * $signed(input_fmap_101[15:0]) +
	( 14'sd 4106) * $signed(input_fmap_102[15:0]) +
	( 15'sd 10927) * $signed(input_fmap_103[15:0]) +
	( 16'sd 23348) * $signed(input_fmap_104[15:0]) +
	( 15'sd 9799) * $signed(input_fmap_105[15:0]) +
	( 16'sd 31973) * $signed(input_fmap_106[15:0]) +
	( 15'sd 14634) * $signed(input_fmap_107[15:0]) +
	( 16'sd 23550) * $signed(input_fmap_108[15:0]) +
	( 16'sd 16504) * $signed(input_fmap_109[15:0]) +
	( 16'sd 30721) * $signed(input_fmap_110[15:0]) +
	( 16'sd 32671) * $signed(input_fmap_111[15:0]) +
	( 16'sd 18037) * $signed(input_fmap_112[15:0]) +
	( 14'sd 7558) * $signed(input_fmap_113[15:0]) +
	( 16'sd 16989) * $signed(input_fmap_114[15:0]) +
	( 15'sd 14320) * $signed(input_fmap_115[15:0]) +
	( 16'sd 24061) * $signed(input_fmap_116[15:0]) +
	( 10'sd 382) * $signed(input_fmap_117[15:0]) +
	( 15'sd 9173) * $signed(input_fmap_118[15:0]) +
	( 16'sd 17625) * $signed(input_fmap_119[15:0]) +
	( 16'sd 28959) * $signed(input_fmap_120[15:0]) +
	( 16'sd 32503) * $signed(input_fmap_121[15:0]) +
	( 16'sd 27837) * $signed(input_fmap_122[15:0]) +
	( 15'sd 12541) * $signed(input_fmap_123[15:0]) +
	( 16'sd 29324) * $signed(input_fmap_124[15:0]) +
	( 14'sd 5833) * $signed(input_fmap_125[15:0]) +
	( 15'sd 14514) * $signed(input_fmap_126[15:0]) +
	( 16'sd 22447) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 14'sd 5387) * $signed(input_fmap_0[15:0]) +
	( 15'sd 14008) * $signed(input_fmap_1[15:0]) +
	( 16'sd 26356) * $signed(input_fmap_2[15:0]) +
	( 16'sd 25127) * $signed(input_fmap_3[15:0]) +
	( 16'sd 17911) * $signed(input_fmap_4[15:0]) +
	( 14'sd 4779) * $signed(input_fmap_5[15:0]) +
	( 16'sd 22166) * $signed(input_fmap_6[15:0]) +
	( 16'sd 17749) * $signed(input_fmap_7[15:0]) +
	( 16'sd 30238) * $signed(input_fmap_8[15:0]) +
	( 16'sd 17528) * $signed(input_fmap_9[15:0]) +
	( 10'sd 504) * $signed(input_fmap_10[15:0]) +
	( 10'sd 276) * $signed(input_fmap_11[15:0]) +
	( 16'sd 30983) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24935) * $signed(input_fmap_13[15:0]) +
	( 15'sd 13213) * $signed(input_fmap_14[15:0]) +
	( 16'sd 32224) * $signed(input_fmap_15[15:0]) +
	( 15'sd 14206) * $signed(input_fmap_16[15:0]) +
	( 15'sd 16104) * $signed(input_fmap_17[15:0]) +
	( 14'sd 6739) * $signed(input_fmap_18[15:0]) +
	( 16'sd 28135) * $signed(input_fmap_19[15:0]) +
	( 10'sd 438) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17599) * $signed(input_fmap_21[15:0]) +
	( 12'sd 1509) * $signed(input_fmap_22[15:0]) +
	( 16'sd 26872) * $signed(input_fmap_23[15:0]) +
	( 10'sd 386) * $signed(input_fmap_24[15:0]) +
	( 16'sd 19075) * $signed(input_fmap_25[15:0]) +
	( 16'sd 16940) * $signed(input_fmap_26[15:0]) +
	( 15'sd 9135) * $signed(input_fmap_27[15:0]) +
	( 13'sd 2799) * $signed(input_fmap_28[15:0]) +
	( 16'sd 23566) * $signed(input_fmap_29[15:0]) +
	( 16'sd 28788) * $signed(input_fmap_30[15:0]) +
	( 16'sd 22899) * $signed(input_fmap_31[15:0]) +
	( 16'sd 23226) * $signed(input_fmap_32[15:0]) +
	( 16'sd 26697) * $signed(input_fmap_33[15:0]) +
	( 15'sd 15381) * $signed(input_fmap_34[15:0]) +
	( 16'sd 25369) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2162) * $signed(input_fmap_36[15:0]) +
	( 16'sd 30938) * $signed(input_fmap_37[15:0]) +
	( 16'sd 22875) * $signed(input_fmap_38[15:0]) +
	( 16'sd 30103) * $signed(input_fmap_39[15:0]) +
	( 16'sd 28079) * $signed(input_fmap_40[15:0]) +
	( 13'sd 2341) * $signed(input_fmap_41[15:0]) +
	( 16'sd 18484) * $signed(input_fmap_42[15:0]) +
	( 16'sd 16417) * $signed(input_fmap_43[15:0]) +
	( 15'sd 8334) * $signed(input_fmap_44[15:0]) +
	( 15'sd 12241) * $signed(input_fmap_45[15:0]) +
	( 16'sd 28323) * $signed(input_fmap_46[15:0]) +
	( 15'sd 12980) * $signed(input_fmap_47[15:0]) +
	( 13'sd 3524) * $signed(input_fmap_48[15:0]) +
	( 16'sd 24391) * $signed(input_fmap_49[15:0]) +
	( 16'sd 24293) * $signed(input_fmap_50[15:0]) +
	( 14'sd 6135) * $signed(input_fmap_51[15:0]) +
	( 14'sd 4312) * $signed(input_fmap_52[15:0]) +
	( 15'sd 14181) * $signed(input_fmap_53[15:0]) +
	( 16'sd 18249) * $signed(input_fmap_54[15:0]) +
	( 10'sd 493) * $signed(input_fmap_55[15:0]) +
	( 16'sd 25280) * $signed(input_fmap_56[15:0]) +
	( 16'sd 21708) * $signed(input_fmap_57[15:0]) +
	( 10'sd 346) * $signed(input_fmap_58[15:0]) +
	( 16'sd 28620) * $signed(input_fmap_59[15:0]) +
	( 16'sd 28884) * $signed(input_fmap_60[15:0]) +
	( 15'sd 9905) * $signed(input_fmap_61[15:0]) +
	( 16'sd 23511) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20425) * $signed(input_fmap_63[15:0]) +
	( 15'sd 13474) * $signed(input_fmap_64[15:0]) +
	( 15'sd 12977) * $signed(input_fmap_65[15:0]) +
	( 16'sd 21269) * $signed(input_fmap_66[15:0]) +
	( 16'sd 30710) * $signed(input_fmap_67[15:0]) +
	( 14'sd 7338) * $signed(input_fmap_68[15:0]) +
	( 16'sd 32731) * $signed(input_fmap_69[15:0]) +
	( 16'sd 18470) * $signed(input_fmap_70[15:0]) +
	( 13'sd 3742) * $signed(input_fmap_71[15:0]) +
	( 16'sd 30181) * $signed(input_fmap_72[15:0]) +
	( 16'sd 21589) * $signed(input_fmap_73[15:0]) +
	( 16'sd 23707) * $signed(input_fmap_74[15:0]) +
	( 15'sd 8648) * $signed(input_fmap_75[15:0]) +
	( 16'sd 25889) * $signed(input_fmap_76[15:0]) +
	( 16'sd 21313) * $signed(input_fmap_77[15:0]) +
	( 16'sd 27828) * $signed(input_fmap_78[15:0]) +
	( 15'sd 9441) * $signed(input_fmap_79[15:0]) +
	( 16'sd 24232) * $signed(input_fmap_80[15:0]) +
	( 15'sd 13667) * $signed(input_fmap_81[15:0]) +
	( 12'sd 1389) * $signed(input_fmap_82[15:0]) +
	( 16'sd 23347) * $signed(input_fmap_83[15:0]) +
	( 16'sd 30065) * $signed(input_fmap_84[15:0]) +
	( 13'sd 2572) * $signed(input_fmap_85[15:0]) +
	( 15'sd 8734) * $signed(input_fmap_86[15:0]) +
	( 16'sd 27237) * $signed(input_fmap_87[15:0]) +
	( 15'sd 11499) * $signed(input_fmap_88[15:0]) +
	( 16'sd 28707) * $signed(input_fmap_89[15:0]) +
	( 15'sd 15358) * $signed(input_fmap_90[15:0]) +
	( 15'sd 9497) * $signed(input_fmap_91[15:0]) +
	( 16'sd 21527) * $signed(input_fmap_92[15:0]) +
	( 16'sd 29107) * $signed(input_fmap_93[15:0]) +
	( 16'sd 17173) * $signed(input_fmap_94[15:0]) +
	( 16'sd 18983) * $signed(input_fmap_95[15:0]) +
	( 15'sd 12652) * $signed(input_fmap_96[15:0]) +
	( 16'sd 32326) * $signed(input_fmap_97[15:0]) +
	( 13'sd 2485) * $signed(input_fmap_98[15:0]) +
	( 15'sd 8229) * $signed(input_fmap_99[15:0]) +
	( 16'sd 22381) * $signed(input_fmap_100[15:0]) +
	( 12'sd 1280) * $signed(input_fmap_101[15:0]) +
	( 16'sd 28020) * $signed(input_fmap_102[15:0]) +
	( 16'sd 29303) * $signed(input_fmap_103[15:0]) +
	( 15'sd 15067) * $signed(input_fmap_104[15:0]) +
	( 16'sd 18391) * $signed(input_fmap_105[15:0]) +
	( 16'sd 16814) * $signed(input_fmap_106[15:0]) +
	( 15'sd 13827) * $signed(input_fmap_107[15:0]) +
	( 16'sd 22734) * $signed(input_fmap_108[15:0]) +
	( 16'sd 16765) * $signed(input_fmap_109[15:0]) +
	( 16'sd 30642) * $signed(input_fmap_110[15:0]) +
	( 14'sd 6910) * $signed(input_fmap_111[15:0]) +
	( 15'sd 15762) * $signed(input_fmap_112[15:0]) +
	( 16'sd 26163) * $signed(input_fmap_113[15:0]) +
	( 15'sd 10755) * $signed(input_fmap_114[15:0]) +
	( 15'sd 12100) * $signed(input_fmap_115[15:0]) +
	( 11'sd 827) * $signed(input_fmap_116[15:0]) +
	( 16'sd 25577) * $signed(input_fmap_117[15:0]) +
	( 16'sd 20967) * $signed(input_fmap_118[15:0]) +
	( 15'sd 13367) * $signed(input_fmap_119[15:0]) +
	( 16'sd 25650) * $signed(input_fmap_120[15:0]) +
	( 16'sd 30958) * $signed(input_fmap_121[15:0]) +
	( 16'sd 25895) * $signed(input_fmap_122[15:0]) +
	( 16'sd 18868) * $signed(input_fmap_123[15:0]) +
	( 16'sd 18228) * $signed(input_fmap_124[15:0]) +
	( 16'sd 27468) * $signed(input_fmap_125[15:0]) +
	( 15'sd 11980) * $signed(input_fmap_126[15:0]) +
	( 16'sd 29922) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 14'sd 6050) * $signed(input_fmap_0[15:0]) +
	( 15'sd 8807) * $signed(input_fmap_1[15:0]) +
	( 16'sd 25393) * $signed(input_fmap_2[15:0]) +
	( 13'sd 2185) * $signed(input_fmap_3[15:0]) +
	( 14'sd 7023) * $signed(input_fmap_4[15:0]) +
	( 16'sd 16674) * $signed(input_fmap_5[15:0]) +
	( 16'sd 23497) * $signed(input_fmap_6[15:0]) +
	( 15'sd 15422) * $signed(input_fmap_7[15:0]) +
	( 15'sd 8598) * $signed(input_fmap_8[15:0]) +
	( 14'sd 6797) * $signed(input_fmap_9[15:0]) +
	( 16'sd 24278) * $signed(input_fmap_10[15:0]) +
	( 11'sd 834) * $signed(input_fmap_11[15:0]) +
	( 16'sd 17955) * $signed(input_fmap_12[15:0]) +
	( 14'sd 5490) * $signed(input_fmap_13[15:0]) +
	( 16'sd 32676) * $signed(input_fmap_14[15:0]) +
	( 16'sd 18193) * $signed(input_fmap_15[15:0]) +
	( 16'sd 25872) * $signed(input_fmap_16[15:0]) +
	( 16'sd 18665) * $signed(input_fmap_17[15:0]) +
	( 15'sd 12603) * $signed(input_fmap_18[15:0]) +
	( 16'sd 28930) * $signed(input_fmap_19[15:0]) +
	( 16'sd 32158) * $signed(input_fmap_20[15:0]) +
	( 16'sd 30652) * $signed(input_fmap_21[15:0]) +
	( 16'sd 26830) * $signed(input_fmap_22[15:0]) +
	( 16'sd 22394) * $signed(input_fmap_23[15:0]) +
	( 15'sd 9385) * $signed(input_fmap_24[15:0]) +
	( 16'sd 32560) * $signed(input_fmap_25[15:0]) +
	( 16'sd 28179) * $signed(input_fmap_26[15:0]) +
	( 15'sd 10042) * $signed(input_fmap_27[15:0]) +
	( 14'sd 6137) * $signed(input_fmap_28[15:0]) +
	( 16'sd 20662) * $signed(input_fmap_29[15:0]) +
	( 16'sd 21761) * $signed(input_fmap_30[15:0]) +
	( 16'sd 20292) * $signed(input_fmap_31[15:0]) +
	( 16'sd 31763) * $signed(input_fmap_32[15:0]) +
	( 15'sd 10934) * $signed(input_fmap_33[15:0]) +
	( 15'sd 11522) * $signed(input_fmap_34[15:0]) +
	( 16'sd 17630) * $signed(input_fmap_35[15:0]) +
	( 16'sd 32038) * $signed(input_fmap_36[15:0]) +
	( 16'sd 29870) * $signed(input_fmap_37[15:0]) +
	( 14'sd 7122) * $signed(input_fmap_38[15:0]) +
	( 16'sd 25311) * $signed(input_fmap_39[15:0]) +
	( 16'sd 18519) * $signed(input_fmap_40[15:0]) +
	( 16'sd 31621) * $signed(input_fmap_41[15:0]) +
	( 14'sd 6252) * $signed(input_fmap_42[15:0]) +
	( 16'sd 21335) * $signed(input_fmap_43[15:0]) +
	( 16'sd 32480) * $signed(input_fmap_44[15:0]) +
	( 16'sd 25013) * $signed(input_fmap_45[15:0]) +
	( 16'sd 31328) * $signed(input_fmap_46[15:0]) +
	( 15'sd 11891) * $signed(input_fmap_47[15:0]) +
	( 16'sd 23196) * $signed(input_fmap_48[15:0]) +
	( 16'sd 21371) * $signed(input_fmap_49[15:0]) +
	( 15'sd 15245) * $signed(input_fmap_50[15:0]) +
	( 16'sd 18243) * $signed(input_fmap_51[15:0]) +
	( 16'sd 29402) * $signed(input_fmap_52[15:0]) +
	( 16'sd 28327) * $signed(input_fmap_53[15:0]) +
	( 16'sd 32186) * $signed(input_fmap_54[15:0]) +
	( 15'sd 11853) * $signed(input_fmap_55[15:0]) +
	( 16'sd 20697) * $signed(input_fmap_56[15:0]) +
	( 16'sd 30915) * $signed(input_fmap_57[15:0]) +
	( 15'sd 15175) * $signed(input_fmap_58[15:0]) +
	( 16'sd 31995) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1253) * $signed(input_fmap_60[15:0]) +
	( 16'sd 18087) * $signed(input_fmap_61[15:0]) +
	( 16'sd 27643) * $signed(input_fmap_62[15:0]) +
	( 14'sd 5926) * $signed(input_fmap_63[15:0]) +
	( 14'sd 7689) * $signed(input_fmap_64[15:0]) +
	( 16'sd 24999) * $signed(input_fmap_65[15:0]) +
	( 15'sd 9845) * $signed(input_fmap_66[15:0]) +
	( 14'sd 4395) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26075) * $signed(input_fmap_68[15:0]) +
	( 16'sd 24633) * $signed(input_fmap_69[15:0]) +
	( 15'sd 12452) * $signed(input_fmap_70[15:0]) +
	( 15'sd 14899) * $signed(input_fmap_71[15:0]) +
	( 16'sd 31924) * $signed(input_fmap_72[15:0]) +
	( 12'sd 2028) * $signed(input_fmap_73[15:0]) +
	( 15'sd 11756) * $signed(input_fmap_74[15:0]) +
	( 15'sd 14448) * $signed(input_fmap_75[15:0]) +
	( 14'sd 7761) * $signed(input_fmap_76[15:0]) +
	( 15'sd 11348) * $signed(input_fmap_77[15:0]) +
	( 16'sd 18319) * $signed(input_fmap_78[15:0]) +
	( 16'sd 24068) * $signed(input_fmap_79[15:0]) +
	( 14'sd 4429) * $signed(input_fmap_80[15:0]) +
	( 16'sd 22319) * $signed(input_fmap_81[15:0]) +
	( 12'sd 2009) * $signed(input_fmap_82[15:0]) +
	( 16'sd 22229) * $signed(input_fmap_83[15:0]) +
	( 14'sd 6884) * $signed(input_fmap_84[15:0]) +
	( 16'sd 25500) * $signed(input_fmap_85[15:0]) +
	( 16'sd 23399) * $signed(input_fmap_86[15:0]) +
	( 16'sd 29090) * $signed(input_fmap_87[15:0]) +
	( 12'sd 2026) * $signed(input_fmap_88[15:0]) +
	( 16'sd 30827) * $signed(input_fmap_89[15:0]) +
	( 14'sd 4991) * $signed(input_fmap_90[15:0]) +
	( 14'sd 7592) * $signed(input_fmap_91[15:0]) +
	( 16'sd 23848) * $signed(input_fmap_92[15:0]) +
	( 13'sd 2881) * $signed(input_fmap_93[15:0]) +
	( 16'sd 29784) * $signed(input_fmap_94[15:0]) +
	( 16'sd 19766) * $signed(input_fmap_95[15:0]) +
	( 15'sd 12447) * $signed(input_fmap_96[15:0]) +
	( 16'sd 31526) * $signed(input_fmap_97[15:0]) +
	( 16'sd 32590) * $signed(input_fmap_98[15:0]) +
	( 15'sd 10632) * $signed(input_fmap_99[15:0]) +
	( 16'sd 26145) * $signed(input_fmap_100[15:0]) +
	( 15'sd 12937) * $signed(input_fmap_101[15:0]) +
	( 13'sd 3600) * $signed(input_fmap_102[15:0]) +
	( 16'sd 31019) * $signed(input_fmap_103[15:0]) +
	( 15'sd 9590) * $signed(input_fmap_104[15:0]) +
	( 16'sd 28713) * $signed(input_fmap_105[15:0]) +
	( 16'sd 17299) * $signed(input_fmap_106[15:0]) +
	( 15'sd 14033) * $signed(input_fmap_107[15:0]) +
	( 14'sd 6667) * $signed(input_fmap_108[15:0]) +
	( 16'sd 29317) * $signed(input_fmap_109[15:0]) +
	( 14'sd 6002) * $signed(input_fmap_110[15:0]) +
	( 13'sd 2664) * $signed(input_fmap_111[15:0]) +
	( 16'sd 18590) * $signed(input_fmap_112[15:0]) +
	( 14'sd 6761) * $signed(input_fmap_113[15:0]) +
	( 16'sd 17675) * $signed(input_fmap_114[15:0]) +
	( 14'sd 7065) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15239) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27004) * $signed(input_fmap_117[15:0]) +
	( 15'sd 9936) * $signed(input_fmap_118[15:0]) +
	( 15'sd 10039) * $signed(input_fmap_119[15:0]) +
	( 16'sd 28537) * $signed(input_fmap_120[15:0]) +
	( 16'sd 29847) * $signed(input_fmap_121[15:0]) +
	( 14'sd 5455) * $signed(input_fmap_122[15:0]) +
	( 15'sd 14535) * $signed(input_fmap_123[15:0]) +
	( 16'sd 21335) * $signed(input_fmap_124[15:0]) +
	( 10'sd 419) * $signed(input_fmap_125[15:0]) +
	( 16'sd 28302) * $signed(input_fmap_126[15:0]) +
	( 15'sd 15039) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 16'sd 16550) * $signed(input_fmap_0[15:0]) +
	( 15'sd 15766) * $signed(input_fmap_1[15:0]) +
	( 14'sd 7884) * $signed(input_fmap_2[15:0]) +
	( 14'sd 4765) * $signed(input_fmap_3[15:0]) +
	( 14'sd 6347) * $signed(input_fmap_4[15:0]) +
	( 16'sd 29171) * $signed(input_fmap_5[15:0]) +
	( 16'sd 29462) * $signed(input_fmap_6[15:0]) +
	( 16'sd 32703) * $signed(input_fmap_7[15:0]) +
	( 15'sd 11424) * $signed(input_fmap_8[15:0]) +
	( 16'sd 27494) * $signed(input_fmap_9[15:0]) +
	( 15'sd 11150) * $signed(input_fmap_10[15:0]) +
	( 12'sd 1127) * $signed(input_fmap_11[15:0]) +
	( 16'sd 32669) * $signed(input_fmap_12[15:0]) +
	( 15'sd 14994) * $signed(input_fmap_13[15:0]) +
	( 15'sd 14484) * $signed(input_fmap_14[15:0]) +
	( 15'sd 9234) * $signed(input_fmap_15[15:0]) +
	( 16'sd 28409) * $signed(input_fmap_16[15:0]) +
	( 16'sd 30993) * $signed(input_fmap_17[15:0]) +
	( 16'sd 29153) * $signed(input_fmap_18[15:0]) +
	( 14'sd 4750) * $signed(input_fmap_19[15:0]) +
	( 15'sd 9870) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17505) * $signed(input_fmap_21[15:0]) +
	( 14'sd 8133) * $signed(input_fmap_22[15:0]) +
	( 16'sd 30162) * $signed(input_fmap_23[15:0]) +
	( 15'sd 10180) * $signed(input_fmap_24[15:0]) +
	( 16'sd 26944) * $signed(input_fmap_25[15:0]) +
	( 16'sd 27288) * $signed(input_fmap_26[15:0]) +
	( 16'sd 19313) * $signed(input_fmap_27[15:0]) +
	( 16'sd 17298) * $signed(input_fmap_28[15:0]) +
	( 15'sd 13970) * $signed(input_fmap_29[15:0]) +
	( 15'sd 9968) * $signed(input_fmap_30[15:0]) +
	( 15'sd 12651) * $signed(input_fmap_31[15:0]) +
	( 15'sd 11528) * $signed(input_fmap_32[15:0]) +
	( 16'sd 23240) * $signed(input_fmap_33[15:0]) +
	( 16'sd 32268) * $signed(input_fmap_34[15:0]) +
	( 15'sd 14936) * $signed(input_fmap_35[15:0]) +
	( 16'sd 19897) * $signed(input_fmap_36[15:0]) +
	( 16'sd 30438) * $signed(input_fmap_37[15:0]) +
	( 16'sd 31650) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24269) * $signed(input_fmap_39[15:0]) +
	( 14'sd 6455) * $signed(input_fmap_40[15:0]) +
	( 15'sd 11330) * $signed(input_fmap_41[15:0]) +
	( 14'sd 5618) * $signed(input_fmap_42[15:0]) +
	( 16'sd 29098) * $signed(input_fmap_43[15:0]) +
	( 12'sd 1272) * $signed(input_fmap_44[15:0]) +
	( 13'sd 4040) * $signed(input_fmap_45[15:0]) +
	( 16'sd 23182) * $signed(input_fmap_46[15:0]) +
	( 15'sd 12165) * $signed(input_fmap_47[15:0]) +
	( 15'sd 14263) * $signed(input_fmap_48[15:0]) +
	( 14'sd 4221) * $signed(input_fmap_49[15:0]) +
	( 13'sd 3492) * $signed(input_fmap_50[15:0]) +
	( 16'sd 24944) * $signed(input_fmap_51[15:0]) +
	( 14'sd 4970) * $signed(input_fmap_52[15:0]) +
	( 14'sd 6955) * $signed(input_fmap_53[15:0]) +
	( 16'sd 20034) * $signed(input_fmap_54[15:0]) +
	( 16'sd 18846) * $signed(input_fmap_55[15:0]) +
	( 16'sd 17232) * $signed(input_fmap_56[15:0]) +
	( 13'sd 2717) * $signed(input_fmap_57[15:0]) +
	( 11'sd 586) * $signed(input_fmap_58[15:0]) +
	( 16'sd 23113) * $signed(input_fmap_59[15:0]) +
	( 16'sd 16817) * $signed(input_fmap_60[15:0]) +
	( 15'sd 14857) * $signed(input_fmap_61[15:0]) +
	( 16'sd 16709) * $signed(input_fmap_62[15:0]) +
	( 16'sd 23044) * $signed(input_fmap_63[15:0]) +
	( 16'sd 31923) * $signed(input_fmap_64[15:0]) +
	( 16'sd 27169) * $signed(input_fmap_65[15:0]) +
	( 16'sd 30927) * $signed(input_fmap_66[15:0]) +
	( 10'sd 414) * $signed(input_fmap_67[15:0]) +
	( 16'sd 25520) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31575) * $signed(input_fmap_69[15:0]) +
	( 13'sd 4091) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31686) * $signed(input_fmap_71[15:0]) +
	( 13'sd 2393) * $signed(input_fmap_72[15:0]) +
	( 15'sd 15630) * $signed(input_fmap_73[15:0]) +
	( 16'sd 30691) * $signed(input_fmap_74[15:0]) +
	( 15'sd 9906) * $signed(input_fmap_75[15:0]) +
	( 14'sd 8158) * $signed(input_fmap_76[15:0]) +
	( 15'sd 8554) * $signed(input_fmap_77[15:0]) +
	( 16'sd 32694) * $signed(input_fmap_78[15:0]) +
	( 14'sd 6819) * $signed(input_fmap_79[15:0]) +
	( 14'sd 4275) * $signed(input_fmap_80[15:0]) +
	( 15'sd 16212) * $signed(input_fmap_81[15:0]) +
	( 15'sd 9666) * $signed(input_fmap_82[15:0]) +
	( 14'sd 7975) * $signed(input_fmap_83[15:0]) +
	( 12'sd 1222) * $signed(input_fmap_84[15:0]) +
	( 14'sd 5617) * $signed(input_fmap_85[15:0]) +
	( 14'sd 7366) * $signed(input_fmap_86[15:0]) +
	( 15'sd 12316) * $signed(input_fmap_87[15:0]) +
	( 15'sd 8524) * $signed(input_fmap_88[15:0]) +
	( 16'sd 26571) * $signed(input_fmap_89[15:0]) +
	( 16'sd 27846) * $signed(input_fmap_90[15:0]) +
	( 16'sd 17992) * $signed(input_fmap_91[15:0]) +
	( 16'sd 28369) * $signed(input_fmap_92[15:0]) +
	( 16'sd 29352) * $signed(input_fmap_93[15:0]) +
	( 16'sd 27135) * $signed(input_fmap_94[15:0]) +
	( 16'sd 22708) * $signed(input_fmap_95[15:0]) +
	( 15'sd 9313) * $signed(input_fmap_96[15:0]) +
	( 16'sd 28911) * $signed(input_fmap_97[15:0]) +
	( 15'sd 14295) * $signed(input_fmap_98[15:0]) +
	( 16'sd 26621) * $signed(input_fmap_99[15:0]) +
	( 15'sd 14281) * $signed(input_fmap_100[15:0]) +
	( 15'sd 11915) * $signed(input_fmap_101[15:0]) +
	( 12'sd 1586) * $signed(input_fmap_102[15:0]) +
	( 12'sd 1084) * $signed(input_fmap_103[15:0]) +
	( 16'sd 17238) * $signed(input_fmap_104[15:0]) +
	( 16'sd 26810) * $signed(input_fmap_105[15:0]) +
	( 14'sd 5263) * $signed(input_fmap_106[15:0]) +
	( 15'sd 14760) * $signed(input_fmap_107[15:0]) +
	( 15'sd 14885) * $signed(input_fmap_108[15:0]) +
	( 14'sd 7796) * $signed(input_fmap_109[15:0]) +
	( 16'sd 31919) * $signed(input_fmap_110[15:0]) +
	( 12'sd 1966) * $signed(input_fmap_111[15:0]) +
	( 15'sd 15158) * $signed(input_fmap_112[15:0]) +
	( 14'sd 4630) * $signed(input_fmap_113[15:0]) +
	( 16'sd 21268) * $signed(input_fmap_114[15:0]) +
	( 16'sd 27950) * $signed(input_fmap_115[15:0]) +
	( 15'sd 9231) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27446) * $signed(input_fmap_117[15:0]) +
	( 13'sd 3905) * $signed(input_fmap_118[15:0]) +
	( 12'sd 1331) * $signed(input_fmap_119[15:0]) +
	( 16'sd 26664) * $signed(input_fmap_120[15:0]) +
	( 15'sd 14878) * $signed(input_fmap_121[15:0]) +
	( 16'sd 28482) * $signed(input_fmap_122[15:0]) +
	( 16'sd 29325) * $signed(input_fmap_123[15:0]) +
	( 13'sd 3086) * $signed(input_fmap_124[15:0]) +
	( 16'sd 30673) * $signed(input_fmap_125[15:0]) +
	( 15'sd 9794) * $signed(input_fmap_126[15:0]) +
	( 14'sd 8132) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 16'sd 21193) * $signed(input_fmap_0[15:0]) +
	( 16'sd 16626) * $signed(input_fmap_1[15:0]) +
	( 16'sd 28928) * $signed(input_fmap_2[15:0]) +
	( 14'sd 5293) * $signed(input_fmap_3[15:0]) +
	( 15'sd 15077) * $signed(input_fmap_4[15:0]) +
	( 12'sd 1888) * $signed(input_fmap_5[15:0]) +
	( 16'sd 22069) * $signed(input_fmap_6[15:0]) +
	( 16'sd 20061) * $signed(input_fmap_7[15:0]) +
	( 15'sd 13809) * $signed(input_fmap_8[15:0]) +
	( 16'sd 22280) * $signed(input_fmap_9[15:0]) +
	( 14'sd 4389) * $signed(input_fmap_10[15:0]) +
	( 14'sd 6598) * $signed(input_fmap_11[15:0]) +
	( 15'sd 15691) * $signed(input_fmap_12[15:0]) +
	( 15'sd 14239) * $signed(input_fmap_13[15:0]) +
	( 16'sd 23890) * $signed(input_fmap_14[15:0]) +
	( 16'sd 18504) * $signed(input_fmap_15[15:0]) +
	( 16'sd 32011) * $signed(input_fmap_16[15:0]) +
	( 14'sd 6993) * $signed(input_fmap_17[15:0]) +
	( 16'sd 30793) * $signed(input_fmap_18[15:0]) +
	( 16'sd 18970) * $signed(input_fmap_19[15:0]) +
	( 16'sd 23533) * $signed(input_fmap_20[15:0]) +
	( 12'sd 1540) * $signed(input_fmap_21[15:0]) +
	( 16'sd 30775) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24929) * $signed(input_fmap_23[15:0]) +
	( 15'sd 11790) * $signed(input_fmap_24[15:0]) +
	( 16'sd 26488) * $signed(input_fmap_25[15:0]) +
	( 14'sd 4569) * $signed(input_fmap_26[15:0]) +
	( 15'sd 12749) * $signed(input_fmap_27[15:0]) +
	( 16'sd 32055) * $signed(input_fmap_28[15:0]) +
	( 16'sd 17217) * $signed(input_fmap_29[15:0]) +
	( 16'sd 25172) * $signed(input_fmap_30[15:0]) +
	( 14'sd 5095) * $signed(input_fmap_31[15:0]) +
	( 16'sd 23491) * $signed(input_fmap_32[15:0]) +
	( 16'sd 27518) * $signed(input_fmap_33[15:0]) +
	( 13'sd 3053) * $signed(input_fmap_34[15:0]) +
	( 15'sd 11075) * $signed(input_fmap_35[15:0]) +
	( 16'sd 26967) * $signed(input_fmap_36[15:0]) +
	( 16'sd 31131) * $signed(input_fmap_37[15:0]) +
	( 12'sd 1972) * $signed(input_fmap_38[15:0]) +
	( 16'sd 26798) * $signed(input_fmap_39[15:0]) +
	( 16'sd 20710) * $signed(input_fmap_40[15:0]) +
	( 16'sd 16992) * $signed(input_fmap_41[15:0]) +
	( 15'sd 15593) * $signed(input_fmap_42[15:0]) +
	( 16'sd 16645) * $signed(input_fmap_43[15:0]) +
	( 15'sd 9303) * $signed(input_fmap_44[15:0]) +
	( 16'sd 26679) * $signed(input_fmap_45[15:0]) +
	( 12'sd 1872) * $signed(input_fmap_46[15:0]) +
	( 16'sd 22739) * $signed(input_fmap_47[15:0]) +
	( 16'sd 17109) * $signed(input_fmap_48[15:0]) +
	( 16'sd 22803) * $signed(input_fmap_49[15:0]) +
	( 15'sd 11512) * $signed(input_fmap_50[15:0]) +
	( 15'sd 11705) * $signed(input_fmap_51[15:0]) +
	( 16'sd 30053) * $signed(input_fmap_52[15:0]) +
	( 16'sd 27742) * $signed(input_fmap_53[15:0]) +
	( 16'sd 18162) * $signed(input_fmap_54[15:0]) +
	( 16'sd 19760) * $signed(input_fmap_55[15:0]) +
	( 15'sd 12383) * $signed(input_fmap_56[15:0]) +
	( 16'sd 29877) * $signed(input_fmap_57[15:0]) +
	( 14'sd 7975) * $signed(input_fmap_58[15:0]) +
	( 14'sd 4218) * $signed(input_fmap_59[15:0]) +
	( 16'sd 16392) * $signed(input_fmap_60[15:0]) +
	( 10'sd 469) * $signed(input_fmap_61[15:0]) +
	( 15'sd 12150) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20896) * $signed(input_fmap_63[15:0]) +
	( 16'sd 16496) * $signed(input_fmap_64[15:0]) +
	( 14'sd 7395) * $signed(input_fmap_65[15:0]) +
	( 14'sd 7288) * $signed(input_fmap_66[15:0]) +
	( 16'sd 25662) * $signed(input_fmap_67[15:0]) +
	( 15'sd 11470) * $signed(input_fmap_68[15:0]) +
	( 16'sd 32329) * $signed(input_fmap_69[15:0]) +
	( 16'sd 20222) * $signed(input_fmap_70[15:0]) +
	( 15'sd 8412) * $signed(input_fmap_71[15:0]) +
	( 16'sd 32001) * $signed(input_fmap_72[15:0]) +
	( 16'sd 30840) * $signed(input_fmap_73[15:0]) +
	( 16'sd 21462) * $signed(input_fmap_74[15:0]) +
	( 15'sd 11582) * $signed(input_fmap_75[15:0]) +
	( 12'sd 1756) * $signed(input_fmap_76[15:0]) +
	( 13'sd 3854) * $signed(input_fmap_77[15:0]) +
	( 16'sd 20147) * $signed(input_fmap_78[15:0]) +
	( 15'sd 11294) * $signed(input_fmap_79[15:0]) +
	( 16'sd 30451) * $signed(input_fmap_80[15:0]) +
	( 15'sd 13657) * $signed(input_fmap_81[15:0]) +
	( 16'sd 16787) * $signed(input_fmap_82[15:0]) +
	( 16'sd 22617) * $signed(input_fmap_83[15:0]) +
	( 13'sd 2293) * $signed(input_fmap_84[15:0]) +
	( 12'sd 1884) * $signed(input_fmap_85[15:0]) +
	( 16'sd 24183) * $signed(input_fmap_86[15:0]) +
	( 16'sd 26132) * $signed(input_fmap_87[15:0]) +
	( 11'sd 530) * $signed(input_fmap_88[15:0]) +
	( 16'sd 31427) * $signed(input_fmap_89[15:0]) +
	( 15'sd 15063) * $signed(input_fmap_90[15:0]) +
	( 15'sd 15153) * $signed(input_fmap_91[15:0]) +
	( 13'sd 2444) * $signed(input_fmap_92[15:0]) +
	( 15'sd 9497) * $signed(input_fmap_93[15:0]) +
	( 15'sd 10788) * $signed(input_fmap_94[15:0]) +
	( 14'sd 8131) * $signed(input_fmap_95[15:0]) +
	( 16'sd 32244) * $signed(input_fmap_96[15:0]) +
	( 15'sd 15610) * $signed(input_fmap_97[15:0]) +
	( 16'sd 24971) * $signed(input_fmap_98[15:0]) +
	( 14'sd 7962) * $signed(input_fmap_99[15:0]) +
	( 15'sd 11058) * $signed(input_fmap_100[15:0]) +
	( 15'sd 14832) * $signed(input_fmap_101[15:0]) +
	( 15'sd 12555) * $signed(input_fmap_102[15:0]) +
	( 14'sd 6344) * $signed(input_fmap_103[15:0]) +
	( 15'sd 8964) * $signed(input_fmap_104[15:0]) +
	( 15'sd 13666) * $signed(input_fmap_105[15:0]) +
	( 16'sd 16955) * $signed(input_fmap_106[15:0]) +
	( 11'sd 611) * $signed(input_fmap_107[15:0]) +
	( 11'sd 580) * $signed(input_fmap_108[15:0]) +
	( 15'sd 9790) * $signed(input_fmap_109[15:0]) +
	( 15'sd 12757) * $signed(input_fmap_110[15:0]) +
	( 16'sd 24339) * $signed(input_fmap_111[15:0]) +
	( 16'sd 23415) * $signed(input_fmap_112[15:0]) +
	( 16'sd 26671) * $signed(input_fmap_113[15:0]) +
	( 16'sd 22525) * $signed(input_fmap_114[15:0]) +
	( 16'sd 18366) * $signed(input_fmap_115[15:0]) +
	( 15'sd 14384) * $signed(input_fmap_116[15:0]) +
	( 16'sd 32168) * $signed(input_fmap_117[15:0]) +
	( 14'sd 4200) * $signed(input_fmap_118[15:0]) +
	( 15'sd 13189) * $signed(input_fmap_119[15:0]) +
	( 16'sd 16987) * $signed(input_fmap_120[15:0]) +
	( 15'sd 13413) * $signed(input_fmap_121[15:0]) +
	( 16'sd 17503) * $signed(input_fmap_122[15:0]) +
	( 16'sd 24520) * $signed(input_fmap_123[15:0]) +
	( 14'sd 6455) * $signed(input_fmap_124[15:0]) +
	( 15'sd 8425) * $signed(input_fmap_125[15:0]) +
	( 12'sd 1255) * $signed(input_fmap_126[15:0]) +
	( 15'sd 14142) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 14'sd 5001) * $signed(input_fmap_0[15:0]) +
	( 14'sd 7205) * $signed(input_fmap_1[15:0]) +
	( 12'sd 1441) * $signed(input_fmap_2[15:0]) +
	( 14'sd 4360) * $signed(input_fmap_3[15:0]) +
	( 14'sd 5358) * $signed(input_fmap_4[15:0]) +
	( 16'sd 24230) * $signed(input_fmap_5[15:0]) +
	( 13'sd 3194) * $signed(input_fmap_6[15:0]) +
	( 15'sd 10685) * $signed(input_fmap_7[15:0]) +
	( 15'sd 12700) * $signed(input_fmap_8[15:0]) +
	( 12'sd 1458) * $signed(input_fmap_9[15:0]) +
	( 15'sd 15236) * $signed(input_fmap_10[15:0]) +
	( 16'sd 25192) * $signed(input_fmap_11[15:0]) +
	( 16'sd 19854) * $signed(input_fmap_12[15:0]) +
	( 16'sd 28970) * $signed(input_fmap_13[15:0]) +
	( 15'sd 12129) * $signed(input_fmap_14[15:0]) +
	( 14'sd 7967) * $signed(input_fmap_15[15:0]) +
	( 15'sd 8560) * $signed(input_fmap_16[15:0]) +
	( 15'sd 12831) * $signed(input_fmap_17[15:0]) +
	( 12'sd 1614) * $signed(input_fmap_18[15:0]) +
	( 15'sd 14273) * $signed(input_fmap_19[15:0]) +
	( 16'sd 31351) * $signed(input_fmap_20[15:0]) +
	( 16'sd 18747) * $signed(input_fmap_21[15:0]) +
	( 13'sd 3331) * $signed(input_fmap_22[15:0]) +
	( 16'sd 30482) * $signed(input_fmap_23[15:0]) +
	( 15'sd 8540) * $signed(input_fmap_24[15:0]) +
	( 13'sd 2144) * $signed(input_fmap_25[15:0]) +
	( 16'sd 29361) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2143) * $signed(input_fmap_27[15:0]) +
	( 16'sd 18740) * $signed(input_fmap_28[15:0]) +
	( 16'sd 25711) * $signed(input_fmap_29[15:0]) +
	( 16'sd 26902) * $signed(input_fmap_30[15:0]) +
	( 16'sd 18758) * $signed(input_fmap_31[15:0]) +
	( 14'sd 4574) * $signed(input_fmap_32[15:0]) +
	( 16'sd 28184) * $signed(input_fmap_33[15:0]) +
	( 15'sd 11932) * $signed(input_fmap_34[15:0]) +
	( 14'sd 4377) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2126) * $signed(input_fmap_36[15:0]) +
	( 15'sd 15135) * $signed(input_fmap_37[15:0]) +
	( 16'sd 29952) * $signed(input_fmap_38[15:0]) +
	( 14'sd 5079) * $signed(input_fmap_39[15:0]) +
	( 16'sd 21695) * $signed(input_fmap_40[15:0]) +
	( 16'sd 19839) * $signed(input_fmap_41[15:0]) +
	( 14'sd 5563) * $signed(input_fmap_42[15:0]) +
	( 15'sd 13040) * $signed(input_fmap_43[15:0]) +
	( 14'sd 7324) * $signed(input_fmap_44[15:0]) +
	( 13'sd 2963) * $signed(input_fmap_45[15:0]) +
	( 16'sd 30456) * $signed(input_fmap_46[15:0]) +
	( 14'sd 7905) * $signed(input_fmap_47[15:0]) +
	( 16'sd 20117) * $signed(input_fmap_48[15:0]) +
	( 15'sd 13607) * $signed(input_fmap_49[15:0]) +
	( 16'sd 19664) * $signed(input_fmap_50[15:0]) +
	( 16'sd 24945) * $signed(input_fmap_51[15:0]) +
	( 16'sd 17782) * $signed(input_fmap_52[15:0]) +
	( 15'sd 13366) * $signed(input_fmap_53[15:0]) +
	( 14'sd 4847) * $signed(input_fmap_54[15:0]) +
	( 16'sd 27722) * $signed(input_fmap_55[15:0]) +
	( 16'sd 31093) * $signed(input_fmap_56[15:0]) +
	( 15'sd 10897) * $signed(input_fmap_57[15:0]) +
	( 13'sd 3809) * $signed(input_fmap_58[15:0]) +
	( 16'sd 25869) * $signed(input_fmap_59[15:0]) +
	( 16'sd 25504) * $signed(input_fmap_60[15:0]) +
	( 13'sd 2351) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29359) * $signed(input_fmap_62[15:0]) +
	( 14'sd 6585) * $signed(input_fmap_63[15:0]) +
	( 16'sd 30641) * $signed(input_fmap_64[15:0]) +
	( 14'sd 4583) * $signed(input_fmap_65[15:0]) +
	( 12'sd 1895) * $signed(input_fmap_66[15:0]) +
	( 15'sd 16229) * $signed(input_fmap_67[15:0]) +
	( 13'sd 2600) * $signed(input_fmap_68[15:0]) +
	( 12'sd 1579) * $signed(input_fmap_69[15:0]) +
	( 12'sd 1595) * $signed(input_fmap_70[15:0]) +
	( 16'sd 16705) * $signed(input_fmap_71[15:0]) +
	( 16'sd 28300) * $signed(input_fmap_72[15:0]) +
	( 16'sd 28850) * $signed(input_fmap_73[15:0]) +
	( 16'sd 32744) * $signed(input_fmap_74[15:0]) +
	( 16'sd 28494) * $signed(input_fmap_75[15:0]) +
	( 16'sd 17090) * $signed(input_fmap_76[15:0]) +
	( 16'sd 28469) * $signed(input_fmap_77[15:0]) +
	( 16'sd 21428) * $signed(input_fmap_78[15:0]) +
	( 12'sd 1330) * $signed(input_fmap_79[15:0]) +
	( 16'sd 29310) * $signed(input_fmap_80[15:0]) +
	( 15'sd 14242) * $signed(input_fmap_81[15:0]) +
	( 16'sd 21119) * $signed(input_fmap_82[15:0]) +
	( 15'sd 12259) * $signed(input_fmap_83[15:0]) +
	( 15'sd 8380) * $signed(input_fmap_84[15:0]) +
	( 16'sd 18197) * $signed(input_fmap_85[15:0]) +
	( 15'sd 10307) * $signed(input_fmap_86[15:0]) +
	( 16'sd 25801) * $signed(input_fmap_87[15:0]) +
	( 15'sd 13116) * $signed(input_fmap_88[15:0]) +
	( 15'sd 13126) * $signed(input_fmap_89[15:0]) +
	( 15'sd 15323) * $signed(input_fmap_90[15:0]) +
	( 16'sd 29801) * $signed(input_fmap_91[15:0]) +
	( 16'sd 23154) * $signed(input_fmap_92[15:0]) +
	( 16'sd 28978) * $signed(input_fmap_93[15:0]) +
	( 16'sd 28844) * $signed(input_fmap_94[15:0]) +
	( 13'sd 2373) * $signed(input_fmap_95[15:0]) +
	( 15'sd 10187) * $signed(input_fmap_96[15:0]) +
	( 15'sd 13754) * $signed(input_fmap_97[15:0]) +
	( 8'sd 89) * $signed(input_fmap_98[15:0]) +
	( 15'sd 12837) * $signed(input_fmap_99[15:0]) +
	( 16'sd 27577) * $signed(input_fmap_100[15:0]) +
	( 16'sd 22294) * $signed(input_fmap_101[15:0]) +
	( 15'sd 10519) * $signed(input_fmap_102[15:0]) +
	( 16'sd 29574) * $signed(input_fmap_103[15:0]) +
	( 14'sd 5724) * $signed(input_fmap_104[15:0]) +
	( 15'sd 13898) * $signed(input_fmap_105[15:0]) +
	( 16'sd 21058) * $signed(input_fmap_106[15:0]) +
	( 16'sd 24219) * $signed(input_fmap_107[15:0]) +
	( 16'sd 16652) * $signed(input_fmap_108[15:0]) +
	( 16'sd 27570) * $signed(input_fmap_109[15:0]) +
	( 14'sd 5355) * $signed(input_fmap_110[15:0]) +
	( 11'sd 648) * $signed(input_fmap_111[15:0]) +
	( 16'sd 28061) * $signed(input_fmap_112[15:0]) +
	( 15'sd 14410) * $signed(input_fmap_113[15:0]) +
	( 15'sd 16224) * $signed(input_fmap_114[15:0]) +
	( 15'sd 13025) * $signed(input_fmap_115[15:0]) +
	( 14'sd 7504) * $signed(input_fmap_116[15:0]) +
	( 9'sd 235) * $signed(input_fmap_117[15:0]) +
	( 16'sd 28315) * $signed(input_fmap_118[15:0]) +
	( 16'sd 22697) * $signed(input_fmap_119[15:0]) +
	( 15'sd 9259) * $signed(input_fmap_120[15:0]) +
	( 15'sd 13857) * $signed(input_fmap_121[15:0]) +
	( 16'sd 24442) * $signed(input_fmap_122[15:0]) +
	( 14'sd 5232) * $signed(input_fmap_123[15:0]) +
	( 14'sd 4902) * $signed(input_fmap_124[15:0]) +
	( 16'sd 25326) * $signed(input_fmap_125[15:0]) +
	( 16'sd 23790) * $signed(input_fmap_126[15:0]) +
	( 15'sd 10820) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 16'sd 21898) * $signed(input_fmap_0[15:0]) +
	( 16'sd 20342) * $signed(input_fmap_1[15:0]) +
	( 16'sd 17850) * $signed(input_fmap_2[15:0]) +
	( 16'sd 30495) * $signed(input_fmap_3[15:0]) +
	( 16'sd 17389) * $signed(input_fmap_4[15:0]) +
	( 13'sd 3780) * $signed(input_fmap_5[15:0]) +
	( 10'sd 444) * $signed(input_fmap_6[15:0]) +
	( 16'sd 16699) * $signed(input_fmap_7[15:0]) +
	( 16'sd 20431) * $signed(input_fmap_8[15:0]) +
	( 15'sd 14498) * $signed(input_fmap_9[15:0]) +
	( 15'sd 12724) * $signed(input_fmap_10[15:0]) +
	( 16'sd 24610) * $signed(input_fmap_11[15:0]) +
	( 16'sd 24812) * $signed(input_fmap_12[15:0]) +
	( 13'sd 2520) * $signed(input_fmap_13[15:0]) +
	( 16'sd 25602) * $signed(input_fmap_14[15:0]) +
	( 13'sd 3858) * $signed(input_fmap_15[15:0]) +
	( 16'sd 20064) * $signed(input_fmap_16[15:0]) +
	( 16'sd 31900) * $signed(input_fmap_17[15:0]) +
	( 14'sd 8045) * $signed(input_fmap_18[15:0]) +
	( 15'sd 15917) * $signed(input_fmap_19[15:0]) +
	( 16'sd 27353) * $signed(input_fmap_20[15:0]) +
	( 13'sd 3238) * $signed(input_fmap_21[15:0]) +
	( 13'sd 3016) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28381) * $signed(input_fmap_23[15:0]) +
	( 14'sd 5801) * $signed(input_fmap_24[15:0]) +
	( 15'sd 15063) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22756) * $signed(input_fmap_26[15:0]) +
	( 16'sd 25770) * $signed(input_fmap_27[15:0]) +
	( 16'sd 27568) * $signed(input_fmap_28[15:0]) +
	( 16'sd 27288) * $signed(input_fmap_29[15:0]) +
	( 15'sd 10591) * $signed(input_fmap_30[15:0]) +
	( 16'sd 24044) * $signed(input_fmap_31[15:0]) +
	( 15'sd 9695) * $signed(input_fmap_32[15:0]) +
	( 16'sd 28791) * $signed(input_fmap_33[15:0]) +
	( 16'sd 32378) * $signed(input_fmap_34[15:0]) +
	( 16'sd 19506) * $signed(input_fmap_35[15:0]) +
	( 15'sd 14391) * $signed(input_fmap_36[15:0]) +
	( 15'sd 9681) * $signed(input_fmap_37[15:0]) +
	( 16'sd 16687) * $signed(input_fmap_38[15:0]) +
	( 13'sd 3850) * $signed(input_fmap_39[15:0]) +
	( 13'sd 2458) * $signed(input_fmap_40[15:0]) +
	( 12'sd 1281) * $signed(input_fmap_41[15:0]) +
	( 15'sd 12169) * $signed(input_fmap_42[15:0]) +
	( 16'sd 29581) * $signed(input_fmap_43[15:0]) +
	( 14'sd 5629) * $signed(input_fmap_44[15:0]) +
	( 14'sd 6720) * $signed(input_fmap_45[15:0]) +
	( 14'sd 7662) * $signed(input_fmap_46[15:0]) +
	( 16'sd 16746) * $signed(input_fmap_47[15:0]) +
	( 16'sd 22851) * $signed(input_fmap_48[15:0]) +
	( 16'sd 31018) * $signed(input_fmap_49[15:0]) +
	( 16'sd 25806) * $signed(input_fmap_50[15:0]) +
	( 15'sd 16011) * $signed(input_fmap_51[15:0]) +
	( 16'sd 22820) * $signed(input_fmap_52[15:0]) +
	( 12'sd 1030) * $signed(input_fmap_53[15:0]) +
	( 14'sd 5275) * $signed(input_fmap_54[15:0]) +
	( 15'sd 11981) * $signed(input_fmap_55[15:0]) +
	( 16'sd 32691) * $signed(input_fmap_56[15:0]) +
	( 15'sd 8801) * $signed(input_fmap_57[15:0]) +
	( 15'sd 12114) * $signed(input_fmap_58[15:0]) +
	( 15'sd 13083) * $signed(input_fmap_59[15:0]) +
	( 16'sd 22157) * $signed(input_fmap_60[15:0]) +
	( 15'sd 14603) * $signed(input_fmap_61[15:0]) +
	( 15'sd 9353) * $signed(input_fmap_62[15:0]) +
	( 14'sd 7145) * $signed(input_fmap_63[15:0]) +
	( 16'sd 18795) * $signed(input_fmap_64[15:0]) +
	( 14'sd 7106) * $signed(input_fmap_65[15:0]) +
	( 13'sd 3984) * $signed(input_fmap_66[15:0]) +
	( 15'sd 9126) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26818) * $signed(input_fmap_68[15:0]) +
	( 13'sd 2366) * $signed(input_fmap_69[15:0]) +
	( 16'sd 23957) * $signed(input_fmap_70[15:0]) +
	( 16'sd 28240) * $signed(input_fmap_71[15:0]) +
	( 16'sd 17527) * $signed(input_fmap_72[15:0]) +
	( 14'sd 5110) * $signed(input_fmap_73[15:0]) +
	( 15'sd 12261) * $signed(input_fmap_74[15:0]) +
	( 16'sd 23021) * $signed(input_fmap_75[15:0]) +
	( 15'sd 12458) * $signed(input_fmap_76[15:0]) +
	( 15'sd 12390) * $signed(input_fmap_77[15:0]) +
	( 15'sd 12421) * $signed(input_fmap_78[15:0]) +
	( 15'sd 13836) * $signed(input_fmap_79[15:0]) +
	( 15'sd 8683) * $signed(input_fmap_80[15:0]) +
	( 16'sd 17257) * $signed(input_fmap_81[15:0]) +
	( 16'sd 21288) * $signed(input_fmap_82[15:0]) +
	( 15'sd 10045) * $signed(input_fmap_83[15:0]) +
	( 13'sd 2114) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24945) * $signed(input_fmap_85[15:0]) +
	( 15'sd 11777) * $signed(input_fmap_86[15:0]) +
	( 16'sd 26252) * $signed(input_fmap_87[15:0]) +
	( 16'sd 30957) * $signed(input_fmap_88[15:0]) +
	( 16'sd 23904) * $signed(input_fmap_89[15:0]) +
	( 15'sd 9983) * $signed(input_fmap_90[15:0]) +
	( 16'sd 27448) * $signed(input_fmap_91[15:0]) +
	( 16'sd 26544) * $signed(input_fmap_92[15:0]) +
	( 15'sd 15290) * $signed(input_fmap_93[15:0]) +
	( 16'sd 25667) * $signed(input_fmap_94[15:0]) +
	( 14'sd 6961) * $signed(input_fmap_95[15:0]) +
	( 15'sd 11911) * $signed(input_fmap_96[15:0]) +
	( 16'sd 17444) * $signed(input_fmap_97[15:0]) +
	( 15'sd 12716) * $signed(input_fmap_98[15:0]) +
	( 16'sd 24179) * $signed(input_fmap_99[15:0]) +
	( 15'sd 15352) * $signed(input_fmap_100[15:0]) +
	( 16'sd 21131) * $signed(input_fmap_101[15:0]) +
	( 12'sd 1338) * $signed(input_fmap_102[15:0]) +
	( 16'sd 18926) * $signed(input_fmap_103[15:0]) +
	( 16'sd 26634) * $signed(input_fmap_104[15:0]) +
	( 16'sd 18943) * $signed(input_fmap_105[15:0]) +
	( 16'sd 28666) * $signed(input_fmap_106[15:0]) +
	( 16'sd 20225) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15022) * $signed(input_fmap_108[15:0]) +
	( 16'sd 16666) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22896) * $signed(input_fmap_110[15:0]) +
	( 13'sd 3063) * $signed(input_fmap_111[15:0]) +
	( 14'sd 5098) * $signed(input_fmap_112[15:0]) +
	( 16'sd 23124) * $signed(input_fmap_113[15:0]) +
	( 15'sd 14641) * $signed(input_fmap_114[15:0]) +
	( 13'sd 3126) * $signed(input_fmap_115[15:0]) +
	( 16'sd 17020) * $signed(input_fmap_116[15:0]) +
	( 16'sd 22303) * $signed(input_fmap_117[15:0]) +
	( 16'sd 17236) * $signed(input_fmap_118[15:0]) +
	( 16'sd 26927) * $signed(input_fmap_119[15:0]) +
	( 16'sd 19874) * $signed(input_fmap_120[15:0]) +
	( 16'sd 21455) * $signed(input_fmap_121[15:0]) +
	( 15'sd 14550) * $signed(input_fmap_122[15:0]) +
	( 15'sd 14230) * $signed(input_fmap_123[15:0]) +
	( 15'sd 14757) * $signed(input_fmap_124[15:0]) +
	( 14'sd 5394) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6882) * $signed(input_fmap_126[15:0]) +
	( 14'sd 7878) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 15'sd 8255) * $signed(input_fmap_0[15:0]) +
	( 16'sd 18222) * $signed(input_fmap_1[15:0]) +
	( 16'sd 16716) * $signed(input_fmap_2[15:0]) +
	( 16'sd 30170) * $signed(input_fmap_3[15:0]) +
	( 13'sd 3601) * $signed(input_fmap_4[15:0]) +
	( 15'sd 16376) * $signed(input_fmap_5[15:0]) +
	( 15'sd 13532) * $signed(input_fmap_6[15:0]) +
	( 16'sd 31209) * $signed(input_fmap_7[15:0]) +
	( 15'sd 13261) * $signed(input_fmap_8[15:0]) +
	( 15'sd 8681) * $signed(input_fmap_9[15:0]) +
	( 13'sd 2674) * $signed(input_fmap_10[15:0]) +
	( 15'sd 8910) * $signed(input_fmap_11[15:0]) +
	( 16'sd 22105) * $signed(input_fmap_12[15:0]) +
	( 16'sd 26114) * $signed(input_fmap_13[15:0]) +
	( 16'sd 28897) * $signed(input_fmap_14[15:0]) +
	( 15'sd 8195) * $signed(input_fmap_15[15:0]) +
	( 14'sd 6451) * $signed(input_fmap_16[15:0]) +
	( 16'sd 19055) * $signed(input_fmap_17[15:0]) +
	( 16'sd 27703) * $signed(input_fmap_18[15:0]) +
	( 13'sd 2584) * $signed(input_fmap_19[15:0]) +
	( 16'sd 24745) * $signed(input_fmap_20[15:0]) +
	( 16'sd 30550) * $signed(input_fmap_21[15:0]) +
	( 16'sd 29252) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28986) * $signed(input_fmap_23[15:0]) +
	( 16'sd 26820) * $signed(input_fmap_24[15:0]) +
	( 15'sd 11226) * $signed(input_fmap_25[15:0]) +
	( 15'sd 14335) * $signed(input_fmap_26[15:0]) +
	( 16'sd 17560) * $signed(input_fmap_27[15:0]) +
	( 15'sd 9458) * $signed(input_fmap_28[15:0]) +
	( 16'sd 24167) * $signed(input_fmap_29[15:0]) +
	( 16'sd 17445) * $signed(input_fmap_30[15:0]) +
	( 16'sd 31963) * $signed(input_fmap_31[15:0]) +
	( 16'sd 26886) * $signed(input_fmap_32[15:0]) +
	( 14'sd 6397) * $signed(input_fmap_33[15:0]) +
	( 15'sd 13727) * $signed(input_fmap_34[15:0]) +
	( 16'sd 27534) * $signed(input_fmap_35[15:0]) +
	( 15'sd 12691) * $signed(input_fmap_36[15:0]) +
	( 15'sd 10656) * $signed(input_fmap_37[15:0]) +
	( 16'sd 27137) * $signed(input_fmap_38[15:0]) +
	( 15'sd 9921) * $signed(input_fmap_39[15:0]) +
	( 16'sd 28089) * $signed(input_fmap_40[15:0]) +
	( 13'sd 2708) * $signed(input_fmap_41[15:0]) +
	( 14'sd 6146) * $signed(input_fmap_42[15:0]) +
	( 16'sd 27653) * $signed(input_fmap_43[15:0]) +
	( 14'sd 4352) * $signed(input_fmap_44[15:0]) +
	( 16'sd 28064) * $signed(input_fmap_45[15:0]) +
	( 15'sd 11817) * $signed(input_fmap_46[15:0]) +
	( 16'sd 31931) * $signed(input_fmap_47[15:0]) +
	( 16'sd 17230) * $signed(input_fmap_48[15:0]) +
	( 16'sd 16953) * $signed(input_fmap_49[15:0]) +
	( 16'sd 18261) * $signed(input_fmap_50[15:0]) +
	( 16'sd 19283) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19436) * $signed(input_fmap_52[15:0]) +
	( 16'sd 18836) * $signed(input_fmap_53[15:0]) +
	( 16'sd 21345) * $signed(input_fmap_54[15:0]) +
	( 12'sd 1583) * $signed(input_fmap_55[15:0]) +
	( 16'sd 19080) * $signed(input_fmap_56[15:0]) +
	( 16'sd 19353) * $signed(input_fmap_57[15:0]) +
	( 16'sd 28110) * $signed(input_fmap_58[15:0]) +
	( 15'sd 9764) * $signed(input_fmap_59[15:0]) +
	( 15'sd 12115) * $signed(input_fmap_60[15:0]) +
	( 5'sd 8) * $signed(input_fmap_61[15:0]) +
	( 14'sd 4317) * $signed(input_fmap_62[15:0]) +
	( 15'sd 9390) * $signed(input_fmap_63[15:0]) +
	( 9'sd 249) * $signed(input_fmap_64[15:0]) +
	( 16'sd 29892) * $signed(input_fmap_65[15:0]) +
	( 16'sd 31916) * $signed(input_fmap_66[15:0]) +
	( 15'sd 14052) * $signed(input_fmap_67[15:0]) +
	( 16'sd 27964) * $signed(input_fmap_68[15:0]) +
	( 16'sd 25427) * $signed(input_fmap_69[15:0]) +
	( 15'sd 10831) * $signed(input_fmap_70[15:0]) +
	( 14'sd 4145) * $signed(input_fmap_71[15:0]) +
	( 16'sd 30558) * $signed(input_fmap_72[15:0]) +
	( 16'sd 22373) * $signed(input_fmap_73[15:0]) +
	( 15'sd 10615) * $signed(input_fmap_74[15:0]) +
	( 15'sd 9618) * $signed(input_fmap_75[15:0]) +
	( 16'sd 30936) * $signed(input_fmap_76[15:0]) +
	( 15'sd 14380) * $signed(input_fmap_77[15:0]) +
	( 14'sd 4716) * $signed(input_fmap_78[15:0]) +
	( 16'sd 20467) * $signed(input_fmap_79[15:0]) +
	( 15'sd 13823) * $signed(input_fmap_80[15:0]) +
	( 15'sd 13858) * $signed(input_fmap_81[15:0]) +
	( 16'sd 20897) * $signed(input_fmap_82[15:0]) +
	( 16'sd 27180) * $signed(input_fmap_83[15:0]) +
	( 16'sd 22511) * $signed(input_fmap_84[15:0]) +
	( 16'sd 17075) * $signed(input_fmap_85[15:0]) +
	( 16'sd 28670) * $signed(input_fmap_86[15:0]) +
	( 15'sd 10292) * $signed(input_fmap_87[15:0]) +
	( 12'sd 1369) * $signed(input_fmap_88[15:0]) +
	( 15'sd 9283) * $signed(input_fmap_89[15:0]) +
	( 16'sd 19221) * $signed(input_fmap_90[15:0]) +
	( 7'sd 51) * $signed(input_fmap_91[15:0]) +
	( 15'sd 12376) * $signed(input_fmap_92[15:0]) +
	( 15'sd 13230) * $signed(input_fmap_93[15:0]) +
	( 15'sd 9011) * $signed(input_fmap_94[15:0]) +
	( 16'sd 22340) * $signed(input_fmap_95[15:0]) +
	( 16'sd 27594) * $signed(input_fmap_96[15:0]) +
	( 16'sd 32239) * $signed(input_fmap_97[15:0]) +
	( 16'sd 30033) * $signed(input_fmap_98[15:0]) +
	( 15'sd 14830) * $signed(input_fmap_99[15:0]) +
	( 15'sd 8518) * $signed(input_fmap_100[15:0]) +
	( 16'sd 24100) * $signed(input_fmap_101[15:0]) +
	( 15'sd 15300) * $signed(input_fmap_102[15:0]) +
	( 16'sd 27645) * $signed(input_fmap_103[15:0]) +
	( 16'sd 27970) * $signed(input_fmap_104[15:0]) +
	( 13'sd 3222) * $signed(input_fmap_105[15:0]) +
	( 15'sd 12896) * $signed(input_fmap_106[15:0]) +
	( 15'sd 15388) * $signed(input_fmap_107[15:0]) +
	( 13'sd 3012) * $signed(input_fmap_108[15:0]) +
	( 16'sd 17155) * $signed(input_fmap_109[15:0]) +
	( 16'sd 29531) * $signed(input_fmap_110[15:0]) +
	( 16'sd 24444) * $signed(input_fmap_111[15:0]) +
	( 14'sd 6993) * $signed(input_fmap_112[15:0]) +
	( 16'sd 26921) * $signed(input_fmap_113[15:0]) +
	( 16'sd 29228) * $signed(input_fmap_114[15:0]) +
	( 15'sd 16018) * $signed(input_fmap_115[15:0]) +
	( 16'sd 30211) * $signed(input_fmap_116[15:0]) +
	( 14'sd 5228) * $signed(input_fmap_117[15:0]) +
	( 16'sd 21405) * $signed(input_fmap_118[15:0]) +
	( 14'sd 6231) * $signed(input_fmap_119[15:0]) +
	( 16'sd 23105) * $signed(input_fmap_120[15:0]) +
	( 14'sd 6743) * $signed(input_fmap_121[15:0]) +
	( 15'sd 15451) * $signed(input_fmap_122[15:0]) +
	( 16'sd 29887) * $signed(input_fmap_123[15:0]) +
	( 15'sd 13990) * $signed(input_fmap_124[15:0]) +
	( 13'sd 3046) * $signed(input_fmap_125[15:0]) +
	( 16'sd 28293) * $signed(input_fmap_126[15:0]) +
	( 15'sd 12573) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 16'sd 26633) * $signed(input_fmap_0[15:0]) +
	( 16'sd 19765) * $signed(input_fmap_1[15:0]) +
	( 16'sd 31697) * $signed(input_fmap_2[15:0]) +
	( 16'sd 22106) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30774) * $signed(input_fmap_4[15:0]) +
	( 16'sd 23630) * $signed(input_fmap_5[15:0]) +
	( 10'sd 370) * $signed(input_fmap_6[15:0]) +
	( 15'sd 8665) * $signed(input_fmap_7[15:0]) +
	( 16'sd 22145) * $signed(input_fmap_8[15:0]) +
	( 16'sd 26497) * $signed(input_fmap_9[15:0]) +
	( 16'sd 28099) * $signed(input_fmap_10[15:0]) +
	( 15'sd 13109) * $signed(input_fmap_11[15:0]) +
	( 16'sd 23243) * $signed(input_fmap_12[15:0]) +
	( 15'sd 10124) * $signed(input_fmap_13[15:0]) +
	( 15'sd 16192) * $signed(input_fmap_14[15:0]) +
	( 14'sd 7301) * $signed(input_fmap_15[15:0]) +
	( 16'sd 24309) * $signed(input_fmap_16[15:0]) +
	( 15'sd 12377) * $signed(input_fmap_17[15:0]) +
	( 14'sd 6391) * $signed(input_fmap_18[15:0]) +
	( 14'sd 8155) * $signed(input_fmap_19[15:0]) +
	( 15'sd 9130) * $signed(input_fmap_20[15:0]) +
	( 10'sd 464) * $signed(input_fmap_21[15:0]) +
	( 12'sd 1627) * $signed(input_fmap_22[15:0]) +
	( 16'sd 18163) * $signed(input_fmap_23[15:0]) +
	( 16'sd 30693) * $signed(input_fmap_24[15:0]) +
	( 16'sd 22595) * $signed(input_fmap_25[15:0]) +
	( 16'sd 18773) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2798) * $signed(input_fmap_27[15:0]) +
	( 16'sd 19488) * $signed(input_fmap_28[15:0]) +
	( 16'sd 23662) * $signed(input_fmap_29[15:0]) +
	( 16'sd 31777) * $signed(input_fmap_30[15:0]) +
	( 10'sd 449) * $signed(input_fmap_31[15:0]) +
	( 16'sd 25966) * $signed(input_fmap_32[15:0]) +
	( 14'sd 4468) * $signed(input_fmap_33[15:0]) +
	( 12'sd 1747) * $signed(input_fmap_34[15:0]) +
	( 15'sd 8821) * $signed(input_fmap_35[15:0]) +
	( 16'sd 28918) * $signed(input_fmap_36[15:0]) +
	( 15'sd 9811) * $signed(input_fmap_37[15:0]) +
	( 16'sd 31810) * $signed(input_fmap_38[15:0]) +
	( 16'sd 30436) * $signed(input_fmap_39[15:0]) +
	( 16'sd 21601) * $signed(input_fmap_40[15:0]) +
	( 16'sd 28353) * $signed(input_fmap_41[15:0]) +
	( 16'sd 16519) * $signed(input_fmap_42[15:0]) +
	( 12'sd 1598) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31996) * $signed(input_fmap_44[15:0]) +
	( 13'sd 3526) * $signed(input_fmap_45[15:0]) +
	( 16'sd 22746) * $signed(input_fmap_46[15:0]) +
	( 16'sd 22304) * $signed(input_fmap_47[15:0]) +
	( 16'sd 17133) * $signed(input_fmap_48[15:0]) +
	( 16'sd 26963) * $signed(input_fmap_49[15:0]) +
	( 16'sd 28261) * $signed(input_fmap_50[15:0]) +
	( 14'sd 8040) * $signed(input_fmap_51[15:0]) +
	( 16'sd 25041) * $signed(input_fmap_52[15:0]) +
	( 16'sd 19538) * $signed(input_fmap_53[15:0]) +
	( 15'sd 9320) * $signed(input_fmap_54[15:0]) +
	( 14'sd 7027) * $signed(input_fmap_55[15:0]) +
	( 15'sd 9501) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17987) * $signed(input_fmap_57[15:0]) +
	( 16'sd 24840) * $signed(input_fmap_58[15:0]) +
	( 15'sd 8813) * $signed(input_fmap_59[15:0]) +
	( 15'sd 9599) * $signed(input_fmap_60[15:0]) +
	( 13'sd 2059) * $signed(input_fmap_61[15:0]) +
	( 16'sd 20512) * $signed(input_fmap_62[15:0]) +
	( 16'sd 19093) * $signed(input_fmap_63[15:0]) +
	( 14'sd 6314) * $signed(input_fmap_64[15:0]) +
	( 16'sd 16502) * $signed(input_fmap_65[15:0]) +
	( 15'sd 8411) * $signed(input_fmap_66[15:0]) +
	( 15'sd 10322) * $signed(input_fmap_67[15:0]) +
	( 16'sd 28209) * $signed(input_fmap_68[15:0]) +
	( 12'sd 1762) * $signed(input_fmap_69[15:0]) +
	( 13'sd 3869) * $signed(input_fmap_70[15:0]) +
	( 16'sd 30903) * $signed(input_fmap_71[15:0]) +
	( 15'sd 9694) * $signed(input_fmap_72[15:0]) +
	( 15'sd 16200) * $signed(input_fmap_73[15:0]) +
	( 16'sd 18628) * $signed(input_fmap_74[15:0]) +
	( 15'sd 12599) * $signed(input_fmap_75[15:0]) +
	( 12'sd 1139) * $signed(input_fmap_76[15:0]) +
	( 16'sd 18198) * $signed(input_fmap_77[15:0]) +
	( 14'sd 7019) * $signed(input_fmap_78[15:0]) +
	( 16'sd 22184) * $signed(input_fmap_79[15:0]) +
	( 16'sd 19206) * $signed(input_fmap_80[15:0]) +
	( 16'sd 20867) * $signed(input_fmap_81[15:0]) +
	( 16'sd 23071) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25429) * $signed(input_fmap_83[15:0]) +
	( 15'sd 15357) * $signed(input_fmap_84[15:0]) +
	( 16'sd 21444) * $signed(input_fmap_85[15:0]) +
	( 16'sd 16868) * $signed(input_fmap_86[15:0]) +
	( 7'sd 53) * $signed(input_fmap_87[15:0]) +
	( 14'sd 5638) * $signed(input_fmap_88[15:0]) +
	( 15'sd 13262) * $signed(input_fmap_89[15:0]) +
	( 16'sd 27827) * $signed(input_fmap_90[15:0]) +
	( 12'sd 1261) * $signed(input_fmap_91[15:0]) +
	( 13'sd 2727) * $signed(input_fmap_92[15:0]) +
	( 14'sd 5787) * $signed(input_fmap_93[15:0]) +
	( 16'sd 29861) * $signed(input_fmap_94[15:0]) +
	( 16'sd 29919) * $signed(input_fmap_95[15:0]) +
	( 16'sd 31918) * $signed(input_fmap_96[15:0]) +
	( 14'sd 7396) * $signed(input_fmap_97[15:0]) +
	( 15'sd 9962) * $signed(input_fmap_98[15:0]) +
	( 15'sd 14962) * $signed(input_fmap_99[15:0]) +
	( 16'sd 27393) * $signed(input_fmap_100[15:0]) +
	( 14'sd 4715) * $signed(input_fmap_101[15:0]) +
	( 15'sd 15145) * $signed(input_fmap_102[15:0]) +
	( 16'sd 29146) * $signed(input_fmap_103[15:0]) +
	( 14'sd 7116) * $signed(input_fmap_104[15:0]) +
	( 12'sd 1198) * $signed(input_fmap_105[15:0]) +
	( 16'sd 19301) * $signed(input_fmap_106[15:0]) +
	( 16'sd 24942) * $signed(input_fmap_107[15:0]) +
	( 15'sd 10314) * $signed(input_fmap_108[15:0]) +
	( 11'sd 607) * $signed(input_fmap_109[15:0]) +
	( 11'sd 643) * $signed(input_fmap_110[15:0]) +
	( 16'sd 24571) * $signed(input_fmap_111[15:0]) +
	( 16'sd 19583) * $signed(input_fmap_112[15:0]) +
	( 14'sd 5122) * $signed(input_fmap_113[15:0]) +
	( 15'sd 12732) * $signed(input_fmap_114[15:0]) +
	( 15'sd 10278) * $signed(input_fmap_115[15:0]) +
	( 14'sd 5976) * $signed(input_fmap_116[15:0]) +
	( 16'sd 22746) * $signed(input_fmap_117[15:0]) +
	( 14'sd 5961) * $signed(input_fmap_118[15:0]) +
	( 16'sd 27390) * $signed(input_fmap_119[15:0]) +
	( 14'sd 6758) * $signed(input_fmap_120[15:0]) +
	( 16'sd 28713) * $signed(input_fmap_121[15:0]) +
	( 12'sd 1331) * $signed(input_fmap_122[15:0]) +
	( 16'sd 31904) * $signed(input_fmap_123[15:0]) +
	( 16'sd 28713) * $signed(input_fmap_124[15:0]) +
	( 16'sd 19350) * $signed(input_fmap_125[15:0]) +
	( 16'sd 29630) * $signed(input_fmap_126[15:0]) +
	( 15'sd 14355) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 16'sd 28129) * $signed(input_fmap_0[15:0]) +
	( 16'sd 28382) * $signed(input_fmap_1[15:0]) +
	( 16'sd 27926) * $signed(input_fmap_2[15:0]) +
	( 16'sd 28414) * $signed(input_fmap_3[15:0]) +
	( 16'sd 31551) * $signed(input_fmap_4[15:0]) +
	( 16'sd 19690) * $signed(input_fmap_5[15:0]) +
	( 16'sd 32581) * $signed(input_fmap_6[15:0]) +
	( 15'sd 9163) * $signed(input_fmap_7[15:0]) +
	( 15'sd 15977) * $signed(input_fmap_8[15:0]) +
	( 15'sd 9003) * $signed(input_fmap_9[15:0]) +
	( 16'sd 23418) * $signed(input_fmap_10[15:0]) +
	( 16'sd 25989) * $signed(input_fmap_11[15:0]) +
	( 16'sd 23500) * $signed(input_fmap_12[15:0]) +
	( 13'sd 2970) * $signed(input_fmap_13[15:0]) +
	( 11'sd 743) * $signed(input_fmap_14[15:0]) +
	( 15'sd 8493) * $signed(input_fmap_15[15:0]) +
	( 15'sd 8196) * $signed(input_fmap_16[15:0]) +
	( 14'sd 4904) * $signed(input_fmap_17[15:0]) +
	( 14'sd 5086) * $signed(input_fmap_18[15:0]) +
	( 16'sd 17044) * $signed(input_fmap_19[15:0]) +
	( 15'sd 11710) * $signed(input_fmap_20[15:0]) +
	( 16'sd 21710) * $signed(input_fmap_21[15:0]) +
	( 14'sd 6480) * $signed(input_fmap_22[15:0]) +
	( 13'sd 3356) * $signed(input_fmap_23[15:0]) +
	( 15'sd 12742) * $signed(input_fmap_24[15:0]) +
	( 16'sd 18747) * $signed(input_fmap_25[15:0]) +
	( 14'sd 6814) * $signed(input_fmap_26[15:0]) +
	( 14'sd 6737) * $signed(input_fmap_27[15:0]) +
	( 16'sd 28814) * $signed(input_fmap_28[15:0]) +
	( 15'sd 12954) * $signed(input_fmap_29[15:0]) +
	( 15'sd 10383) * $signed(input_fmap_30[15:0]) +
	( 16'sd 19063) * $signed(input_fmap_31[15:0]) +
	( 14'sd 6087) * $signed(input_fmap_32[15:0]) +
	( 15'sd 12692) * $signed(input_fmap_33[15:0]) +
	( 13'sd 3600) * $signed(input_fmap_34[15:0]) +
	( 16'sd 22171) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11397) * $signed(input_fmap_36[15:0]) +
	( 16'sd 21937) * $signed(input_fmap_37[15:0]) +
	( 16'sd 21768) * $signed(input_fmap_38[15:0]) +
	( 16'sd 21771) * $signed(input_fmap_39[15:0]) +
	( 15'sd 10595) * $signed(input_fmap_40[15:0]) +
	( 15'sd 12507) * $signed(input_fmap_41[15:0]) +
	( 14'sd 7503) * $signed(input_fmap_42[15:0]) +
	( 15'sd 13760) * $signed(input_fmap_43[15:0]) +
	( 16'sd 24170) * $signed(input_fmap_44[15:0]) +
	( 16'sd 18212) * $signed(input_fmap_45[15:0]) +
	( 16'sd 16623) * $signed(input_fmap_46[15:0]) +
	( 15'sd 8434) * $signed(input_fmap_47[15:0]) +
	( 13'sd 3559) * $signed(input_fmap_48[15:0]) +
	( 12'sd 1967) * $signed(input_fmap_49[15:0]) +
	( 16'sd 32282) * $signed(input_fmap_50[15:0]) +
	( 13'sd 3522) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19261) * $signed(input_fmap_52[15:0]) +
	( 15'sd 9009) * $signed(input_fmap_53[15:0]) +
	( 10'sd 437) * $signed(input_fmap_54[15:0]) +
	( 15'sd 12081) * $signed(input_fmap_55[15:0]) +
	( 16'sd 31713) * $signed(input_fmap_56[15:0]) +
	( 13'sd 2200) * $signed(input_fmap_57[15:0]) +
	( 16'sd 29778) * $signed(input_fmap_58[15:0]) +
	( 16'sd 29810) * $signed(input_fmap_59[15:0]) +
	( 16'sd 31168) * $signed(input_fmap_60[15:0]) +
	( 16'sd 23806) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3100) * $signed(input_fmap_62[15:0]) +
	( 15'sd 9962) * $signed(input_fmap_63[15:0]) +
	( 16'sd 22068) * $signed(input_fmap_64[15:0]) +
	( 14'sd 7203) * $signed(input_fmap_65[15:0]) +
	( 13'sd 3946) * $signed(input_fmap_66[15:0]) +
	( 16'sd 19691) * $signed(input_fmap_67[15:0]) +
	( 11'sd 614) * $signed(input_fmap_68[15:0]) +
	( 16'sd 26895) * $signed(input_fmap_69[15:0]) +
	( 11'sd 991) * $signed(input_fmap_70[15:0]) +
	( 14'sd 6148) * $signed(input_fmap_71[15:0]) +
	( 12'sd 1359) * $signed(input_fmap_72[15:0]) +
	( 13'sd 3187) * $signed(input_fmap_73[15:0]) +
	( 16'sd 23832) * $signed(input_fmap_74[15:0]) +
	( 14'sd 6557) * $signed(input_fmap_75[15:0]) +
	( 16'sd 20131) * $signed(input_fmap_76[15:0]) +
	( 15'sd 13817) * $signed(input_fmap_77[15:0]) +
	( 14'sd 5782) * $signed(input_fmap_78[15:0]) +
	( 16'sd 27174) * $signed(input_fmap_79[15:0]) +
	( 8'sd 111) * $signed(input_fmap_80[15:0]) +
	( 15'sd 8247) * $signed(input_fmap_81[15:0]) +
	( 16'sd 17489) * $signed(input_fmap_82[15:0]) +
	( 16'sd 24851) * $signed(input_fmap_83[15:0]) +
	( 16'sd 27073) * $signed(input_fmap_84[15:0]) +
	( 16'sd 26657) * $signed(input_fmap_85[15:0]) +
	( 14'sd 6777) * $signed(input_fmap_86[15:0]) +
	( 6'sd 22) * $signed(input_fmap_87[15:0]) +
	( 16'sd 23074) * $signed(input_fmap_88[15:0]) +
	( 14'sd 6688) * $signed(input_fmap_89[15:0]) +
	( 16'sd 16708) * $signed(input_fmap_90[15:0]) +
	( 16'sd 32539) * $signed(input_fmap_91[15:0]) +
	( 16'sd 31277) * $signed(input_fmap_92[15:0]) +
	( 16'sd 30675) * $signed(input_fmap_93[15:0]) +
	( 16'sd 27342) * $signed(input_fmap_94[15:0]) +
	( 14'sd 7556) * $signed(input_fmap_95[15:0]) +
	( 13'sd 2664) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27401) * $signed(input_fmap_97[15:0]) +
	( 14'sd 8145) * $signed(input_fmap_98[15:0]) +
	( 16'sd 25374) * $signed(input_fmap_99[15:0]) +
	( 9'sd 155) * $signed(input_fmap_100[15:0]) +
	( 12'sd 1210) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5383) * $signed(input_fmap_102[15:0]) +
	( 16'sd 25997) * $signed(input_fmap_103[15:0]) +
	( 14'sd 5362) * $signed(input_fmap_104[15:0]) +
	( 14'sd 4818) * $signed(input_fmap_105[15:0]) +
	( 16'sd 30670) * $signed(input_fmap_106[15:0]) +
	( 16'sd 31768) * $signed(input_fmap_107[15:0]) +
	( 16'sd 31701) * $signed(input_fmap_108[15:0]) +
	( 12'sd 1166) * $signed(input_fmap_109[15:0]) +
	( 12'sd 1458) * $signed(input_fmap_110[15:0]) +
	( 14'sd 7861) * $signed(input_fmap_111[15:0]) +
	( 15'sd 8354) * $signed(input_fmap_112[15:0]) +
	( 14'sd 4807) * $signed(input_fmap_113[15:0]) +
	( 16'sd 25511) * $signed(input_fmap_114[15:0]) +
	( 16'sd 25290) * $signed(input_fmap_115[15:0]) +
	( 16'sd 21950) * $signed(input_fmap_116[15:0]) +
	( 16'sd 26247) * $signed(input_fmap_117[15:0]) +
	( 16'sd 29510) * $signed(input_fmap_118[15:0]) +
	( 16'sd 23159) * $signed(input_fmap_119[15:0]) +
	( 14'sd 5221) * $signed(input_fmap_120[15:0]) +
	( 16'sd 23799) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9422) * $signed(input_fmap_122[15:0]) +
	( 12'sd 1590) * $signed(input_fmap_123[15:0]) +
	( 13'sd 3148) * $signed(input_fmap_124[15:0]) +
	( 15'sd 11292) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6694) * $signed(input_fmap_126[15:0]) +
	( 16'sd 19392) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 16'sd 25620) * $signed(input_fmap_0[15:0]) +
	( 15'sd 14252) * $signed(input_fmap_1[15:0]) +
	( 15'sd 9281) * $signed(input_fmap_2[15:0]) +
	( 14'sd 5702) * $signed(input_fmap_3[15:0]) +
	( 16'sd 19205) * $signed(input_fmap_4[15:0]) +
	( 16'sd 23044) * $signed(input_fmap_5[15:0]) +
	( 16'sd 17518) * $signed(input_fmap_6[15:0]) +
	( 13'sd 2350) * $signed(input_fmap_7[15:0]) +
	( 16'sd 31521) * $signed(input_fmap_8[15:0]) +
	( 14'sd 6697) * $signed(input_fmap_9[15:0]) +
	( 16'sd 32187) * $signed(input_fmap_10[15:0]) +
	( 16'sd 21840) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20756) * $signed(input_fmap_12[15:0]) +
	( 15'sd 11433) * $signed(input_fmap_13[15:0]) +
	( 15'sd 15686) * $signed(input_fmap_14[15:0]) +
	( 15'sd 13886) * $signed(input_fmap_15[15:0]) +
	( 16'sd 25335) * $signed(input_fmap_16[15:0]) +
	( 16'sd 22571) * $signed(input_fmap_17[15:0]) +
	( 12'sd 1029) * $signed(input_fmap_18[15:0]) +
	( 10'sd 354) * $signed(input_fmap_19[15:0]) +
	( 16'sd 18077) * $signed(input_fmap_20[15:0]) +
	( 16'sd 22634) * $signed(input_fmap_21[15:0]) +
	( 16'sd 22822) * $signed(input_fmap_22[15:0]) +
	( 15'sd 12837) * $signed(input_fmap_23[15:0]) +
	( 15'sd 11911) * $signed(input_fmap_24[15:0]) +
	( 16'sd 23993) * $signed(input_fmap_25[15:0]) +
	( 16'sd 20509) * $signed(input_fmap_26[15:0]) +
	( 15'sd 15362) * $signed(input_fmap_27[15:0]) +
	( 15'sd 11856) * $signed(input_fmap_28[15:0]) +
	( 16'sd 19521) * $signed(input_fmap_29[15:0]) +
	( 16'sd 31740) * $signed(input_fmap_30[15:0]) +
	( 16'sd 18884) * $signed(input_fmap_31[15:0]) +
	( 15'sd 12255) * $signed(input_fmap_32[15:0]) +
	( 13'sd 3167) * $signed(input_fmap_33[15:0]) +
	( 16'sd 22657) * $signed(input_fmap_34[15:0]) +
	( 16'sd 21138) * $signed(input_fmap_35[15:0]) +
	( 15'sd 12616) * $signed(input_fmap_36[15:0]) +
	( 15'sd 13033) * $signed(input_fmap_37[15:0]) +
	( 12'sd 2006) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24922) * $signed(input_fmap_39[15:0]) +
	( 16'sd 19319) * $signed(input_fmap_40[15:0]) +
	( 16'sd 16611) * $signed(input_fmap_41[15:0]) +
	( 16'sd 31436) * $signed(input_fmap_42[15:0]) +
	( 16'sd 28906) * $signed(input_fmap_43[15:0]) +
	( 15'sd 10896) * $signed(input_fmap_44[15:0]) +
	( 16'sd 25265) * $signed(input_fmap_45[15:0]) +
	( 16'sd 25121) * $signed(input_fmap_46[15:0]) +
	( 16'sd 31641) * $signed(input_fmap_47[15:0]) +
	( 15'sd 9264) * $signed(input_fmap_48[15:0]) +
	( 16'sd 19447) * $signed(input_fmap_49[15:0]) +
	( 14'sd 7458) * $signed(input_fmap_50[15:0]) +
	( 16'sd 18190) * $signed(input_fmap_51[15:0]) +
	( 13'sd 2362) * $signed(input_fmap_52[15:0]) +
	( 16'sd 17688) * $signed(input_fmap_53[15:0]) +
	( 16'sd 18133) * $signed(input_fmap_54[15:0]) +
	( 15'sd 13809) * $signed(input_fmap_55[15:0]) +
	( 12'sd 1386) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17331) * $signed(input_fmap_57[15:0]) +
	( 16'sd 31468) * $signed(input_fmap_58[15:0]) +
	( 16'sd 28404) * $signed(input_fmap_59[15:0]) +
	( 14'sd 6875) * $signed(input_fmap_60[15:0]) +
	( 15'sd 13654) * $signed(input_fmap_61[15:0]) +
	( 15'sd 13694) * $signed(input_fmap_62[15:0]) +
	( 16'sd 25592) * $signed(input_fmap_63[15:0]) +
	( 16'sd 19052) * $signed(input_fmap_64[15:0]) +
	( 16'sd 24121) * $signed(input_fmap_65[15:0]) +
	( 13'sd 2958) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28830) * $signed(input_fmap_67[15:0]) +
	( 15'sd 8237) * $signed(input_fmap_68[15:0]) +
	( 14'sd 6946) * $signed(input_fmap_69[15:0]) +
	( 14'sd 5199) * $signed(input_fmap_70[15:0]) +
	( 13'sd 3158) * $signed(input_fmap_71[15:0]) +
	( 14'sd 6562) * $signed(input_fmap_72[15:0]) +
	( 15'sd 13533) * $signed(input_fmap_73[15:0]) +
	( 14'sd 5749) * $signed(input_fmap_74[15:0]) +
	( 15'sd 13598) * $signed(input_fmap_75[15:0]) +
	( 14'sd 4314) * $signed(input_fmap_76[15:0]) +
	( 14'sd 6580) * $signed(input_fmap_77[15:0]) +
	( 16'sd 20395) * $signed(input_fmap_78[15:0]) +
	( 14'sd 5134) * $signed(input_fmap_79[15:0]) +
	( 10'sd 289) * $signed(input_fmap_80[15:0]) +
	( 16'sd 26431) * $signed(input_fmap_81[15:0]) +
	( 16'sd 23196) * $signed(input_fmap_82[15:0]) +
	( 16'sd 28860) * $signed(input_fmap_83[15:0]) +
	( 11'sd 709) * $signed(input_fmap_84[15:0]) +
	( 15'sd 14311) * $signed(input_fmap_85[15:0]) +
	( 16'sd 26070) * $signed(input_fmap_86[15:0]) +
	( 15'sd 12982) * $signed(input_fmap_87[15:0]) +
	( 16'sd 25496) * $signed(input_fmap_88[15:0]) +
	( 15'sd 12346) * $signed(input_fmap_89[15:0]) +
	( 15'sd 15336) * $signed(input_fmap_90[15:0]) +
	( 15'sd 11133) * $signed(input_fmap_91[15:0]) +
	( 12'sd 1128) * $signed(input_fmap_92[15:0]) +
	( 14'sd 6087) * $signed(input_fmap_93[15:0]) +
	( 13'sd 2780) * $signed(input_fmap_94[15:0]) +
	( 13'sd 2808) * $signed(input_fmap_95[15:0]) +
	( 15'sd 13646) * $signed(input_fmap_96[15:0]) +
	( 16'sd 28456) * $signed(input_fmap_97[15:0]) +
	( 16'sd 16862) * $signed(input_fmap_98[15:0]) +
	( 14'sd 4991) * $signed(input_fmap_99[15:0]) +
	( 14'sd 4783) * $signed(input_fmap_100[15:0]) +
	( 16'sd 31737) * $signed(input_fmap_101[15:0]) +
	( 12'sd 1275) * $signed(input_fmap_102[15:0]) +
	( 14'sd 6394) * $signed(input_fmap_103[15:0]) +
	( 13'sd 4028) * $signed(input_fmap_104[15:0]) +
	( 15'sd 15767) * $signed(input_fmap_105[15:0]) +
	( 15'sd 10575) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27022) * $signed(input_fmap_107[15:0]) +
	( 16'sd 30403) * $signed(input_fmap_108[15:0]) +
	( 16'sd 27410) * $signed(input_fmap_109[15:0]) +
	( 15'sd 15913) * $signed(input_fmap_110[15:0]) +
	( 16'sd 24593) * $signed(input_fmap_111[15:0]) +
	( 14'sd 7582) * $signed(input_fmap_112[15:0]) +
	( 16'sd 25591) * $signed(input_fmap_113[15:0]) +
	( 14'sd 6344) * $signed(input_fmap_114[15:0]) +
	( 16'sd 27308) * $signed(input_fmap_115[15:0]) +
	( 13'sd 2557) * $signed(input_fmap_116[15:0]) +
	( 13'sd 3278) * $signed(input_fmap_117[15:0]) +
	( 13'sd 3918) * $signed(input_fmap_118[15:0]) +
	( 14'sd 7418) * $signed(input_fmap_119[15:0]) +
	( 6'sd 25) * $signed(input_fmap_120[15:0]) +
	( 12'sd 1522) * $signed(input_fmap_121[15:0]) +
	( 15'sd 14825) * $signed(input_fmap_122[15:0]) +
	( 16'sd 24819) * $signed(input_fmap_123[15:0]) +
	( 15'sd 15692) * $signed(input_fmap_124[15:0]) +
	( 15'sd 13971) * $signed(input_fmap_125[15:0]) +
	( 16'sd 19438) * $signed(input_fmap_126[15:0]) +
	( 13'sd 2892) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 15'sd 8430) * $signed(input_fmap_0[15:0]) +
	( 16'sd 32284) * $signed(input_fmap_1[15:0]) +
	( 15'sd 13660) * $signed(input_fmap_2[15:0]) +
	( 15'sd 15176) * $signed(input_fmap_3[15:0]) +
	( 16'sd 21116) * $signed(input_fmap_4[15:0]) +
	( 15'sd 12484) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2445) * $signed(input_fmap_6[15:0]) +
	( 16'sd 30931) * $signed(input_fmap_7[15:0]) +
	( 16'sd 24967) * $signed(input_fmap_8[15:0]) +
	( 14'sd 4524) * $signed(input_fmap_9[15:0]) +
	( 15'sd 15819) * $signed(input_fmap_10[15:0]) +
	( 14'sd 7830) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20209) * $signed(input_fmap_12[15:0]) +
	( 16'sd 23751) * $signed(input_fmap_13[15:0]) +
	( 16'sd 26866) * $signed(input_fmap_14[15:0]) +
	( 15'sd 11282) * $signed(input_fmap_15[15:0]) +
	( 16'sd 25753) * $signed(input_fmap_16[15:0]) +
	( 15'sd 15652) * $signed(input_fmap_17[15:0]) +
	( 14'sd 7218) * $signed(input_fmap_18[15:0]) +
	( 13'sd 3116) * $signed(input_fmap_19[15:0]) +
	( 16'sd 18415) * $signed(input_fmap_20[15:0]) +
	( 16'sd 23339) * $signed(input_fmap_21[15:0]) +
	( 15'sd 14862) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28424) * $signed(input_fmap_23[15:0]) +
	( 15'sd 11784) * $signed(input_fmap_24[15:0]) +
	( 16'sd 27949) * $signed(input_fmap_25[15:0]) +
	( 16'sd 28754) * $signed(input_fmap_26[15:0]) +
	( 16'sd 19951) * $signed(input_fmap_27[15:0]) +
	( 16'sd 18922) * $signed(input_fmap_28[15:0]) +
	( 15'sd 10321) * $signed(input_fmap_29[15:0]) +
	( 14'sd 5486) * $signed(input_fmap_30[15:0]) +
	( 15'sd 15136) * $signed(input_fmap_31[15:0]) +
	( 14'sd 4515) * $signed(input_fmap_32[15:0]) +
	( 16'sd 28878) * $signed(input_fmap_33[15:0]) +
	( 16'sd 17672) * $signed(input_fmap_34[15:0]) +
	( 16'sd 20184) * $signed(input_fmap_35[15:0]) +
	( 16'sd 18026) * $signed(input_fmap_36[15:0]) +
	( 16'sd 21987) * $signed(input_fmap_37[15:0]) +
	( 14'sd 7196) * $signed(input_fmap_38[15:0]) +
	( 14'sd 6974) * $signed(input_fmap_39[15:0]) +
	( 15'sd 12452) * $signed(input_fmap_40[15:0]) +
	( 16'sd 30287) * $signed(input_fmap_41[15:0]) +
	( 16'sd 29420) * $signed(input_fmap_42[15:0]) +
	( 16'sd 27386) * $signed(input_fmap_43[15:0]) +
	( 14'sd 5326) * $signed(input_fmap_44[15:0]) +
	( 15'sd 14339) * $signed(input_fmap_45[15:0]) +
	( 13'sd 3973) * $signed(input_fmap_46[15:0]) +
	( 16'sd 18044) * $signed(input_fmap_47[15:0]) +
	( 8'sd 72) * $signed(input_fmap_48[15:0]) +
	( 14'sd 7776) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22222) * $signed(input_fmap_50[15:0]) +
	( 12'sd 1602) * $signed(input_fmap_51[15:0]) +
	( 15'sd 13509) * $signed(input_fmap_52[15:0]) +
	( 16'sd 21131) * $signed(input_fmap_53[15:0]) +
	( 16'sd 16819) * $signed(input_fmap_54[15:0]) +
	( 14'sd 6014) * $signed(input_fmap_55[15:0]) +
	( 16'sd 20280) * $signed(input_fmap_56[15:0]) +
	( 16'sd 21604) * $signed(input_fmap_57[15:0]) +
	( 16'sd 21283) * $signed(input_fmap_58[15:0]) +
	( 16'sd 18658) * $signed(input_fmap_59[15:0]) +
	( 15'sd 12970) * $signed(input_fmap_60[15:0]) +
	( 15'sd 12197) * $signed(input_fmap_61[15:0]) +
	( 14'sd 6519) * $signed(input_fmap_62[15:0]) +
	( 16'sd 28932) * $signed(input_fmap_63[15:0]) +
	( 15'sd 15568) * $signed(input_fmap_64[15:0]) +
	( 14'sd 6384) * $signed(input_fmap_65[15:0]) +
	( 16'sd 17080) * $signed(input_fmap_66[15:0]) +
	( 13'sd 2879) * $signed(input_fmap_67[15:0]) +
	( 7'sd 39) * $signed(input_fmap_68[15:0]) +
	( 16'sd 25428) * $signed(input_fmap_69[15:0]) +
	( 14'sd 7127) * $signed(input_fmap_70[15:0]) +
	( 15'sd 9119) * $signed(input_fmap_71[15:0]) +
	( 11'sd 903) * $signed(input_fmap_72[15:0]) +
	( 16'sd 26521) * $signed(input_fmap_73[15:0]) +
	( 16'sd 31530) * $signed(input_fmap_74[15:0]) +
	( 15'sd 8440) * $signed(input_fmap_75[15:0]) +
	( 16'sd 20350) * $signed(input_fmap_76[15:0]) +
	( 16'sd 18767) * $signed(input_fmap_77[15:0]) +
	( 13'sd 4066) * $signed(input_fmap_78[15:0]) +
	( 15'sd 8979) * $signed(input_fmap_79[15:0]) +
	( 13'sd 3836) * $signed(input_fmap_80[15:0]) +
	( 16'sd 29419) * $signed(input_fmap_81[15:0]) +
	( 9'sd 153) * $signed(input_fmap_82[15:0]) +
	( 16'sd 23713) * $signed(input_fmap_83[15:0]) +
	( 15'sd 10143) * $signed(input_fmap_84[15:0]) +
	( 16'sd 30011) * $signed(input_fmap_85[15:0]) +
	( 16'sd 24613) * $signed(input_fmap_86[15:0]) +
	( 16'sd 25354) * $signed(input_fmap_87[15:0]) +
	( 15'sd 11476) * $signed(input_fmap_88[15:0]) +
	( 16'sd 19194) * $signed(input_fmap_89[15:0]) +
	( 16'sd 19331) * $signed(input_fmap_90[15:0]) +
	( 11'sd 558) * $signed(input_fmap_91[15:0]) +
	( 12'sd 1127) * $signed(input_fmap_92[15:0]) +
	( 13'sd 3106) * $signed(input_fmap_93[15:0]) +
	( 14'sd 6510) * $signed(input_fmap_94[15:0]) +
	( 16'sd 20487) * $signed(input_fmap_95[15:0]) +
	( 13'sd 2129) * $signed(input_fmap_96[15:0]) +
	( 15'sd 11159) * $signed(input_fmap_97[15:0]) +
	( 15'sd 11935) * $signed(input_fmap_98[15:0]) +
	( 16'sd 27611) * $signed(input_fmap_99[15:0]) +
	( 16'sd 23963) * $signed(input_fmap_100[15:0]) +
	( 15'sd 13050) * $signed(input_fmap_101[15:0]) +
	( 16'sd 24191) * $signed(input_fmap_102[15:0]) +
	( 14'sd 7910) * $signed(input_fmap_103[15:0]) +
	( 16'sd 30624) * $signed(input_fmap_104[15:0]) +
	( 15'sd 10039) * $signed(input_fmap_105[15:0]) +
	( 16'sd 20547) * $signed(input_fmap_106[15:0]) +
	( 15'sd 11189) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15708) * $signed(input_fmap_108[15:0]) +
	( 14'sd 6163) * $signed(input_fmap_109[15:0]) +
	( 15'sd 12853) * $signed(input_fmap_110[15:0]) +
	( 16'sd 23239) * $signed(input_fmap_111[15:0]) +
	( 16'sd 29649) * $signed(input_fmap_112[15:0]) +
	( 14'sd 5629) * $signed(input_fmap_113[15:0]) +
	( 15'sd 8864) * $signed(input_fmap_114[15:0]) +
	( 16'sd 25141) * $signed(input_fmap_115[15:0]) +
	( 13'sd 2121) * $signed(input_fmap_116[15:0]) +
	( 16'sd 19041) * $signed(input_fmap_117[15:0]) +
	( 16'sd 28091) * $signed(input_fmap_118[15:0]) +
	( 16'sd 31854) * $signed(input_fmap_119[15:0]) +
	( 16'sd 32305) * $signed(input_fmap_120[15:0]) +
	( 16'sd 18622) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9565) * $signed(input_fmap_122[15:0]) +
	( 15'sd 11787) * $signed(input_fmap_123[15:0]) +
	( 16'sd 25036) * $signed(input_fmap_124[15:0]) +
	( 16'sd 25916) * $signed(input_fmap_125[15:0]) +
	( 15'sd 11898) * $signed(input_fmap_126[15:0]) +
	( 16'sd 28428) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 15'sd 14067) * $signed(input_fmap_0[15:0]) +
	( 16'sd 19138) * $signed(input_fmap_1[15:0]) +
	( 16'sd 26926) * $signed(input_fmap_2[15:0]) +
	( 12'sd 1844) * $signed(input_fmap_3[15:0]) +
	( 15'sd 15250) * $signed(input_fmap_4[15:0]) +
	( 16'sd 19273) * $signed(input_fmap_5[15:0]) +
	( 15'sd 15779) * $signed(input_fmap_6[15:0]) +
	( 16'sd 17401) * $signed(input_fmap_7[15:0]) +
	( 15'sd 12130) * $signed(input_fmap_8[15:0]) +
	( 16'sd 27739) * $signed(input_fmap_9[15:0]) +
	( 16'sd 20365) * $signed(input_fmap_10[15:0]) +
	( 16'sd 26434) * $signed(input_fmap_11[15:0]) +
	( 15'sd 13847) * $signed(input_fmap_12[15:0]) +
	( 16'sd 26987) * $signed(input_fmap_13[15:0]) +
	( 16'sd 31927) * $signed(input_fmap_14[15:0]) +
	( 13'sd 2417) * $signed(input_fmap_15[15:0]) +
	( 16'sd 23026) * $signed(input_fmap_16[15:0]) +
	( 16'sd 31718) * $signed(input_fmap_17[15:0]) +
	( 16'sd 31625) * $signed(input_fmap_18[15:0]) +
	( 16'sd 28073) * $signed(input_fmap_19[15:0]) +
	( 13'sd 2506) * $signed(input_fmap_20[15:0]) +
	( 16'sd 20887) * $signed(input_fmap_21[15:0]) +
	( 14'sd 5170) * $signed(input_fmap_22[15:0]) +
	( 15'sd 15822) * $signed(input_fmap_23[15:0]) +
	( 15'sd 9967) * $signed(input_fmap_24[15:0]) +
	( 16'sd 23919) * $signed(input_fmap_25[15:0]) +
	( 13'sd 2081) * $signed(input_fmap_26[15:0]) +
	( 16'sd 22667) * $signed(input_fmap_27[15:0]) +
	( 16'sd 30683) * $signed(input_fmap_28[15:0]) +
	( 15'sd 9906) * $signed(input_fmap_29[15:0]) +
	( 16'sd 25208) * $signed(input_fmap_30[15:0]) +
	( 16'sd 24128) * $signed(input_fmap_31[15:0]) +
	( 15'sd 12082) * $signed(input_fmap_32[15:0]) +
	( 13'sd 2132) * $signed(input_fmap_33[15:0]) +
	( 15'sd 16094) * $signed(input_fmap_34[15:0]) +
	( 14'sd 7401) * $signed(input_fmap_35[15:0]) +
	( 12'sd 1441) * $signed(input_fmap_36[15:0]) +
	( 14'sd 5506) * $signed(input_fmap_37[15:0]) +
	( 14'sd 5514) * $signed(input_fmap_38[15:0]) +
	( 16'sd 17407) * $signed(input_fmap_39[15:0]) +
	( 16'sd 17203) * $signed(input_fmap_40[15:0]) +
	( 14'sd 7105) * $signed(input_fmap_41[15:0]) +
	( 15'sd 13234) * $signed(input_fmap_42[15:0]) +
	( 16'sd 31794) * $signed(input_fmap_43[15:0]) +
	( 13'sd 2670) * $signed(input_fmap_44[15:0]) +
	( 15'sd 10912) * $signed(input_fmap_45[15:0]) +
	( 16'sd 22312) * $signed(input_fmap_46[15:0]) +
	( 16'sd 32181) * $signed(input_fmap_47[15:0]) +
	( 14'sd 4543) * $signed(input_fmap_48[15:0]) +
	( 16'sd 20679) * $signed(input_fmap_49[15:0]) +
	( 16'sd 17509) * $signed(input_fmap_50[15:0]) +
	( 16'sd 22376) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19351) * $signed(input_fmap_52[15:0]) +
	( 16'sd 31365) * $signed(input_fmap_53[15:0]) +
	( 13'sd 2706) * $signed(input_fmap_54[15:0]) +
	( 15'sd 9838) * $signed(input_fmap_55[15:0]) +
	( 16'sd 29895) * $signed(input_fmap_56[15:0]) +
	( 16'sd 24352) * $signed(input_fmap_57[15:0]) +
	( 16'sd 19875) * $signed(input_fmap_58[15:0]) +
	( 16'sd 22374) * $signed(input_fmap_59[15:0]) +
	( 16'sd 17659) * $signed(input_fmap_60[15:0]) +
	( 16'sd 26255) * $signed(input_fmap_61[15:0]) +
	( 15'sd 16293) * $signed(input_fmap_62[15:0]) +
	( 14'sd 7069) * $signed(input_fmap_63[15:0]) +
	( 13'sd 3054) * $signed(input_fmap_64[15:0]) +
	( 14'sd 5913) * $signed(input_fmap_65[15:0]) +
	( 16'sd 18615) * $signed(input_fmap_66[15:0]) +
	( 16'sd 31566) * $signed(input_fmap_67[15:0]) +
	( 16'sd 17469) * $signed(input_fmap_68[15:0]) +
	( 16'sd 25129) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31501) * $signed(input_fmap_70[15:0]) +
	( 14'sd 6923) * $signed(input_fmap_71[15:0]) +
	( 12'sd 2032) * $signed(input_fmap_72[15:0]) +
	( 14'sd 4325) * $signed(input_fmap_73[15:0]) +
	( 15'sd 9067) * $signed(input_fmap_74[15:0]) +
	( 16'sd 19517) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19724) * $signed(input_fmap_76[15:0]) +
	( 16'sd 27366) * $signed(input_fmap_77[15:0]) +
	( 16'sd 20901) * $signed(input_fmap_78[15:0]) +
	( 15'sd 11338) * $signed(input_fmap_79[15:0]) +
	( 15'sd 14567) * $signed(input_fmap_80[15:0]) +
	( 15'sd 13274) * $signed(input_fmap_81[15:0]) +
	( 15'sd 15763) * $signed(input_fmap_82[15:0]) +
	( 14'sd 4953) * $signed(input_fmap_83[15:0]) +
	( 16'sd 16568) * $signed(input_fmap_84[15:0]) +
	( 16'sd 17106) * $signed(input_fmap_85[15:0]) +
	( 16'sd 32462) * $signed(input_fmap_86[15:0]) +
	( 15'sd 10906) * $signed(input_fmap_87[15:0]) +
	( 16'sd 25679) * $signed(input_fmap_88[15:0]) +
	( 15'sd 15650) * $signed(input_fmap_89[15:0]) +
	( 16'sd 22860) * $signed(input_fmap_90[15:0]) +
	( 14'sd 6863) * $signed(input_fmap_91[15:0]) +
	( 16'sd 20337) * $signed(input_fmap_92[15:0]) +
	( 15'sd 10159) * $signed(input_fmap_93[15:0]) +
	( 15'sd 11972) * $signed(input_fmap_94[15:0]) +
	( 16'sd 27209) * $signed(input_fmap_95[15:0]) +
	( 14'sd 6381) * $signed(input_fmap_96[15:0]) +
	( 16'sd 19053) * $signed(input_fmap_97[15:0]) +
	( 16'sd 24360) * $signed(input_fmap_98[15:0]) +
	( 13'sd 2703) * $signed(input_fmap_99[15:0]) +
	( 16'sd 26663) * $signed(input_fmap_100[15:0]) +
	( 16'sd 27742) * $signed(input_fmap_101[15:0]) +
	( 15'sd 8843) * $signed(input_fmap_102[15:0]) +
	( 16'sd 22657) * $signed(input_fmap_103[15:0]) +
	( 16'sd 19679) * $signed(input_fmap_104[15:0]) +
	( 16'sd 24765) * $signed(input_fmap_105[15:0]) +
	( 15'sd 16075) * $signed(input_fmap_106[15:0]) +
	( 15'sd 9837) * $signed(input_fmap_107[15:0]) +
	( 16'sd 28459) * $signed(input_fmap_108[15:0]) +
	( 15'sd 15029) * $signed(input_fmap_109[15:0]) +
	( 16'sd 18804) * $signed(input_fmap_110[15:0]) +
	( 16'sd 27215) * $signed(input_fmap_111[15:0]) +
	( 15'sd 10443) * $signed(input_fmap_112[15:0]) +
	( 16'sd 27326) * $signed(input_fmap_113[15:0]) +
	( 16'sd 17186) * $signed(input_fmap_114[15:0]) +
	( 16'sd 25852) * $signed(input_fmap_115[15:0]) +
	( 14'sd 7163) * $signed(input_fmap_116[15:0]) +
	( 14'sd 4919) * $signed(input_fmap_117[15:0]) +
	( 16'sd 18553) * $signed(input_fmap_118[15:0]) +
	( 16'sd 27719) * $signed(input_fmap_119[15:0]) +
	( 16'sd 30389) * $signed(input_fmap_120[15:0]) +
	( 15'sd 10906) * $signed(input_fmap_121[15:0]) +
	( 16'sd 16435) * $signed(input_fmap_122[15:0]) +
	( 16'sd 19113) * $signed(input_fmap_123[15:0]) +
	( 15'sd 8901) * $signed(input_fmap_124[15:0]) +
	( 16'sd 23869) * $signed(input_fmap_125[15:0]) +
	( 11'sd 703) * $signed(input_fmap_126[15:0]) +
	( 16'sd 23408) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 15'sd 12911) * $signed(input_fmap_0[15:0]) +
	( 16'sd 32574) * $signed(input_fmap_1[15:0]) +
	( 15'sd 12392) * $signed(input_fmap_2[15:0]) +
	( 15'sd 8280) * $signed(input_fmap_3[15:0]) +
	( 14'sd 6673) * $signed(input_fmap_4[15:0]) +
	( 15'sd 16341) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2886) * $signed(input_fmap_6[15:0]) +
	( 14'sd 5033) * $signed(input_fmap_7[15:0]) +
	( 14'sd 4406) * $signed(input_fmap_8[15:0]) +
	( 16'sd 23242) * $signed(input_fmap_9[15:0]) +
	( 16'sd 17013) * $signed(input_fmap_10[15:0]) +
	( 15'sd 12500) * $signed(input_fmap_11[15:0]) +
	( 14'sd 5094) * $signed(input_fmap_12[15:0]) +
	( 15'sd 10566) * $signed(input_fmap_13[15:0]) +
	( 16'sd 28211) * $signed(input_fmap_14[15:0]) +
	( 16'sd 30648) * $signed(input_fmap_15[15:0]) +
	( 15'sd 11333) * $signed(input_fmap_16[15:0]) +
	( 16'sd 29785) * $signed(input_fmap_17[15:0]) +
	( 14'sd 6994) * $signed(input_fmap_18[15:0]) +
	( 16'sd 22010) * $signed(input_fmap_19[15:0]) +
	( 16'sd 25619) * $signed(input_fmap_20[15:0]) +
	( 14'sd 6398) * $signed(input_fmap_21[15:0]) +
	( 14'sd 6381) * $signed(input_fmap_22[15:0]) +
	( 16'sd 20330) * $signed(input_fmap_23[15:0]) +
	( 16'sd 23065) * $signed(input_fmap_24[15:0]) +
	( 16'sd 30112) * $signed(input_fmap_25[15:0]) +
	( 15'sd 15837) * $signed(input_fmap_26[15:0]) +
	( 16'sd 16659) * $signed(input_fmap_27[15:0]) +
	( 16'sd 23748) * $signed(input_fmap_28[15:0]) +
	( 15'sd 15986) * $signed(input_fmap_29[15:0]) +
	( 14'sd 7299) * $signed(input_fmap_30[15:0]) +
	( 15'sd 8871) * $signed(input_fmap_31[15:0]) +
	( 14'sd 5272) * $signed(input_fmap_32[15:0]) +
	( 12'sd 1220) * $signed(input_fmap_33[15:0]) +
	( 16'sd 20435) * $signed(input_fmap_34[15:0]) +
	( 16'sd 19286) * $signed(input_fmap_35[15:0]) +
	( 16'sd 30810) * $signed(input_fmap_36[15:0]) +
	( 16'sd 22066) * $signed(input_fmap_37[15:0]) +
	( 16'sd 19331) * $signed(input_fmap_38[15:0]) +
	( 16'sd 28073) * $signed(input_fmap_39[15:0]) +
	( 15'sd 15121) * $signed(input_fmap_40[15:0]) +
	( 16'sd 29072) * $signed(input_fmap_41[15:0]) +
	( 15'sd 12058) * $signed(input_fmap_42[15:0]) +
	( 16'sd 20071) * $signed(input_fmap_43[15:0]) +
	( 16'sd 17651) * $signed(input_fmap_44[15:0]) +
	( 12'sd 1606) * $signed(input_fmap_45[15:0]) +
	( 15'sd 8453) * $signed(input_fmap_46[15:0]) +
	( 15'sd 8405) * $signed(input_fmap_47[15:0]) +
	( 16'sd 29694) * $signed(input_fmap_48[15:0]) +
	( 15'sd 15548) * $signed(input_fmap_49[15:0]) +
	( 12'sd 1759) * $signed(input_fmap_50[15:0]) +
	( 16'sd 30714) * $signed(input_fmap_51[15:0]) +
	( 10'sd 503) * $signed(input_fmap_52[15:0]) +
	( 16'sd 22949) * $signed(input_fmap_53[15:0]) +
	( 16'sd 25056) * $signed(input_fmap_54[15:0]) +
	( 16'sd 17423) * $signed(input_fmap_55[15:0]) +
	( 15'sd 12043) * $signed(input_fmap_56[15:0]) +
	( 16'sd 32436) * $signed(input_fmap_57[15:0]) +
	( 11'sd 646) * $signed(input_fmap_58[15:0]) +
	( 16'sd 18283) * $signed(input_fmap_59[15:0]) +
	( 16'sd 18479) * $signed(input_fmap_60[15:0]) +
	( 15'sd 8896) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3665) * $signed(input_fmap_62[15:0]) +
	( 13'sd 2556) * $signed(input_fmap_63[15:0]) +
	( 16'sd 17862) * $signed(input_fmap_64[15:0]) +
	( 15'sd 12549) * $signed(input_fmap_65[15:0]) +
	( 16'sd 23240) * $signed(input_fmap_66[15:0]) +
	( 16'sd 18072) * $signed(input_fmap_67[15:0]) +
	( 15'sd 13999) * $signed(input_fmap_68[15:0]) +
	( 15'sd 11333) * $signed(input_fmap_69[15:0]) +
	( 16'sd 32289) * $signed(input_fmap_70[15:0]) +
	( 10'sd 338) * $signed(input_fmap_71[15:0]) +
	( 15'sd 9148) * $signed(input_fmap_72[15:0]) +
	( 14'sd 6700) * $signed(input_fmap_73[15:0]) +
	( 13'sd 2664) * $signed(input_fmap_74[15:0]) +
	( 15'sd 9903) * $signed(input_fmap_75[15:0]) +
	( 14'sd 5447) * $signed(input_fmap_76[15:0]) +
	( 14'sd 5915) * $signed(input_fmap_77[15:0]) +
	( 16'sd 30128) * $signed(input_fmap_78[15:0]) +
	( 12'sd 1832) * $signed(input_fmap_79[15:0]) +
	( 16'sd 31502) * $signed(input_fmap_80[15:0]) +
	( 16'sd 23527) * $signed(input_fmap_81[15:0]) +
	( 14'sd 5459) * $signed(input_fmap_82[15:0]) +
	( 11'sd 803) * $signed(input_fmap_83[15:0]) +
	( 16'sd 21764) * $signed(input_fmap_84[15:0]) +
	( 14'sd 4682) * $signed(input_fmap_85[15:0]) +
	( 16'sd 18020) * $signed(input_fmap_86[15:0]) +
	( 16'sd 16864) * $signed(input_fmap_87[15:0]) +
	( 14'sd 4200) * $signed(input_fmap_88[15:0]) +
	( 16'sd 24048) * $signed(input_fmap_89[15:0]) +
	( 13'sd 2230) * $signed(input_fmap_90[15:0]) +
	( 16'sd 25352) * $signed(input_fmap_91[15:0]) +
	( 15'sd 10458) * $signed(input_fmap_92[15:0]) +
	( 15'sd 15204) * $signed(input_fmap_93[15:0]) +
	( 14'sd 7681) * $signed(input_fmap_94[15:0]) +
	( 16'sd 24521) * $signed(input_fmap_95[15:0]) +
	( 15'sd 14065) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27586) * $signed(input_fmap_97[15:0]) +
	( 13'sd 2926) * $signed(input_fmap_98[15:0]) +
	( 13'sd 2111) * $signed(input_fmap_99[15:0]) +
	( 16'sd 25104) * $signed(input_fmap_100[15:0]) +
	( 16'sd 16650) * $signed(input_fmap_101[15:0]) +
	( 16'sd 17374) * $signed(input_fmap_102[15:0]) +
	( 15'sd 10595) * $signed(input_fmap_103[15:0]) +
	( 16'sd 27842) * $signed(input_fmap_104[15:0]) +
	( 16'sd 24036) * $signed(input_fmap_105[15:0]) +
	( 15'sd 11646) * $signed(input_fmap_106[15:0]) +
	( 16'sd 21486) * $signed(input_fmap_107[15:0]) +
	( 15'sd 9058) * $signed(input_fmap_108[15:0]) +
	( 15'sd 13538) * $signed(input_fmap_109[15:0]) +
	( 15'sd 12131) * $signed(input_fmap_110[15:0]) +
	( 15'sd 13317) * $signed(input_fmap_111[15:0]) +
	( 13'sd 4072) * $signed(input_fmap_112[15:0]) +
	( 16'sd 24080) * $signed(input_fmap_113[15:0]) +
	( 16'sd 27682) * $signed(input_fmap_114[15:0]) +
	( 16'sd 20523) * $signed(input_fmap_115[15:0]) +
	( 15'sd 14413) * $signed(input_fmap_116[15:0]) +
	( 16'sd 19493) * $signed(input_fmap_117[15:0]) +
	( 16'sd 23654) * $signed(input_fmap_118[15:0]) +
	( 14'sd 7373) * $signed(input_fmap_119[15:0]) +
	( 16'sd 29626) * $signed(input_fmap_120[15:0]) +
	( 16'sd 24231) * $signed(input_fmap_121[15:0]) +
	( 16'sd 30474) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21512) * $signed(input_fmap_123[15:0]) +
	( 16'sd 29704) * $signed(input_fmap_124[15:0]) +
	( 12'sd 1151) * $signed(input_fmap_125[15:0]) +
	( 16'sd 26123) * $signed(input_fmap_126[15:0]) +
	( 15'sd 15764) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 15'sd 12990) * $signed(input_fmap_0[15:0]) +
	( 16'sd 20306) * $signed(input_fmap_1[15:0]) +
	( 14'sd 4748) * $signed(input_fmap_2[15:0]) +
	( 16'sd 17874) * $signed(input_fmap_3[15:0]) +
	( 14'sd 5826) * $signed(input_fmap_4[15:0]) +
	( 15'sd 10571) * $signed(input_fmap_5[15:0]) +
	( 15'sd 8535) * $signed(input_fmap_6[15:0]) +
	( 15'sd 9709) * $signed(input_fmap_7[15:0]) +
	( 16'sd 16514) * $signed(input_fmap_8[15:0]) +
	( 16'sd 28855) * $signed(input_fmap_9[15:0]) +
	( 16'sd 16690) * $signed(input_fmap_10[15:0]) +
	( 14'sd 7853) * $signed(input_fmap_11[15:0]) +
	( 16'sd 17317) * $signed(input_fmap_12[15:0]) +
	( 16'sd 26720) * $signed(input_fmap_13[15:0]) +
	( 16'sd 20875) * $signed(input_fmap_14[15:0]) +
	( 16'sd 27967) * $signed(input_fmap_15[15:0]) +
	( 11'sd 997) * $signed(input_fmap_16[15:0]) +
	( 16'sd 27696) * $signed(input_fmap_17[15:0]) +
	( 15'sd 14734) * $signed(input_fmap_18[15:0]) +
	( 16'sd 29598) * $signed(input_fmap_19[15:0]) +
	( 13'sd 2239) * $signed(input_fmap_20[15:0]) +
	( 16'sd 21723) * $signed(input_fmap_21[15:0]) +
	( 16'sd 27436) * $signed(input_fmap_22[15:0]) +
	( 16'sd 18801) * $signed(input_fmap_23[15:0]) +
	( 15'sd 10722) * $signed(input_fmap_24[15:0]) +
	( 16'sd 27292) * $signed(input_fmap_25[15:0]) +
	( 13'sd 3661) * $signed(input_fmap_26[15:0]) +
	( 16'sd 31600) * $signed(input_fmap_27[15:0]) +
	( 15'sd 13301) * $signed(input_fmap_28[15:0]) +
	( 16'sd 16737) * $signed(input_fmap_29[15:0]) +
	( 16'sd 18790) * $signed(input_fmap_30[15:0]) +
	( 15'sd 11170) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28420) * $signed(input_fmap_32[15:0]) +
	( 16'sd 29556) * $signed(input_fmap_33[15:0]) +
	( 16'sd 17313) * $signed(input_fmap_34[15:0]) +
	( 16'sd 25077) * $signed(input_fmap_35[15:0]) +
	( 14'sd 6012) * $signed(input_fmap_36[15:0]) +
	( 14'sd 4238) * $signed(input_fmap_37[15:0]) +
	( 14'sd 4765) * $signed(input_fmap_38[15:0]) +
	( 16'sd 31320) * $signed(input_fmap_39[15:0]) +
	( 15'sd 15327) * $signed(input_fmap_40[15:0]) +
	( 15'sd 14250) * $signed(input_fmap_41[15:0]) +
	( 15'sd 10022) * $signed(input_fmap_42[15:0]) +
	( 15'sd 12023) * $signed(input_fmap_43[15:0]) +
	( 16'sd 26138) * $signed(input_fmap_44[15:0]) +
	( 16'sd 20491) * $signed(input_fmap_45[15:0]) +
	( 16'sd 22130) * $signed(input_fmap_46[15:0]) +
	( 14'sd 5805) * $signed(input_fmap_47[15:0]) +
	( 16'sd 26426) * $signed(input_fmap_48[15:0]) +
	( 16'sd 16941) * $signed(input_fmap_49[15:0]) +
	( 15'sd 15717) * $signed(input_fmap_50[15:0]) +
	( 13'sd 3112) * $signed(input_fmap_51[15:0]) +
	( 15'sd 12272) * $signed(input_fmap_52[15:0]) +
	( 14'sd 4535) * $signed(input_fmap_53[15:0]) +
	( 16'sd 19125) * $signed(input_fmap_54[15:0]) +
	( 15'sd 13623) * $signed(input_fmap_55[15:0]) +
	( 15'sd 8674) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17592) * $signed(input_fmap_57[15:0]) +
	( 14'sd 5244) * $signed(input_fmap_58[15:0]) +
	( 16'sd 29143) * $signed(input_fmap_59[15:0]) +
	( 16'sd 21917) * $signed(input_fmap_60[15:0]) +
	( 13'sd 2653) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29264) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20138) * $signed(input_fmap_63[15:0]) +
	( 15'sd 15655) * $signed(input_fmap_64[15:0]) +
	( 16'sd 27869) * $signed(input_fmap_65[15:0]) +
	( 16'sd 31241) * $signed(input_fmap_66[15:0]) +
	( 16'sd 23089) * $signed(input_fmap_67[15:0]) +
	( 16'sd 23720) * $signed(input_fmap_68[15:0]) +
	( 15'sd 13174) * $signed(input_fmap_69[15:0]) +
	( 15'sd 11374) * $signed(input_fmap_70[15:0]) +
	( 12'sd 1422) * $signed(input_fmap_71[15:0]) +
	( 12'sd 1566) * $signed(input_fmap_72[15:0]) +
	( 16'sd 22595) * $signed(input_fmap_73[15:0]) +
	( 15'sd 15523) * $signed(input_fmap_74[15:0]) +
	( 15'sd 16243) * $signed(input_fmap_75[15:0]) +
	( 15'sd 12251) * $signed(input_fmap_76[15:0]) +
	( 16'sd 30363) * $signed(input_fmap_77[15:0]) +
	( 16'sd 28575) * $signed(input_fmap_78[15:0]) +
	( 16'sd 24854) * $signed(input_fmap_79[15:0]) +
	( 16'sd 29038) * $signed(input_fmap_80[15:0]) +
	( 16'sd 18913) * $signed(input_fmap_81[15:0]) +
	( 15'sd 12918) * $signed(input_fmap_82[15:0]) +
	( 12'sd 1943) * $signed(input_fmap_83[15:0]) +
	( 15'sd 13485) * $signed(input_fmap_84[15:0]) +
	( 16'sd 16590) * $signed(input_fmap_85[15:0]) +
	( 16'sd 16441) * $signed(input_fmap_86[15:0]) +
	( 15'sd 10282) * $signed(input_fmap_87[15:0]) +
	( 16'sd 26130) * $signed(input_fmap_88[15:0]) +
	( 15'sd 9552) * $signed(input_fmap_89[15:0]) +
	( 15'sd 16173) * $signed(input_fmap_90[15:0]) +
	( 16'sd 29160) * $signed(input_fmap_91[15:0]) +
	( 14'sd 7722) * $signed(input_fmap_92[15:0]) +
	( 16'sd 21923) * $signed(input_fmap_93[15:0]) +
	( 14'sd 5947) * $signed(input_fmap_94[15:0]) +
	( 12'sd 1915) * $signed(input_fmap_95[15:0]) +
	( 15'sd 14841) * $signed(input_fmap_96[15:0]) +
	( 15'sd 8503) * $signed(input_fmap_97[15:0]) +
	( 15'sd 10798) * $signed(input_fmap_98[15:0]) +
	( 15'sd 9826) * $signed(input_fmap_99[15:0]) +
	( 16'sd 29859) * $signed(input_fmap_100[15:0]) +
	( 15'sd 13740) * $signed(input_fmap_101[15:0]) +
	( 15'sd 10925) * $signed(input_fmap_102[15:0]) +
	( 14'sd 6148) * $signed(input_fmap_103[15:0]) +
	( 14'sd 7397) * $signed(input_fmap_104[15:0]) +
	( 13'sd 2744) * $signed(input_fmap_105[15:0]) +
	( 16'sd 27169) * $signed(input_fmap_106[15:0]) +
	( 11'sd 945) * $signed(input_fmap_107[15:0]) +
	( 16'sd 24908) * $signed(input_fmap_108[15:0]) +
	( 16'sd 32295) * $signed(input_fmap_109[15:0]) +
	( 14'sd 7410) * $signed(input_fmap_110[15:0]) +
	( 14'sd 7289) * $signed(input_fmap_111[15:0]) +
	( 13'sd 2441) * $signed(input_fmap_112[15:0]) +
	( 15'sd 10726) * $signed(input_fmap_113[15:0]) +
	( 14'sd 4629) * $signed(input_fmap_114[15:0]) +
	( 13'sd 2887) * $signed(input_fmap_115[15:0]) +
	( 16'sd 27070) * $signed(input_fmap_116[15:0]) +
	( 16'sd 25802) * $signed(input_fmap_117[15:0]) +
	( 15'sd 11429) * $signed(input_fmap_118[15:0]) +
	( 16'sd 17489) * $signed(input_fmap_119[15:0]) +
	( 15'sd 9451) * $signed(input_fmap_120[15:0]) +
	( 15'sd 9949) * $signed(input_fmap_121[15:0]) +
	( 16'sd 29332) * $signed(input_fmap_122[15:0]) +
	( 12'sd 1086) * $signed(input_fmap_123[15:0]) +
	( 16'sd 28231) * $signed(input_fmap_124[15:0]) +
	( 16'sd 23833) * $signed(input_fmap_125[15:0]) +
	( 13'sd 3710) * $signed(input_fmap_126[15:0]) +
	( 15'sd 13935) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 16'sd 26606) * $signed(input_fmap_0[15:0]) +
	( 16'sd 22187) * $signed(input_fmap_1[15:0]) +
	( 16'sd 17384) * $signed(input_fmap_2[15:0]) +
	( 16'sd 26032) * $signed(input_fmap_3[15:0]) +
	( 15'sd 8227) * $signed(input_fmap_4[15:0]) +
	( 16'sd 24503) * $signed(input_fmap_5[15:0]) +
	( 15'sd 14035) * $signed(input_fmap_6[15:0]) +
	( 13'sd 2747) * $signed(input_fmap_7[15:0]) +
	( 16'sd 28278) * $signed(input_fmap_8[15:0]) +
	( 14'sd 5604) * $signed(input_fmap_9[15:0]) +
	( 14'sd 5475) * $signed(input_fmap_10[15:0]) +
	( 16'sd 19408) * $signed(input_fmap_11[15:0]) +
	( 14'sd 7496) * $signed(input_fmap_12[15:0]) +
	( 16'sd 23678) * $signed(input_fmap_13[15:0]) +
	( 16'sd 31932) * $signed(input_fmap_14[15:0]) +
	( 14'sd 6084) * $signed(input_fmap_15[15:0]) +
	( 15'sd 14947) * $signed(input_fmap_16[15:0]) +
	( 11'sd 746) * $signed(input_fmap_17[15:0]) +
	( 13'sd 2419) * $signed(input_fmap_18[15:0]) +
	( 16'sd 31331) * $signed(input_fmap_19[15:0]) +
	( 13'sd 4053) * $signed(input_fmap_20[15:0]) +
	( 16'sd 18270) * $signed(input_fmap_21[15:0]) +
	( 16'sd 22165) * $signed(input_fmap_22[15:0]) +
	( 13'sd 3433) * $signed(input_fmap_23[15:0]) +
	( 16'sd 19657) * $signed(input_fmap_24[15:0]) +
	( 15'sd 15295) * $signed(input_fmap_25[15:0]) +
	( 14'sd 6028) * $signed(input_fmap_26[15:0]) +
	( 10'sd 320) * $signed(input_fmap_27[15:0]) +
	( 13'sd 4033) * $signed(input_fmap_28[15:0]) +
	( 16'sd 22837) * $signed(input_fmap_29[15:0]) +
	( 16'sd 22431) * $signed(input_fmap_30[15:0]) +
	( 16'sd 28696) * $signed(input_fmap_31[15:0]) +
	( 16'sd 30501) * $signed(input_fmap_32[15:0]) +
	( 15'sd 14674) * $signed(input_fmap_33[15:0]) +
	( 15'sd 12742) * $signed(input_fmap_34[15:0]) +
	( 16'sd 27732) * $signed(input_fmap_35[15:0]) +
	( 15'sd 13039) * $signed(input_fmap_36[15:0]) +
	( 14'sd 6452) * $signed(input_fmap_37[15:0]) +
	( 16'sd 31591) * $signed(input_fmap_38[15:0]) +
	( 16'sd 26448) * $signed(input_fmap_39[15:0]) +
	( 12'sd 1541) * $signed(input_fmap_40[15:0]) +
	( 11'sd 738) * $signed(input_fmap_41[15:0]) +
	( 16'sd 27261) * $signed(input_fmap_42[15:0]) +
	( 15'sd 10115) * $signed(input_fmap_43[15:0]) +
	( 16'sd 20196) * $signed(input_fmap_44[15:0]) +
	( 14'sd 7625) * $signed(input_fmap_45[15:0]) +
	( 15'sd 14980) * $signed(input_fmap_46[15:0]) +
	( 16'sd 17301) * $signed(input_fmap_47[15:0]) +
	( 16'sd 18804) * $signed(input_fmap_48[15:0]) +
	( 16'sd 19886) * $signed(input_fmap_49[15:0]) +
	( 16'sd 17164) * $signed(input_fmap_50[15:0]) +
	( 16'sd 27703) * $signed(input_fmap_51[15:0]) +
	( 16'sd 31372) * $signed(input_fmap_52[15:0]) +
	( 15'sd 12735) * $signed(input_fmap_53[15:0]) +
	( 16'sd 26706) * $signed(input_fmap_54[15:0]) +
	( 15'sd 12279) * $signed(input_fmap_55[15:0]) +
	( 14'sd 4760) * $signed(input_fmap_56[15:0]) +
	( 16'sd 20287) * $signed(input_fmap_57[15:0]) +
	( 15'sd 15289) * $signed(input_fmap_58[15:0]) +
	( 16'sd 24787) * $signed(input_fmap_59[15:0]) +
	( 16'sd 24399) * $signed(input_fmap_60[15:0]) +
	( 10'sd 404) * $signed(input_fmap_61[15:0]) +
	( 16'sd 31442) * $signed(input_fmap_62[15:0]) +
	( 15'sd 11476) * $signed(input_fmap_63[15:0]) +
	( 16'sd 31951) * $signed(input_fmap_64[15:0]) +
	( 16'sd 31969) * $signed(input_fmap_65[15:0]) +
	( 16'sd 28486) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28291) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26233) * $signed(input_fmap_68[15:0]) +
	( 15'sd 12840) * $signed(input_fmap_69[15:0]) +
	( 15'sd 15988) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11360) * $signed(input_fmap_71[15:0]) +
	( 16'sd 20359) * $signed(input_fmap_72[15:0]) +
	( 16'sd 21738) * $signed(input_fmap_73[15:0]) +
	( 10'sd 310) * $signed(input_fmap_74[15:0]) +
	( 15'sd 15283) * $signed(input_fmap_75[15:0]) +
	( 15'sd 11694) * $signed(input_fmap_76[15:0]) +
	( 15'sd 11819) * $signed(input_fmap_77[15:0]) +
	( 15'sd 11505) * $signed(input_fmap_78[15:0]) +
	( 15'sd 12007) * $signed(input_fmap_79[15:0]) +
	( 15'sd 11736) * $signed(input_fmap_80[15:0]) +
	( 14'sd 6050) * $signed(input_fmap_81[15:0]) +
	( 15'sd 9856) * $signed(input_fmap_82[15:0]) +
	( 16'sd 30663) * $signed(input_fmap_83[15:0]) +
	( 14'sd 5413) * $signed(input_fmap_84[15:0]) +
	( 15'sd 8411) * $signed(input_fmap_85[15:0]) +
	( 15'sd 15889) * $signed(input_fmap_86[15:0]) +
	( 13'sd 3097) * $signed(input_fmap_87[15:0]) +
	( 15'sd 11279) * $signed(input_fmap_88[15:0]) +
	( 16'sd 29748) * $signed(input_fmap_89[15:0]) +
	( 14'sd 7024) * $signed(input_fmap_90[15:0]) +
	( 14'sd 5056) * $signed(input_fmap_91[15:0]) +
	( 15'sd 13992) * $signed(input_fmap_92[15:0]) +
	( 11'sd 660) * $signed(input_fmap_93[15:0]) +
	( 13'sd 3178) * $signed(input_fmap_94[15:0]) +
	( 15'sd 15154) * $signed(input_fmap_95[15:0]) +
	( 14'sd 5231) * $signed(input_fmap_96[15:0]) +
	( 16'sd 26122) * $signed(input_fmap_97[15:0]) +
	( 11'sd 589) * $signed(input_fmap_98[15:0]) +
	( 14'sd 7086) * $signed(input_fmap_99[15:0]) +
	( 15'sd 11576) * $signed(input_fmap_100[15:0]) +
	( 14'sd 4389) * $signed(input_fmap_101[15:0]) +
	( 16'sd 24058) * $signed(input_fmap_102[15:0]) +
	( 16'sd 20546) * $signed(input_fmap_103[15:0]) +
	( 16'sd 26884) * $signed(input_fmap_104[15:0]) +
	( 15'sd 10052) * $signed(input_fmap_105[15:0]) +
	( 12'sd 1130) * $signed(input_fmap_106[15:0]) +
	( 16'sd 28725) * $signed(input_fmap_107[15:0]) +
	( 15'sd 13468) * $signed(input_fmap_108[15:0]) +
	( 16'sd 16555) * $signed(input_fmap_109[15:0]) +
	( 14'sd 6922) * $signed(input_fmap_110[15:0]) +
	( 14'sd 6804) * $signed(input_fmap_111[15:0]) +
	( 14'sd 7807) * $signed(input_fmap_112[15:0]) +
	( 16'sd 28349) * $signed(input_fmap_113[15:0]) +
	( 15'sd 9652) * $signed(input_fmap_114[15:0]) +
	( 16'sd 24811) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26692) * $signed(input_fmap_116[15:0]) +
	( 16'sd 30825) * $signed(input_fmap_117[15:0]) +
	( 15'sd 8915) * $signed(input_fmap_118[15:0]) +
	( 15'sd 10858) * $signed(input_fmap_119[15:0]) +
	( 15'sd 16160) * $signed(input_fmap_120[15:0]) +
	( 15'sd 16300) * $signed(input_fmap_121[15:0]) +
	( 16'sd 18436) * $signed(input_fmap_122[15:0]) +
	( 16'sd 32720) * $signed(input_fmap_123[15:0]) +
	( 16'sd 27250) * $signed(input_fmap_124[15:0]) +
	( 14'sd 4537) * $signed(input_fmap_125[15:0]) +
	( 16'sd 25751) * $signed(input_fmap_126[15:0]) +
	( 14'sd 4717) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 16'sd 27885) * $signed(input_fmap_0[15:0]) +
	( 15'sd 12856) * $signed(input_fmap_1[15:0]) +
	( 15'sd 9332) * $signed(input_fmap_2[15:0]) +
	( 16'sd 20541) * $signed(input_fmap_3[15:0]) +
	( 16'sd 27246) * $signed(input_fmap_4[15:0]) +
	( 14'sd 8015) * $signed(input_fmap_5[15:0]) +
	( 16'sd 31620) * $signed(input_fmap_6[15:0]) +
	( 15'sd 9832) * $signed(input_fmap_7[15:0]) +
	( 15'sd 11120) * $signed(input_fmap_8[15:0]) +
	( 16'sd 18064) * $signed(input_fmap_9[15:0]) +
	( 14'sd 6202) * $signed(input_fmap_10[15:0]) +
	( 16'sd 21377) * $signed(input_fmap_11[15:0]) +
	( 15'sd 11018) * $signed(input_fmap_12[15:0]) +
	( 15'sd 14170) * $signed(input_fmap_13[15:0]) +
	( 16'sd 17912) * $signed(input_fmap_14[15:0]) +
	( 16'sd 24821) * $signed(input_fmap_15[15:0]) +
	( 16'sd 28186) * $signed(input_fmap_16[15:0]) +
	( 13'sd 2872) * $signed(input_fmap_17[15:0]) +
	( 14'sd 4145) * $signed(input_fmap_18[15:0]) +
	( 16'sd 22083) * $signed(input_fmap_19[15:0]) +
	( 14'sd 6328) * $signed(input_fmap_20[15:0]) +
	( 16'sd 25593) * $signed(input_fmap_21[15:0]) +
	( 14'sd 7839) * $signed(input_fmap_22[15:0]) +
	( 14'sd 4495) * $signed(input_fmap_23[15:0]) +
	( 14'sd 6232) * $signed(input_fmap_24[15:0]) +
	( 16'sd 30722) * $signed(input_fmap_25[15:0]) +
	( 16'sd 25399) * $signed(input_fmap_26[15:0]) +
	( 16'sd 22827) * $signed(input_fmap_27[15:0]) +
	( 16'sd 17812) * $signed(input_fmap_28[15:0]) +
	( 14'sd 5125) * $signed(input_fmap_29[15:0]) +
	( 14'sd 8029) * $signed(input_fmap_30[15:0]) +
	( 13'sd 3205) * $signed(input_fmap_31[15:0]) +
	( 13'sd 3806) * $signed(input_fmap_32[15:0]) +
	( 16'sd 26547) * $signed(input_fmap_33[15:0]) +
	( 16'sd 29809) * $signed(input_fmap_34[15:0]) +
	( 14'sd 7640) * $signed(input_fmap_35[15:0]) +
	( 16'sd 18829) * $signed(input_fmap_36[15:0]) +
	( 16'sd 25341) * $signed(input_fmap_37[15:0]) +
	( 16'sd 19150) * $signed(input_fmap_38[15:0]) +
	( 16'sd 20526) * $signed(input_fmap_39[15:0]) +
	( 16'sd 30722) * $signed(input_fmap_40[15:0]) +
	( 16'sd 23086) * $signed(input_fmap_41[15:0]) +
	( 14'sd 5250) * $signed(input_fmap_42[15:0]) +
	( 14'sd 4471) * $signed(input_fmap_43[15:0]) +
	( 14'sd 6383) * $signed(input_fmap_44[15:0]) +
	( 13'sd 2052) * $signed(input_fmap_45[15:0]) +
	( 15'sd 14050) * $signed(input_fmap_46[15:0]) +
	( 15'sd 14374) * $signed(input_fmap_47[15:0]) +
	( 16'sd 27811) * $signed(input_fmap_48[15:0]) +
	( 14'sd 6529) * $signed(input_fmap_49[15:0]) +
	( 15'sd 10364) * $signed(input_fmap_50[15:0]) +
	( 15'sd 9639) * $signed(input_fmap_51[15:0]) +
	( 16'sd 32215) * $signed(input_fmap_52[15:0]) +
	( 16'sd 22471) * $signed(input_fmap_53[15:0]) +
	( 16'sd 18958) * $signed(input_fmap_54[15:0]) +
	( 16'sd 22794) * $signed(input_fmap_55[15:0]) +
	( 16'sd 32408) * $signed(input_fmap_56[15:0]) +
	( 16'sd 27998) * $signed(input_fmap_57[15:0]) +
	( 14'sd 7889) * $signed(input_fmap_58[15:0]) +
	( 15'sd 16110) * $signed(input_fmap_59[15:0]) +
	( 11'sd 896) * $signed(input_fmap_60[15:0]) +
	( 16'sd 32244) * $signed(input_fmap_61[15:0]) +
	( 16'sd 22417) * $signed(input_fmap_62[15:0]) +
	( 16'sd 19882) * $signed(input_fmap_63[15:0]) +
	( 16'sd 20966) * $signed(input_fmap_64[15:0]) +
	( 16'sd 29709) * $signed(input_fmap_65[15:0]) +
	( 16'sd 16933) * $signed(input_fmap_66[15:0]) +
	( 12'sd 1195) * $signed(input_fmap_67[15:0]) +
	( 13'sd 2286) * $signed(input_fmap_68[15:0]) +
	( 15'sd 8745) * $signed(input_fmap_69[15:0]) +
	( 13'sd 3022) * $signed(input_fmap_70[15:0]) +
	( 12'sd 1775) * $signed(input_fmap_71[15:0]) +
	( 16'sd 25334) * $signed(input_fmap_72[15:0]) +
	( 16'sd 30409) * $signed(input_fmap_73[15:0]) +
	( 12'sd 1684) * $signed(input_fmap_74[15:0]) +
	( 15'sd 11819) * $signed(input_fmap_75[15:0]) +
	( 16'sd 17533) * $signed(input_fmap_76[15:0]) +
	( 15'sd 14569) * $signed(input_fmap_77[15:0]) +
	( 15'sd 12795) * $signed(input_fmap_78[15:0]) +
	( 16'sd 22004) * $signed(input_fmap_79[15:0]) +
	( 16'sd 19575) * $signed(input_fmap_80[15:0]) +
	( 16'sd 25946) * $signed(input_fmap_81[15:0]) +
	( 15'sd 11972) * $signed(input_fmap_82[15:0]) +
	( 16'sd 32022) * $signed(input_fmap_83[15:0]) +
	( 16'sd 28084) * $signed(input_fmap_84[15:0]) +
	( 16'sd 27577) * $signed(input_fmap_85[15:0]) +
	( 15'sd 14841) * $signed(input_fmap_86[15:0]) +
	( 16'sd 24379) * $signed(input_fmap_87[15:0]) +
	( 16'sd 25291) * $signed(input_fmap_88[15:0]) +
	( 16'sd 17342) * $signed(input_fmap_89[15:0]) +
	( 13'sd 3833) * $signed(input_fmap_90[15:0]) +
	( 15'sd 8946) * $signed(input_fmap_91[15:0]) +
	( 14'sd 7618) * $signed(input_fmap_92[15:0]) +
	( 8'sd 97) * $signed(input_fmap_93[15:0]) +
	( 16'sd 17701) * $signed(input_fmap_94[15:0]) +
	( 16'sd 32129) * $signed(input_fmap_95[15:0]) +
	( 16'sd 16780) * $signed(input_fmap_96[15:0]) +
	( 12'sd 1512) * $signed(input_fmap_97[15:0]) +
	( 15'sd 14237) * $signed(input_fmap_98[15:0]) +
	( 11'sd 874) * $signed(input_fmap_99[15:0]) +
	( 16'sd 28514) * $signed(input_fmap_100[15:0]) +
	( 16'sd 18042) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5071) * $signed(input_fmap_102[15:0]) +
	( 11'sd 621) * $signed(input_fmap_103[15:0]) +
	( 16'sd 31453) * $signed(input_fmap_104[15:0]) +
	( 13'sd 3729) * $signed(input_fmap_105[15:0]) +
	( 13'sd 2105) * $signed(input_fmap_106[15:0]) +
	( 16'sd 26074) * $signed(input_fmap_107[15:0]) +
	( 16'sd 21681) * $signed(input_fmap_108[15:0]) +
	( 16'sd 30064) * $signed(input_fmap_109[15:0]) +
	( 15'sd 11657) * $signed(input_fmap_110[15:0]) +
	( 15'sd 12648) * $signed(input_fmap_111[15:0]) +
	( 14'sd 6922) * $signed(input_fmap_112[15:0]) +
	( 16'sd 22301) * $signed(input_fmap_113[15:0]) +
	( 16'sd 21428) * $signed(input_fmap_114[15:0]) +
	( 12'sd 1118) * $signed(input_fmap_115[15:0]) +
	( 13'sd 2776) * $signed(input_fmap_116[15:0]) +
	( 13'sd 3863) * $signed(input_fmap_117[15:0]) +
	( 16'sd 18411) * $signed(input_fmap_118[15:0]) +
	( 15'sd 9997) * $signed(input_fmap_119[15:0]) +
	( 16'sd 17121) * $signed(input_fmap_120[15:0]) +
	( 13'sd 2789) * $signed(input_fmap_121[15:0]) +
	( 15'sd 11172) * $signed(input_fmap_122[15:0]) +
	( 16'sd 16610) * $signed(input_fmap_123[15:0]) +
	( 16'sd 20960) * $signed(input_fmap_124[15:0]) +
	( 15'sd 13032) * $signed(input_fmap_125[15:0]) +
	( 14'sd 5838) * $signed(input_fmap_126[15:0]) +
	( 16'sd 23887) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 16'sd 25056) * $signed(input_fmap_0[15:0]) +
	( 15'sd 14744) * $signed(input_fmap_1[15:0]) +
	( 15'sd 11293) * $signed(input_fmap_2[15:0]) +
	( 14'sd 5491) * $signed(input_fmap_3[15:0]) +
	( 14'sd 6741) * $signed(input_fmap_4[15:0]) +
	( 16'sd 22235) * $signed(input_fmap_5[15:0]) +
	( 16'sd 23492) * $signed(input_fmap_6[15:0]) +
	( 16'sd 24692) * $signed(input_fmap_7[15:0]) +
	( 16'sd 29046) * $signed(input_fmap_8[15:0]) +
	( 15'sd 8739) * $signed(input_fmap_9[15:0]) +
	( 16'sd 21442) * $signed(input_fmap_10[15:0]) +
	( 16'sd 25276) * $signed(input_fmap_11[15:0]) +
	( 14'sd 4433) * $signed(input_fmap_12[15:0]) +
	( 16'sd 30953) * $signed(input_fmap_13[15:0]) +
	( 14'sd 5208) * $signed(input_fmap_14[15:0]) +
	( 16'sd 16727) * $signed(input_fmap_15[15:0]) +
	( 16'sd 27916) * $signed(input_fmap_16[15:0]) +
	( 16'sd 26201) * $signed(input_fmap_17[15:0]) +
	( 15'sd 11468) * $signed(input_fmap_18[15:0]) +
	( 16'sd 26796) * $signed(input_fmap_19[15:0]) +
	( 14'sd 7217) * $signed(input_fmap_20[15:0]) +
	( 14'sd 4893) * $signed(input_fmap_21[15:0]) +
	( 16'sd 31930) * $signed(input_fmap_22[15:0]) +
	( 16'sd 25360) * $signed(input_fmap_23[15:0]) +
	( 15'sd 11841) * $signed(input_fmap_24[15:0]) +
	( 11'sd 571) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22456) * $signed(input_fmap_26[15:0]) +
	( 14'sd 5880) * $signed(input_fmap_27[15:0]) +
	( 15'sd 15628) * $signed(input_fmap_28[15:0]) +
	( 15'sd 11258) * $signed(input_fmap_29[15:0]) +
	( 15'sd 16192) * $signed(input_fmap_30[15:0]) +
	( 16'sd 30586) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28073) * $signed(input_fmap_32[15:0]) +
	( 11'sd 694) * $signed(input_fmap_33[15:0]) +
	( 16'sd 24835) * $signed(input_fmap_34[15:0]) +
	( 16'sd 21630) * $signed(input_fmap_35[15:0]) +
	( 14'sd 5115) * $signed(input_fmap_36[15:0]) +
	( 14'sd 4594) * $signed(input_fmap_37[15:0]) +
	( 16'sd 32361) * $signed(input_fmap_38[15:0]) +
	( 16'sd 18133) * $signed(input_fmap_39[15:0]) +
	( 16'sd 21927) * $signed(input_fmap_40[15:0]) +
	( 16'sd 25741) * $signed(input_fmap_41[15:0]) +
	( 16'sd 31724) * $signed(input_fmap_42[15:0]) +
	( 16'sd 25635) * $signed(input_fmap_43[15:0]) +
	( 16'sd 32365) * $signed(input_fmap_44[15:0]) +
	( 15'sd 13193) * $signed(input_fmap_45[15:0]) +
	( 16'sd 22961) * $signed(input_fmap_46[15:0]) +
	( 15'sd 8913) * $signed(input_fmap_47[15:0]) +
	( 14'sd 7067) * $signed(input_fmap_48[15:0]) +
	( 16'sd 16668) * $signed(input_fmap_49[15:0]) +
	( 16'sd 30188) * $signed(input_fmap_50[15:0]) +
	( 15'sd 10262) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3082) * $signed(input_fmap_52[15:0]) +
	( 15'sd 13828) * $signed(input_fmap_53[15:0]) +
	( 14'sd 6792) * $signed(input_fmap_54[15:0]) +
	( 14'sd 5920) * $signed(input_fmap_55[15:0]) +
	( 16'sd 21951) * $signed(input_fmap_56[15:0]) +
	( 16'sd 31502) * $signed(input_fmap_57[15:0]) +
	( 16'sd 21284) * $signed(input_fmap_58[15:0]) +
	( 16'sd 20099) * $signed(input_fmap_59[15:0]) +
	( 16'sd 30755) * $signed(input_fmap_60[15:0]) +
	( 15'sd 12115) * $signed(input_fmap_61[15:0]) +
	( 16'sd 20979) * $signed(input_fmap_62[15:0]) +
	( 14'sd 5595) * $signed(input_fmap_63[15:0]) +
	( 16'sd 22922) * $signed(input_fmap_64[15:0]) +
	( 16'sd 22064) * $signed(input_fmap_65[15:0]) +
	( 16'sd 20332) * $signed(input_fmap_66[15:0]) +
	( 13'sd 2614) * $signed(input_fmap_67[15:0]) +
	( 15'sd 10455) * $signed(input_fmap_68[15:0]) +
	( 15'sd 15987) * $signed(input_fmap_69[15:0]) +
	( 15'sd 14665) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31711) * $signed(input_fmap_71[15:0]) +
	( 14'sd 6906) * $signed(input_fmap_72[15:0]) +
	( 11'sd 888) * $signed(input_fmap_73[15:0]) +
	( 16'sd 21640) * $signed(input_fmap_74[15:0]) +
	( 16'sd 22395) * $signed(input_fmap_75[15:0]) +
	( 16'sd 28976) * $signed(input_fmap_76[15:0]) +
	( 14'sd 5552) * $signed(input_fmap_77[15:0]) +
	( 14'sd 6636) * $signed(input_fmap_78[15:0]) +
	( 14'sd 7251) * $signed(input_fmap_79[15:0]) +
	( 14'sd 6613) * $signed(input_fmap_80[15:0]) +
	( 16'sd 30850) * $signed(input_fmap_81[15:0]) +
	( 12'sd 1582) * $signed(input_fmap_82[15:0]) +
	( 16'sd 21890) * $signed(input_fmap_83[15:0]) +
	( 10'sd 472) * $signed(input_fmap_84[15:0]) +
	( 16'sd 19703) * $signed(input_fmap_85[15:0]) +
	( 15'sd 8467) * $signed(input_fmap_86[15:0]) +
	( 16'sd 28878) * $signed(input_fmap_87[15:0]) +
	( 16'sd 26265) * $signed(input_fmap_88[15:0]) +
	( 13'sd 3533) * $signed(input_fmap_89[15:0]) +
	( 15'sd 14165) * $signed(input_fmap_90[15:0]) +
	( 15'sd 12011) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25705) * $signed(input_fmap_92[15:0]) +
	( 15'sd 12729) * $signed(input_fmap_93[15:0]) +
	( 15'sd 10615) * $signed(input_fmap_94[15:0]) +
	( 14'sd 7533) * $signed(input_fmap_95[15:0]) +
	( 15'sd 10768) * $signed(input_fmap_96[15:0]) +
	( 16'sd 19605) * $signed(input_fmap_97[15:0]) +
	( 13'sd 4047) * $signed(input_fmap_98[15:0]) +
	( 16'sd 31102) * $signed(input_fmap_99[15:0]) +
	( 16'sd 32600) * $signed(input_fmap_100[15:0]) +
	( 16'sd 25413) * $signed(input_fmap_101[15:0]) +
	( 16'sd 26016) * $signed(input_fmap_102[15:0]) +
	( 11'sd 663) * $signed(input_fmap_103[15:0]) +
	( 16'sd 17956) * $signed(input_fmap_104[15:0]) +
	( 15'sd 15004) * $signed(input_fmap_105[15:0]) +
	( 15'sd 11199) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27179) * $signed(input_fmap_107[15:0]) +
	( 16'sd 17003) * $signed(input_fmap_108[15:0]) +
	( 16'sd 31758) * $signed(input_fmap_109[15:0]) +
	( 14'sd 7688) * $signed(input_fmap_110[15:0]) +
	( 16'sd 19230) * $signed(input_fmap_111[15:0]) +
	( 15'sd 8980) * $signed(input_fmap_112[15:0]) +
	( 11'sd 884) * $signed(input_fmap_113[15:0]) +
	( 16'sd 29345) * $signed(input_fmap_114[15:0]) +
	( 16'sd 20490) * $signed(input_fmap_115[15:0]) +
	( 16'sd 24961) * $signed(input_fmap_116[15:0]) +
	( 15'sd 8280) * $signed(input_fmap_117[15:0]) +
	( 16'sd 30387) * $signed(input_fmap_118[15:0]) +
	( 16'sd 22073) * $signed(input_fmap_119[15:0]) +
	( 16'sd 18295) * $signed(input_fmap_120[15:0]) +
	( 15'sd 14295) * $signed(input_fmap_121[15:0]) +
	( 15'sd 15513) * $signed(input_fmap_122[15:0]) +
	( 16'sd 28956) * $signed(input_fmap_123[15:0]) +
	( 16'sd 29101) * $signed(input_fmap_124[15:0]) +
	( 15'sd 8760) * $signed(input_fmap_125[15:0]) +
	( 16'sd 27342) * $signed(input_fmap_126[15:0]) +
	( 13'sd 2071) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 16'sd 20422) * $signed(input_fmap_0[15:0]) +
	( 16'sd 22851) * $signed(input_fmap_1[15:0]) +
	( 16'sd 26742) * $signed(input_fmap_2[15:0]) +
	( 16'sd 26875) * $signed(input_fmap_3[15:0]) +
	( 15'sd 11062) * $signed(input_fmap_4[15:0]) +
	( 16'sd 26356) * $signed(input_fmap_5[15:0]) +
	( 16'sd 22589) * $signed(input_fmap_6[15:0]) +
	( 16'sd 21113) * $signed(input_fmap_7[15:0]) +
	( 14'sd 7261) * $signed(input_fmap_8[15:0]) +
	( 16'sd 30959) * $signed(input_fmap_9[15:0]) +
	( 16'sd 25368) * $signed(input_fmap_10[15:0]) +
	( 16'sd 18111) * $signed(input_fmap_11[15:0]) +
	( 15'sd 14719) * $signed(input_fmap_12[15:0]) +
	( 15'sd 9156) * $signed(input_fmap_13[15:0]) +
	( 16'sd 26459) * $signed(input_fmap_14[15:0]) +
	( 16'sd 23340) * $signed(input_fmap_15[15:0]) +
	( 14'sd 8008) * $signed(input_fmap_16[15:0]) +
	( 16'sd 26637) * $signed(input_fmap_17[15:0]) +
	( 16'sd 17860) * $signed(input_fmap_18[15:0]) +
	( 14'sd 5809) * $signed(input_fmap_19[15:0]) +
	( 16'sd 31462) * $signed(input_fmap_20[15:0]) +
	( 15'sd 8928) * $signed(input_fmap_21[15:0]) +
	( 15'sd 14601) * $signed(input_fmap_22[15:0]) +
	( 16'sd 26068) * $signed(input_fmap_23[15:0]) +
	( 16'sd 32212) * $signed(input_fmap_24[15:0]) +
	( 15'sd 10578) * $signed(input_fmap_25[15:0]) +
	( 13'sd 2889) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2455) * $signed(input_fmap_27[15:0]) +
	( 16'sd 27573) * $signed(input_fmap_28[15:0]) +
	( 16'sd 27640) * $signed(input_fmap_29[15:0]) +
	( 14'sd 7400) * $signed(input_fmap_30[15:0]) +
	( 14'sd 6948) * $signed(input_fmap_31[15:0]) +
	( 16'sd 28548) * $signed(input_fmap_32[15:0]) +
	( 15'sd 12685) * $signed(input_fmap_33[15:0]) +
	( 16'sd 24060) * $signed(input_fmap_34[15:0]) +
	( 13'sd 2748) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11035) * $signed(input_fmap_36[15:0]) +
	( 16'sd 29536) * $signed(input_fmap_37[15:0]) +
	( 15'sd 11806) * $signed(input_fmap_38[15:0]) +
	( 16'sd 21837) * $signed(input_fmap_39[15:0]) +
	( 14'sd 4813) * $signed(input_fmap_40[15:0]) +
	( 16'sd 26530) * $signed(input_fmap_41[15:0]) +
	( 16'sd 22612) * $signed(input_fmap_42[15:0]) +
	( 16'sd 25292) * $signed(input_fmap_43[15:0]) +
	( 15'sd 8259) * $signed(input_fmap_44[15:0]) +
	( 15'sd 14173) * $signed(input_fmap_45[15:0]) +
	( 16'sd 27671) * $signed(input_fmap_46[15:0]) +
	( 15'sd 8863) * $signed(input_fmap_47[15:0]) +
	( 14'sd 4928) * $signed(input_fmap_48[15:0]) +
	( 16'sd 29324) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26277) * $signed(input_fmap_50[15:0]) +
	( 14'sd 6764) * $signed(input_fmap_51[15:0]) +
	( 16'sd 26085) * $signed(input_fmap_52[15:0]) +
	( 16'sd 17090) * $signed(input_fmap_53[15:0]) +
	( 16'sd 17828) * $signed(input_fmap_54[15:0]) +
	( 15'sd 14404) * $signed(input_fmap_55[15:0]) +
	( 16'sd 29982) * $signed(input_fmap_56[15:0]) +
	( 14'sd 5966) * $signed(input_fmap_57[15:0]) +
	( 16'sd 31422) * $signed(input_fmap_58[15:0]) +
	( 16'sd 31760) * $signed(input_fmap_59[15:0]) +
	( 15'sd 15995) * $signed(input_fmap_60[15:0]) +
	( 16'sd 22623) * $signed(input_fmap_61[15:0]) +
	( 15'sd 9927) * $signed(input_fmap_62[15:0]) +
	( 14'sd 7050) * $signed(input_fmap_63[15:0]) +
	( 16'sd 21467) * $signed(input_fmap_64[15:0]) +
	( 15'sd 13274) * $signed(input_fmap_65[15:0]) +
	( 11'sd 784) * $signed(input_fmap_66[15:0]) +
	( 16'sd 19378) * $signed(input_fmap_67[15:0]) +
	( 16'sd 30469) * $signed(input_fmap_68[15:0]) +
	( 14'sd 6686) * $signed(input_fmap_69[15:0]) +
	( 16'sd 16544) * $signed(input_fmap_70[15:0]) +
	( 16'sd 29407) * $signed(input_fmap_71[15:0]) +
	( 16'sd 20886) * $signed(input_fmap_72[15:0]) +
	( 16'sd 17969) * $signed(input_fmap_73[15:0]) +
	( 14'sd 7221) * $signed(input_fmap_74[15:0]) +
	( 16'sd 30812) * $signed(input_fmap_75[15:0]) +
	( 16'sd 25936) * $signed(input_fmap_76[15:0]) +
	( 16'sd 20352) * $signed(input_fmap_77[15:0]) +
	( 12'sd 1908) * $signed(input_fmap_78[15:0]) +
	( 15'sd 15623) * $signed(input_fmap_79[15:0]) +
	( 13'sd 2705) * $signed(input_fmap_80[15:0]) +
	( 16'sd 18587) * $signed(input_fmap_81[15:0]) +
	( 16'sd 31589) * $signed(input_fmap_82[15:0]) +
	( 14'sd 5840) * $signed(input_fmap_83[15:0]) +
	( 15'sd 10980) * $signed(input_fmap_84[15:0]) +
	( 16'sd 20771) * $signed(input_fmap_85[15:0]) +
	( 16'sd 21004) * $signed(input_fmap_86[15:0]) +
	( 14'sd 7326) * $signed(input_fmap_87[15:0]) +
	( 14'sd 5993) * $signed(input_fmap_88[15:0]) +
	( 15'sd 13314) * $signed(input_fmap_89[15:0]) +
	( 16'sd 28245) * $signed(input_fmap_90[15:0]) +
	( 16'sd 18567) * $signed(input_fmap_91[15:0]) +
	( 13'sd 2659) * $signed(input_fmap_92[15:0]) +
	( 13'sd 2666) * $signed(input_fmap_93[15:0]) +
	( 16'sd 21334) * $signed(input_fmap_94[15:0]) +
	( 16'sd 31376) * $signed(input_fmap_95[15:0]) +
	( 16'sd 27201) * $signed(input_fmap_96[15:0]) +
	( 16'sd 17725) * $signed(input_fmap_97[15:0]) +
	( 16'sd 30279) * $signed(input_fmap_98[15:0]) +
	( 16'sd 32193) * $signed(input_fmap_99[15:0]) +
	( 14'sd 5089) * $signed(input_fmap_100[15:0]) +
	( 16'sd 28372) * $signed(input_fmap_101[15:0]) +
	( 14'sd 5921) * $signed(input_fmap_102[15:0]) +
	( 12'sd 1929) * $signed(input_fmap_103[15:0]) +
	( 16'sd 19894) * $signed(input_fmap_104[15:0]) +
	( 16'sd 28932) * $signed(input_fmap_105[15:0]) +
	( 12'sd 1667) * $signed(input_fmap_106[15:0]) +
	( 16'sd 26600) * $signed(input_fmap_107[15:0]) +
	( 16'sd 19389) * $signed(input_fmap_108[15:0]) +
	( 16'sd 20682) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22422) * $signed(input_fmap_110[15:0]) +
	( 15'sd 13620) * $signed(input_fmap_111[15:0]) +
	( 15'sd 15269) * $signed(input_fmap_112[15:0]) +
	( 15'sd 16144) * $signed(input_fmap_113[15:0]) +
	( 13'sd 3062) * $signed(input_fmap_114[15:0]) +
	( 16'sd 26864) * $signed(input_fmap_115[15:0]) +
	( 12'sd 1214) * $signed(input_fmap_116[15:0]) +
	( 16'sd 28529) * $signed(input_fmap_117[15:0]) +
	( 15'sd 15324) * $signed(input_fmap_118[15:0]) +
	( 16'sd 31904) * $signed(input_fmap_119[15:0]) +
	( 15'sd 11097) * $signed(input_fmap_120[15:0]) +
	( 13'sd 2527) * $signed(input_fmap_121[15:0]) +
	( 16'sd 30564) * $signed(input_fmap_122[15:0]) +
	( 16'sd 17488) * $signed(input_fmap_123[15:0]) +
	( 16'sd 22645) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24277) * $signed(input_fmap_125[15:0]) +
	( 15'sd 12109) * $signed(input_fmap_126[15:0]) +
	( 16'sd 29795) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 16'sd 27336) * $signed(input_fmap_0[15:0]) +
	( 12'sd 1316) * $signed(input_fmap_1[15:0]) +
	( 15'sd 11684) * $signed(input_fmap_2[15:0]) +
	( 15'sd 10773) * $signed(input_fmap_3[15:0]) +
	( 16'sd 31784) * $signed(input_fmap_4[15:0]) +
	( 16'sd 29053) * $signed(input_fmap_5[15:0]) +
	( 16'sd 26342) * $signed(input_fmap_6[15:0]) +
	( 16'sd 19941) * $signed(input_fmap_7[15:0]) +
	( 16'sd 27808) * $signed(input_fmap_8[15:0]) +
	( 14'sd 5395) * $signed(input_fmap_9[15:0]) +
	( 16'sd 22125) * $signed(input_fmap_10[15:0]) +
	( 16'sd 26131) * $signed(input_fmap_11[15:0]) +
	( 15'sd 11117) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24968) * $signed(input_fmap_13[15:0]) +
	( 16'sd 29093) * $signed(input_fmap_14[15:0]) +
	( 15'sd 8917) * $signed(input_fmap_15[15:0]) +
	( 16'sd 19497) * $signed(input_fmap_16[15:0]) +
	( 15'sd 11603) * $signed(input_fmap_17[15:0]) +
	( 11'sd 916) * $signed(input_fmap_18[15:0]) +
	( 16'sd 23347) * $signed(input_fmap_19[15:0]) +
	( 16'sd 19762) * $signed(input_fmap_20[15:0]) +
	( 16'sd 30017) * $signed(input_fmap_21[15:0]) +
	( 15'sd 10466) * $signed(input_fmap_22[15:0]) +
	( 14'sd 5294) * $signed(input_fmap_23[15:0]) +
	( 16'sd 24556) * $signed(input_fmap_24[15:0]) +
	( 12'sd 1209) * $signed(input_fmap_25[15:0]) +
	( 16'sd 25191) * $signed(input_fmap_26[15:0]) +
	( 16'sd 29750) * $signed(input_fmap_27[15:0]) +
	( 14'sd 7154) * $signed(input_fmap_28[15:0]) +
	( 16'sd 29106) * $signed(input_fmap_29[15:0]) +
	( 16'sd 26487) * $signed(input_fmap_30[15:0]) +
	( 16'sd 20296) * $signed(input_fmap_31[15:0]) +
	( 14'sd 6405) * $signed(input_fmap_32[15:0]) +
	( 16'sd 26408) * $signed(input_fmap_33[15:0]) +
	( 16'sd 29884) * $signed(input_fmap_34[15:0]) +
	( 13'sd 3572) * $signed(input_fmap_35[15:0]) +
	( 16'sd 30886) * $signed(input_fmap_36[15:0]) +
	( 15'sd 15548) * $signed(input_fmap_37[15:0]) +
	( 16'sd 29792) * $signed(input_fmap_38[15:0]) +
	( 16'sd 21708) * $signed(input_fmap_39[15:0]) +
	( 14'sd 4565) * $signed(input_fmap_40[15:0]) +
	( 14'sd 5471) * $signed(input_fmap_41[15:0]) +
	( 15'sd 8990) * $signed(input_fmap_42[15:0]) +
	( 16'sd 27160) * $signed(input_fmap_43[15:0]) +
	( 13'sd 2365) * $signed(input_fmap_44[15:0]) +
	( 15'sd 11899) * $signed(input_fmap_45[15:0]) +
	( 15'sd 15998) * $signed(input_fmap_46[15:0]) +
	( 16'sd 32010) * $signed(input_fmap_47[15:0]) +
	( 14'sd 4511) * $signed(input_fmap_48[15:0]) +
	( 15'sd 11330) * $signed(input_fmap_49[15:0]) +
	( 16'sd 30123) * $signed(input_fmap_50[15:0]) +
	( 15'sd 9719) * $signed(input_fmap_51[15:0]) +
	( 14'sd 7904) * $signed(input_fmap_52[15:0]) +
	( 15'sd 13240) * $signed(input_fmap_53[15:0]) +
	( 15'sd 12039) * $signed(input_fmap_54[15:0]) +
	( 15'sd 8682) * $signed(input_fmap_55[15:0]) +
	( 16'sd 27203) * $signed(input_fmap_56[15:0]) +
	( 15'sd 16045) * $signed(input_fmap_57[15:0]) +
	( 16'sd 25618) * $signed(input_fmap_58[15:0]) +
	( 15'sd 15740) * $signed(input_fmap_59[15:0]) +
	( 16'sd 22984) * $signed(input_fmap_60[15:0]) +
	( 12'sd 1854) * $signed(input_fmap_61[15:0]) +
	( 16'sd 24763) * $signed(input_fmap_62[15:0]) +
	( 16'sd 18999) * $signed(input_fmap_63[15:0]) +
	( 16'sd 30910) * $signed(input_fmap_64[15:0]) +
	( 13'sd 3794) * $signed(input_fmap_65[15:0]) +
	( 15'sd 11370) * $signed(input_fmap_66[15:0]) +
	( 16'sd 29302) * $signed(input_fmap_67[15:0]) +
	( 16'sd 29586) * $signed(input_fmap_68[15:0]) +
	( 14'sd 4649) * $signed(input_fmap_69[15:0]) +
	( 16'sd 30982) * $signed(input_fmap_70[15:0]) +
	( 16'sd 26226) * $signed(input_fmap_71[15:0]) +
	( 16'sd 26280) * $signed(input_fmap_72[15:0]) +
	( 15'sd 13615) * $signed(input_fmap_73[15:0]) +
	( 10'sd 324) * $signed(input_fmap_74[15:0]) +
	( 16'sd 26326) * $signed(input_fmap_75[15:0]) +
	( 9'sd 129) * $signed(input_fmap_76[15:0]) +
	( 16'sd 32680) * $signed(input_fmap_77[15:0]) +
	( 16'sd 18829) * $signed(input_fmap_78[15:0]) +
	( 12'sd 1751) * $signed(input_fmap_79[15:0]) +
	( 14'sd 5051) * $signed(input_fmap_80[15:0]) +
	( 16'sd 25994) * $signed(input_fmap_81[15:0]) +
	( 16'sd 23910) * $signed(input_fmap_82[15:0]) +
	( 16'sd 22585) * $signed(input_fmap_83[15:0]) +
	( 15'sd 10683) * $signed(input_fmap_84[15:0]) +
	( 16'sd 28821) * $signed(input_fmap_85[15:0]) +
	( 15'sd 14844) * $signed(input_fmap_86[15:0]) +
	( 14'sd 7670) * $signed(input_fmap_87[15:0]) +
	( 16'sd 32712) * $signed(input_fmap_88[15:0]) +
	( 15'sd 15912) * $signed(input_fmap_89[15:0]) +
	( 16'sd 22604) * $signed(input_fmap_90[15:0]) +
	( 16'sd 25600) * $signed(input_fmap_91[15:0]) +
	( 16'sd 19433) * $signed(input_fmap_92[15:0]) +
	( 14'sd 6809) * $signed(input_fmap_93[15:0]) +
	( 16'sd 23024) * $signed(input_fmap_94[15:0]) +
	( 14'sd 5672) * $signed(input_fmap_95[15:0]) +
	( 15'sd 8910) * $signed(input_fmap_96[15:0]) +
	( 15'sd 13123) * $signed(input_fmap_97[15:0]) +
	( 16'sd 20911) * $signed(input_fmap_98[15:0]) +
	( 16'sd 16863) * $signed(input_fmap_99[15:0]) +
	( 13'sd 2275) * $signed(input_fmap_100[15:0]) +
	( 16'sd 19838) * $signed(input_fmap_101[15:0]) +
	( 16'sd 22625) * $signed(input_fmap_102[15:0]) +
	( 16'sd 30562) * $signed(input_fmap_103[15:0]) +
	( 16'sd 19129) * $signed(input_fmap_104[15:0]) +
	( 12'sd 1899) * $signed(input_fmap_105[15:0]) +
	( 15'sd 11927) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27844) * $signed(input_fmap_107[15:0]) +
	( 14'sd 5103) * $signed(input_fmap_108[15:0]) +
	( 13'sd 3657) * $signed(input_fmap_109[15:0]) +
	( 16'sd 30013) * $signed(input_fmap_110[15:0]) +
	( 16'sd 26015) * $signed(input_fmap_111[15:0]) +
	( 15'sd 11825) * $signed(input_fmap_112[15:0]) +
	( 15'sd 12311) * $signed(input_fmap_113[15:0]) +
	( 16'sd 25518) * $signed(input_fmap_114[15:0]) +
	( 16'sd 31839) * $signed(input_fmap_115[15:0]) +
	( 14'sd 4931) * $signed(input_fmap_116[15:0]) +
	( 16'sd 32007) * $signed(input_fmap_117[15:0]) +
	( 16'sd 30037) * $signed(input_fmap_118[15:0]) +
	( 15'sd 10069) * $signed(input_fmap_119[15:0]) +
	( 16'sd 25918) * $signed(input_fmap_120[15:0]) +
	( 16'sd 19529) * $signed(input_fmap_121[15:0]) +
	( 16'sd 31334) * $signed(input_fmap_122[15:0]) +
	( 16'sd 20879) * $signed(input_fmap_123[15:0]) +
	( 15'sd 12799) * $signed(input_fmap_124[15:0]) +
	( 16'sd 19755) * $signed(input_fmap_125[15:0]) +
	( 15'sd 15798) * $signed(input_fmap_126[15:0]) +
	( 16'sd 30215) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 15'sd 12527) * $signed(input_fmap_0[15:0]) +
	( 16'sd 17215) * $signed(input_fmap_1[15:0]) +
	( 15'sd 14248) * $signed(input_fmap_2[15:0]) +
	( 15'sd 14548) * $signed(input_fmap_3[15:0]) +
	( 15'sd 8279) * $signed(input_fmap_4[15:0]) +
	( 15'sd 13446) * $signed(input_fmap_5[15:0]) +
	( 15'sd 15230) * $signed(input_fmap_6[15:0]) +
	( 15'sd 8392) * $signed(input_fmap_7[15:0]) +
	( 16'sd 19669) * $signed(input_fmap_8[15:0]) +
	( 13'sd 2860) * $signed(input_fmap_9[15:0]) +
	( 16'sd 17770) * $signed(input_fmap_10[15:0]) +
	( 14'sd 4213) * $signed(input_fmap_11[15:0]) +
	( 16'sd 31084) * $signed(input_fmap_12[15:0]) +
	( 16'sd 19415) * $signed(input_fmap_13[15:0]) +
	( 16'sd 27208) * $signed(input_fmap_14[15:0]) +
	( 16'sd 17796) * $signed(input_fmap_15[15:0]) +
	( 15'sd 12756) * $signed(input_fmap_16[15:0]) +
	( 13'sd 2898) * $signed(input_fmap_17[15:0]) +
	( 16'sd 20021) * $signed(input_fmap_18[15:0]) +
	( 16'sd 26989) * $signed(input_fmap_19[15:0]) +
	( 16'sd 20185) * $signed(input_fmap_20[15:0]) +
	( 16'sd 31757) * $signed(input_fmap_21[15:0]) +
	( 14'sd 7252) * $signed(input_fmap_22[15:0]) +
	( 16'sd 19517) * $signed(input_fmap_23[15:0]) +
	( 15'sd 11818) * $signed(input_fmap_24[15:0]) +
	( 15'sd 15351) * $signed(input_fmap_25[15:0]) +
	( 16'sd 21141) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1749) * $signed(input_fmap_27[15:0]) +
	( 15'sd 14423) * $signed(input_fmap_28[15:0]) +
	( 16'sd 25031) * $signed(input_fmap_29[15:0]) +
	( 12'sd 1226) * $signed(input_fmap_30[15:0]) +
	( 16'sd 16447) * $signed(input_fmap_31[15:0]) +
	( 16'sd 20810) * $signed(input_fmap_32[15:0]) +
	( 14'sd 6266) * $signed(input_fmap_33[15:0]) +
	( 15'sd 16191) * $signed(input_fmap_34[15:0]) +
	( 16'sd 24906) * $signed(input_fmap_35[15:0]) +
	( 11'sd 746) * $signed(input_fmap_36[15:0]) +
	( 16'sd 28683) * $signed(input_fmap_37[15:0]) +
	( 16'sd 19112) * $signed(input_fmap_38[15:0]) +
	( 16'sd 18085) * $signed(input_fmap_39[15:0]) +
	( 16'sd 26509) * $signed(input_fmap_40[15:0]) +
	( 14'sd 6340) * $signed(input_fmap_41[15:0]) +
	( 15'sd 13070) * $signed(input_fmap_42[15:0]) +
	( 16'sd 24308) * $signed(input_fmap_43[15:0]) +
	( 11'sd 541) * $signed(input_fmap_44[15:0]) +
	( 15'sd 10428) * $signed(input_fmap_45[15:0]) +
	( 15'sd 10279) * $signed(input_fmap_46[15:0]) +
	( 16'sd 27197) * $signed(input_fmap_47[15:0]) +
	( 15'sd 10157) * $signed(input_fmap_48[15:0]) +
	( 15'sd 10648) * $signed(input_fmap_49[15:0]) +
	( 16'sd 18380) * $signed(input_fmap_50[15:0]) +
	( 16'sd 26108) * $signed(input_fmap_51[15:0]) +
	( 16'sd 16910) * $signed(input_fmap_52[15:0]) +
	( 15'sd 15118) * $signed(input_fmap_53[15:0]) +
	( 16'sd 21755) * $signed(input_fmap_54[15:0]) +
	( 16'sd 16432) * $signed(input_fmap_55[15:0]) +
	( 16'sd 16835) * $signed(input_fmap_56[15:0]) +
	( 14'sd 7249) * $signed(input_fmap_57[15:0]) +
	( 16'sd 16415) * $signed(input_fmap_58[15:0]) +
	( 15'sd 14411) * $signed(input_fmap_59[15:0]) +
	( 14'sd 5715) * $signed(input_fmap_60[15:0]) +
	( 16'sd 32609) * $signed(input_fmap_61[15:0]) +
	( 16'sd 32293) * $signed(input_fmap_62[15:0]) +
	( 16'sd 29956) * $signed(input_fmap_63[15:0]) +
	( 14'sd 4627) * $signed(input_fmap_64[15:0]) +
	( 15'sd 14325) * $signed(input_fmap_65[15:0]) +
	( 10'sd 424) * $signed(input_fmap_66[15:0]) +
	( 16'sd 26008) * $signed(input_fmap_67[15:0]) +
	( 14'sd 7385) * $signed(input_fmap_68[15:0]) +
	( 16'sd 17419) * $signed(input_fmap_69[15:0]) +
	( 13'sd 3215) * $signed(input_fmap_70[15:0]) +
	( 16'sd 21557) * $signed(input_fmap_71[15:0]) +
	( 16'sd 19539) * $signed(input_fmap_72[15:0]) +
	( 16'sd 26458) * $signed(input_fmap_73[15:0]) +
	( 16'sd 24381) * $signed(input_fmap_74[15:0]) +
	( 16'sd 21469) * $signed(input_fmap_75[15:0]) +
	( 16'sd 27154) * $signed(input_fmap_76[15:0]) +
	( 13'sd 2767) * $signed(input_fmap_77[15:0]) +
	( 16'sd 26869) * $signed(input_fmap_78[15:0]) +
	( 16'sd 19126) * $signed(input_fmap_79[15:0]) +
	( 15'sd 14846) * $signed(input_fmap_80[15:0]) +
	( 13'sd 2894) * $signed(input_fmap_81[15:0]) +
	( 16'sd 17960) * $signed(input_fmap_82[15:0]) +
	( 15'sd 14771) * $signed(input_fmap_83[15:0]) +
	( 16'sd 28811) * $signed(input_fmap_84[15:0]) +
	( 15'sd 10379) * $signed(input_fmap_85[15:0]) +
	( 9'sd 188) * $signed(input_fmap_86[15:0]) +
	( 16'sd 27073) * $signed(input_fmap_87[15:0]) +
	( 16'sd 27296) * $signed(input_fmap_88[15:0]) +
	( 11'sd 881) * $signed(input_fmap_89[15:0]) +
	( 16'sd 17801) * $signed(input_fmap_90[15:0]) +
	( 12'sd 1061) * $signed(input_fmap_91[15:0]) +
	( 13'sd 2877) * $signed(input_fmap_92[15:0]) +
	( 15'sd 9348) * $signed(input_fmap_93[15:0]) +
	( 16'sd 32112) * $signed(input_fmap_94[15:0]) +
	( 14'sd 7532) * $signed(input_fmap_95[15:0]) +
	( 14'sd 5373) * $signed(input_fmap_96[15:0]) +
	( 16'sd 31117) * $signed(input_fmap_97[15:0]) +
	( 10'sd 327) * $signed(input_fmap_98[15:0]) +
	( 16'sd 25683) * $signed(input_fmap_99[15:0]) +
	( 11'sd 620) * $signed(input_fmap_100[15:0]) +
	( 14'sd 7489) * $signed(input_fmap_101[15:0]) +
	( 16'sd 29222) * $signed(input_fmap_102[15:0]) +
	( 16'sd 20330) * $signed(input_fmap_103[15:0]) +
	( 14'sd 4506) * $signed(input_fmap_104[15:0]) +
	( 16'sd 30166) * $signed(input_fmap_105[15:0]) +
	( 15'sd 15505) * $signed(input_fmap_106[15:0]) +
	( 15'sd 12597) * $signed(input_fmap_107[15:0]) +
	( 14'sd 4727) * $signed(input_fmap_108[15:0]) +
	( 16'sd 16952) * $signed(input_fmap_109[15:0]) +
	( 8'sd 126) * $signed(input_fmap_110[15:0]) +
	( 16'sd 26564) * $signed(input_fmap_111[15:0]) +
	( 16'sd 22545) * $signed(input_fmap_112[15:0]) +
	( 16'sd 17075) * $signed(input_fmap_113[15:0]) +
	( 15'sd 14788) * $signed(input_fmap_114[15:0]) +
	( 16'sd 31220) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26380) * $signed(input_fmap_116[15:0]) +
	( 16'sd 20499) * $signed(input_fmap_117[15:0]) +
	( 16'sd 20046) * $signed(input_fmap_118[15:0]) +
	( 9'sd 130) * $signed(input_fmap_119[15:0]) +
	( 14'sd 5170) * $signed(input_fmap_120[15:0]) +
	( 16'sd 24825) * $signed(input_fmap_121[15:0]) +
	( 16'sd 20484) * $signed(input_fmap_122[15:0]) +
	( 16'sd 18422) * $signed(input_fmap_123[15:0]) +
	( 12'sd 1823) * $signed(input_fmap_124[15:0]) +
	( 16'sd 17915) * $signed(input_fmap_125[15:0]) +
	( 14'sd 7910) * $signed(input_fmap_126[15:0]) +
	( 15'sd 16177) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 12'sd 1794) * $signed(input_fmap_0[15:0]) +
	( 13'sd 2178) * $signed(input_fmap_1[15:0]) +
	( 14'sd 5163) * $signed(input_fmap_2[15:0]) +
	( 16'sd 22750) * $signed(input_fmap_3[15:0]) +
	( 16'sd 28746) * $signed(input_fmap_4[15:0]) +
	( 13'sd 2710) * $signed(input_fmap_5[15:0]) +
	( 15'sd 10478) * $signed(input_fmap_6[15:0]) +
	( 16'sd 27349) * $signed(input_fmap_7[15:0]) +
	( 14'sd 6194) * $signed(input_fmap_8[15:0]) +
	( 16'sd 27722) * $signed(input_fmap_9[15:0]) +
	( 15'sd 8684) * $signed(input_fmap_10[15:0]) +
	( 13'sd 3038) * $signed(input_fmap_11[15:0]) +
	( 15'sd 14101) * $signed(input_fmap_12[15:0]) +
	( 15'sd 10412) * $signed(input_fmap_13[15:0]) +
	( 12'sd 1616) * $signed(input_fmap_14[15:0]) +
	( 15'sd 13472) * $signed(input_fmap_15[15:0]) +
	( 16'sd 20478) * $signed(input_fmap_16[15:0]) +
	( 13'sd 2655) * $signed(input_fmap_17[15:0]) +
	( 15'sd 12263) * $signed(input_fmap_18[15:0]) +
	( 16'sd 20131) * $signed(input_fmap_19[15:0]) +
	( 15'sd 15027) * $signed(input_fmap_20[15:0]) +
	( 15'sd 10814) * $signed(input_fmap_21[15:0]) +
	( 12'sd 1748) * $signed(input_fmap_22[15:0]) +
	( 16'sd 20427) * $signed(input_fmap_23[15:0]) +
	( 16'sd 25888) * $signed(input_fmap_24[15:0]) +
	( 16'sd 17924) * $signed(input_fmap_25[15:0]) +
	( 16'sd 21627) * $signed(input_fmap_26[15:0]) +
	( 14'sd 7841) * $signed(input_fmap_27[15:0]) +
	( 16'sd 29792) * $signed(input_fmap_28[15:0]) +
	( 14'sd 8006) * $signed(input_fmap_29[15:0]) +
	( 12'sd 1101) * $signed(input_fmap_30[15:0]) +
	( 16'sd 17946) * $signed(input_fmap_31[15:0]) +
	( 16'sd 25893) * $signed(input_fmap_32[15:0]) +
	( 16'sd 22042) * $signed(input_fmap_33[15:0]) +
	( 13'sd 3254) * $signed(input_fmap_34[15:0]) +
	( 16'sd 19771) * $signed(input_fmap_35[15:0]) +
	( 16'sd 19969) * $signed(input_fmap_36[15:0]) +
	( 12'sd 1879) * $signed(input_fmap_37[15:0]) +
	( 16'sd 28011) * $signed(input_fmap_38[15:0]) +
	( 15'sd 9889) * $signed(input_fmap_39[15:0]) +
	( 16'sd 21724) * $signed(input_fmap_40[15:0]) +
	( 16'sd 32035) * $signed(input_fmap_41[15:0]) +
	( 15'sd 12114) * $signed(input_fmap_42[15:0]) +
	( 16'sd 29667) * $signed(input_fmap_43[15:0]) +
	( 15'sd 12142) * $signed(input_fmap_44[15:0]) +
	( 16'sd 16593) * $signed(input_fmap_45[15:0]) +
	( 16'sd 23220) * $signed(input_fmap_46[15:0]) +
	( 16'sd 17021) * $signed(input_fmap_47[15:0]) +
	( 16'sd 17911) * $signed(input_fmap_48[15:0]) +
	( 15'sd 15671) * $signed(input_fmap_49[15:0]) +
	( 13'sd 2916) * $signed(input_fmap_50[15:0]) +
	( 14'sd 7105) * $signed(input_fmap_51[15:0]) +
	( 11'sd 755) * $signed(input_fmap_52[15:0]) +
	( 16'sd 27850) * $signed(input_fmap_53[15:0]) +
	( 16'sd 26896) * $signed(input_fmap_54[15:0]) +
	( 13'sd 2328) * $signed(input_fmap_55[15:0]) +
	( 16'sd 27066) * $signed(input_fmap_56[15:0]) +
	( 15'sd 10133) * $signed(input_fmap_57[15:0]) +
	( 15'sd 14457) * $signed(input_fmap_58[15:0]) +
	( 16'sd 19176) * $signed(input_fmap_59[15:0]) +
	( 15'sd 15301) * $signed(input_fmap_60[15:0]) +
	( 16'sd 18147) * $signed(input_fmap_61[15:0]) +
	( 16'sd 17789) * $signed(input_fmap_62[15:0]) +
	( 15'sd 11840) * $signed(input_fmap_63[15:0]) +
	( 13'sd 3410) * $signed(input_fmap_64[15:0]) +
	( 14'sd 6773) * $signed(input_fmap_65[15:0]) +
	( 12'sd 1403) * $signed(input_fmap_66[15:0]) +
	( 16'sd 24556) * $signed(input_fmap_67[15:0]) +
	( 16'sd 23940) * $signed(input_fmap_68[15:0]) +
	( 16'sd 29174) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31309) * $signed(input_fmap_70[15:0]) +
	( 14'sd 7058) * $signed(input_fmap_71[15:0]) +
	( 10'sd 328) * $signed(input_fmap_72[15:0]) +
	( 15'sd 14942) * $signed(input_fmap_73[15:0]) +
	( 12'sd 1698) * $signed(input_fmap_74[15:0]) +
	( 10'sd 270) * $signed(input_fmap_75[15:0]) +
	( 16'sd 21336) * $signed(input_fmap_76[15:0]) +
	( 15'sd 8946) * $signed(input_fmap_77[15:0]) +
	( 16'sd 17852) * $signed(input_fmap_78[15:0]) +
	( 14'sd 7592) * $signed(input_fmap_79[15:0]) +
	( 15'sd 13003) * $signed(input_fmap_80[15:0]) +
	( 15'sd 13588) * $signed(input_fmap_81[15:0]) +
	( 16'sd 25608) * $signed(input_fmap_82[15:0]) +
	( 14'sd 4540) * $signed(input_fmap_83[15:0]) +
	( 15'sd 12534) * $signed(input_fmap_84[15:0]) +
	( 15'sd 10344) * $signed(input_fmap_85[15:0]) +
	( 16'sd 27959) * $signed(input_fmap_86[15:0]) +
	( 16'sd 17767) * $signed(input_fmap_87[15:0]) +
	( 16'sd 25504) * $signed(input_fmap_88[15:0]) +
	( 15'sd 14835) * $signed(input_fmap_89[15:0]) +
	( 16'sd 23626) * $signed(input_fmap_90[15:0]) +
	( 16'sd 27044) * $signed(input_fmap_91[15:0]) +
	( 16'sd 20251) * $signed(input_fmap_92[15:0]) +
	( 14'sd 5509) * $signed(input_fmap_93[15:0]) +
	( 15'sd 9944) * $signed(input_fmap_94[15:0]) +
	( 16'sd 21306) * $signed(input_fmap_95[15:0]) +
	( 7'sd 57) * $signed(input_fmap_96[15:0]) +
	( 16'sd 17269) * $signed(input_fmap_97[15:0]) +
	( 13'sd 4093) * $signed(input_fmap_98[15:0]) +
	( 14'sd 6247) * $signed(input_fmap_99[15:0]) +
	( 16'sd 31118) * $signed(input_fmap_100[15:0]) +
	( 16'sd 30150) * $signed(input_fmap_101[15:0]) +
	( 16'sd 25009) * $signed(input_fmap_102[15:0]) +
	( 16'sd 26337) * $signed(input_fmap_103[15:0]) +
	( 16'sd 22093) * $signed(input_fmap_104[15:0]) +
	( 16'sd 22024) * $signed(input_fmap_105[15:0]) +
	( 16'sd 27243) * $signed(input_fmap_106[15:0]) +
	( 16'sd 28432) * $signed(input_fmap_107[15:0]) +
	( 16'sd 18654) * $signed(input_fmap_108[15:0]) +
	( 16'sd 26870) * $signed(input_fmap_109[15:0]) +
	( 14'sd 7541) * $signed(input_fmap_110[15:0]) +
	( 16'sd 25995) * $signed(input_fmap_111[15:0]) +
	( 16'sd 18926) * $signed(input_fmap_112[15:0]) +
	( 13'sd 3215) * $signed(input_fmap_113[15:0]) +
	( 15'sd 14134) * $signed(input_fmap_114[15:0]) +
	( 15'sd 12934) * $signed(input_fmap_115[15:0]) +
	( 16'sd 21142) * $signed(input_fmap_116[15:0]) +
	( 16'sd 16412) * $signed(input_fmap_117[15:0]) +
	( 14'sd 8088) * $signed(input_fmap_118[15:0]) +
	( 16'sd 21724) * $signed(input_fmap_119[15:0]) +
	( 16'sd 20699) * $signed(input_fmap_120[15:0]) +
	( 15'sd 11803) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9555) * $signed(input_fmap_122[15:0]) +
	( 13'sd 3938) * $signed(input_fmap_123[15:0]) +
	( 14'sd 5537) * $signed(input_fmap_124[15:0]) +
	( 16'sd 27499) * $signed(input_fmap_125[15:0]) +
	( 13'sd 2280) * $signed(input_fmap_126[15:0]) +
	( 15'sd 14487) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 16'sd 29927) * $signed(input_fmap_0[15:0]) +
	( 16'sd 19800) * $signed(input_fmap_1[15:0]) +
	( 16'sd 18860) * $signed(input_fmap_2[15:0]) +
	( 16'sd 19985) * $signed(input_fmap_3[15:0]) +
	( 14'sd 7582) * $signed(input_fmap_4[15:0]) +
	( 16'sd 23822) * $signed(input_fmap_5[15:0]) +
	( 13'sd 3358) * $signed(input_fmap_6[15:0]) +
	( 15'sd 15617) * $signed(input_fmap_7[15:0]) +
	( 15'sd 11487) * $signed(input_fmap_8[15:0]) +
	( 15'sd 12849) * $signed(input_fmap_9[15:0]) +
	( 16'sd 21305) * $signed(input_fmap_10[15:0]) +
	( 16'sd 28444) * $signed(input_fmap_11[15:0]) +
	( 15'sd 9961) * $signed(input_fmap_12[15:0]) +
	( 16'sd 19991) * $signed(input_fmap_13[15:0]) +
	( 15'sd 9296) * $signed(input_fmap_14[15:0]) +
	( 14'sd 7362) * $signed(input_fmap_15[15:0]) +
	( 14'sd 6669) * $signed(input_fmap_16[15:0]) +
	( 16'sd 20994) * $signed(input_fmap_17[15:0]) +
	( 16'sd 27569) * $signed(input_fmap_18[15:0]) +
	( 10'sd 411) * $signed(input_fmap_19[15:0]) +
	( 16'sd 23175) * $signed(input_fmap_20[15:0]) +
	( 16'sd 23994) * $signed(input_fmap_21[15:0]) +
	( 16'sd 24000) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24584) * $signed(input_fmap_23[15:0]) +
	( 16'sd 31074) * $signed(input_fmap_24[15:0]) +
	( 16'sd 32506) * $signed(input_fmap_25[15:0]) +
	( 16'sd 28889) * $signed(input_fmap_26[15:0]) +
	( 11'sd 617) * $signed(input_fmap_27[15:0]) +
	( 14'sd 6112) * $signed(input_fmap_28[15:0]) +
	( 16'sd 17311) * $signed(input_fmap_29[15:0]) +
	( 15'sd 10825) * $signed(input_fmap_30[15:0]) +
	( 16'sd 17213) * $signed(input_fmap_31[15:0]) +
	( 12'sd 2016) * $signed(input_fmap_32[15:0]) +
	( 16'sd 31757) * $signed(input_fmap_33[15:0]) +
	( 16'sd 17863) * $signed(input_fmap_34[15:0]) +
	( 16'sd 17976) * $signed(input_fmap_35[15:0]) +
	( 16'sd 25005) * $signed(input_fmap_36[15:0]) +
	( 16'sd 26292) * $signed(input_fmap_37[15:0]) +
	( 16'sd 29619) * $signed(input_fmap_38[15:0]) +
	( 14'sd 6693) * $signed(input_fmap_39[15:0]) +
	( 16'sd 22450) * $signed(input_fmap_40[15:0]) +
	( 13'sd 3589) * $signed(input_fmap_41[15:0]) +
	( 16'sd 23430) * $signed(input_fmap_42[15:0]) +
	( 14'sd 4932) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31091) * $signed(input_fmap_44[15:0]) +
	( 16'sd 26679) * $signed(input_fmap_45[15:0]) +
	( 16'sd 32488) * $signed(input_fmap_46[15:0]) +
	( 16'sd 29231) * $signed(input_fmap_47[15:0]) +
	( 14'sd 6237) * $signed(input_fmap_48[15:0]) +
	( 15'sd 11086) * $signed(input_fmap_49[15:0]) +
	( 14'sd 7734) * $signed(input_fmap_50[15:0]) +
	( 14'sd 5564) * $signed(input_fmap_51[15:0]) +
	( 15'sd 10687) * $signed(input_fmap_52[15:0]) +
	( 15'sd 15777) * $signed(input_fmap_53[15:0]) +
	( 16'sd 23841) * $signed(input_fmap_54[15:0]) +
	( 16'sd 27657) * $signed(input_fmap_55[15:0]) +
	( 9'sd 233) * $signed(input_fmap_56[15:0]) +
	( 15'sd 8984) * $signed(input_fmap_57[15:0]) +
	( 15'sd 14572) * $signed(input_fmap_58[15:0]) +
	( 16'sd 27280) * $signed(input_fmap_59[15:0]) +
	( 16'sd 27805) * $signed(input_fmap_60[15:0]) +
	( 14'sd 7023) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29129) * $signed(input_fmap_62[15:0]) +
	( 16'sd 29307) * $signed(input_fmap_63[15:0]) +
	( 16'sd 16754) * $signed(input_fmap_64[15:0]) +
	( 15'sd 14851) * $signed(input_fmap_65[15:0]) +
	( 13'sd 3841) * $signed(input_fmap_66[15:0]) +
	( 15'sd 13303) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26943) * $signed(input_fmap_68[15:0]) +
	( 16'sd 17807) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31268) * $signed(input_fmap_70[15:0]) +
	( 15'sd 12904) * $signed(input_fmap_71[15:0]) +
	( 13'sd 3762) * $signed(input_fmap_72[15:0]) +
	( 15'sd 12238) * $signed(input_fmap_73[15:0]) +
	( 16'sd 20916) * $signed(input_fmap_74[15:0]) +
	( 15'sd 8527) * $signed(input_fmap_75[15:0]) +
	( 16'sd 16854) * $signed(input_fmap_76[15:0]) +
	( 16'sd 30752) * $signed(input_fmap_77[15:0]) +
	( 15'sd 14378) * $signed(input_fmap_78[15:0]) +
	( 14'sd 7311) * $signed(input_fmap_79[15:0]) +
	( 15'sd 11093) * $signed(input_fmap_80[15:0]) +
	( 16'sd 23152) * $signed(input_fmap_81[15:0]) +
	( 15'sd 16240) * $signed(input_fmap_82[15:0]) +
	( 16'sd 19516) * $signed(input_fmap_83[15:0]) +
	( 16'sd 20792) * $signed(input_fmap_84[15:0]) +
	( 16'sd 21430) * $signed(input_fmap_85[15:0]) +
	( 13'sd 2782) * $signed(input_fmap_86[15:0]) +
	( 15'sd 12843) * $signed(input_fmap_87[15:0]) +
	( 13'sd 3961) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5221) * $signed(input_fmap_89[15:0]) +
	( 13'sd 2611) * $signed(input_fmap_90[15:0]) +
	( 16'sd 17934) * $signed(input_fmap_91[15:0]) +
	( 15'sd 12013) * $signed(input_fmap_92[15:0]) +
	( 15'sd 9295) * $signed(input_fmap_93[15:0]) +
	( 16'sd 31951) * $signed(input_fmap_94[15:0]) +
	( 16'sd 19900) * $signed(input_fmap_95[15:0]) +
	( 16'sd 30931) * $signed(input_fmap_96[15:0]) +
	( 14'sd 7117) * $signed(input_fmap_97[15:0]) +
	( 16'sd 21552) * $signed(input_fmap_98[15:0]) +
	( 15'sd 8393) * $signed(input_fmap_99[15:0]) +
	( 16'sd 16411) * $signed(input_fmap_100[15:0]) +
	( 16'sd 26620) * $signed(input_fmap_101[15:0]) +
	( 15'sd 8420) * $signed(input_fmap_102[15:0]) +
	( 16'sd 28588) * $signed(input_fmap_103[15:0]) +
	( 16'sd 29316) * $signed(input_fmap_104[15:0]) +
	( 16'sd 20309) * $signed(input_fmap_105[15:0]) +
	( 14'sd 4129) * $signed(input_fmap_106[15:0]) +
	( 16'sd 17333) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15881) * $signed(input_fmap_108[15:0]) +
	( 14'sd 4837) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22195) * $signed(input_fmap_110[15:0]) +
	( 15'sd 9948) * $signed(input_fmap_111[15:0]) +
	( 16'sd 19206) * $signed(input_fmap_112[15:0]) +
	( 15'sd 8724) * $signed(input_fmap_113[15:0]) +
	( 15'sd 8504) * $signed(input_fmap_114[15:0]) +
	( 15'sd 15777) * $signed(input_fmap_115[15:0]) +
	( 16'sd 23185) * $signed(input_fmap_116[15:0]) +
	( 16'sd 32120) * $signed(input_fmap_117[15:0]) +
	( 15'sd 8772) * $signed(input_fmap_118[15:0]) +
	( 16'sd 19661) * $signed(input_fmap_119[15:0]) +
	( 16'sd 28731) * $signed(input_fmap_120[15:0]) +
	( 15'sd 8299) * $signed(input_fmap_121[15:0]) +
	( 16'sd 28745) * $signed(input_fmap_122[15:0]) +
	( 16'sd 16690) * $signed(input_fmap_123[15:0]) +
	( 15'sd 10130) * $signed(input_fmap_124[15:0]) +
	( 13'sd 2243) * $signed(input_fmap_125[15:0]) +
	( 16'sd 28443) * $signed(input_fmap_126[15:0]) +
	( 16'sd 23330) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 16'sd 20618) * $signed(input_fmap_0[15:0]) +
	( 15'sd 9725) * $signed(input_fmap_1[15:0]) +
	( 8'sd 127) * $signed(input_fmap_2[15:0]) +
	( 13'sd 2720) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30995) * $signed(input_fmap_4[15:0]) +
	( 16'sd 19637) * $signed(input_fmap_5[15:0]) +
	( 15'sd 8657) * $signed(input_fmap_6[15:0]) +
	( 16'sd 28796) * $signed(input_fmap_7[15:0]) +
	( 16'sd 19989) * $signed(input_fmap_8[15:0]) +
	( 16'sd 30705) * $signed(input_fmap_9[15:0]) +
	( 16'sd 21942) * $signed(input_fmap_10[15:0]) +
	( 15'sd 11628) * $signed(input_fmap_11[15:0]) +
	( 13'sd 3207) * $signed(input_fmap_12[15:0]) +
	( 15'sd 11358) * $signed(input_fmap_13[15:0]) +
	( 16'sd 19744) * $signed(input_fmap_14[15:0]) +
	( 13'sd 2739) * $signed(input_fmap_15[15:0]) +
	( 16'sd 16979) * $signed(input_fmap_16[15:0]) +
	( 16'sd 28686) * $signed(input_fmap_17[15:0]) +
	( 14'sd 4993) * $signed(input_fmap_18[15:0]) +
	( 15'sd 13386) * $signed(input_fmap_19[15:0]) +
	( 13'sd 2361) * $signed(input_fmap_20[15:0]) +
	( 16'sd 18020) * $signed(input_fmap_21[15:0]) +
	( 14'sd 5301) * $signed(input_fmap_22[15:0]) +
	( 14'sd 5106) * $signed(input_fmap_23[15:0]) +
	( 15'sd 15432) * $signed(input_fmap_24[15:0]) +
	( 14'sd 6071) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22200) * $signed(input_fmap_26[15:0]) +
	( 13'sd 3177) * $signed(input_fmap_27[15:0]) +
	( 13'sd 3648) * $signed(input_fmap_28[15:0]) +
	( 15'sd 11859) * $signed(input_fmap_29[15:0]) +
	( 15'sd 13354) * $signed(input_fmap_30[15:0]) +
	( 16'sd 26401) * $signed(input_fmap_31[15:0]) +
	( 16'sd 22743) * $signed(input_fmap_32[15:0]) +
	( 16'sd 17153) * $signed(input_fmap_33[15:0]) +
	( 16'sd 17910) * $signed(input_fmap_34[15:0]) +
	( 16'sd 21990) * $signed(input_fmap_35[15:0]) +
	( 16'sd 27167) * $signed(input_fmap_36[15:0]) +
	( 16'sd 16932) * $signed(input_fmap_37[15:0]) +
	( 16'sd 19538) * $signed(input_fmap_38[15:0]) +
	( 16'sd 28907) * $signed(input_fmap_39[15:0]) +
	( 16'sd 21813) * $signed(input_fmap_40[15:0]) +
	( 15'sd 12327) * $signed(input_fmap_41[15:0]) +
	( 16'sd 21331) * $signed(input_fmap_42[15:0]) +
	( 16'sd 21342) * $signed(input_fmap_43[15:0]) +
	( 11'sd 794) * $signed(input_fmap_44[15:0]) +
	( 16'sd 23900) * $signed(input_fmap_45[15:0]) +
	( 14'sd 5624) * $signed(input_fmap_46[15:0]) +
	( 16'sd 31478) * $signed(input_fmap_47[15:0]) +
	( 14'sd 6035) * $signed(input_fmap_48[15:0]) +
	( 16'sd 30148) * $signed(input_fmap_49[15:0]) +
	( 16'sd 18584) * $signed(input_fmap_50[15:0]) +
	( 16'sd 31286) * $signed(input_fmap_51[15:0]) +
	( 15'sd 9622) * $signed(input_fmap_52[15:0]) +
	( 16'sd 32083) * $signed(input_fmap_53[15:0]) +
	( 16'sd 32738) * $signed(input_fmap_54[15:0]) +
	( 16'sd 29380) * $signed(input_fmap_55[15:0]) +
	( 10'sd 306) * $signed(input_fmap_56[15:0]) +
	( 15'sd 15574) * $signed(input_fmap_57[15:0]) +
	( 16'sd 30308) * $signed(input_fmap_58[15:0]) +
	( 12'sd 1780) * $signed(input_fmap_59[15:0]) +
	( 15'sd 12460) * $signed(input_fmap_60[15:0]) +
	( 15'sd 8703) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29512) * $signed(input_fmap_62[15:0]) +
	( 15'sd 9376) * $signed(input_fmap_63[15:0]) +
	( 14'sd 6573) * $signed(input_fmap_64[15:0]) +
	( 16'sd 27285) * $signed(input_fmap_65[15:0]) +
	( 16'sd 28745) * $signed(input_fmap_66[15:0]) +
	( 16'sd 16736) * $signed(input_fmap_67[15:0]) +
	( 11'sd 512) * $signed(input_fmap_68[15:0]) +
	( 12'sd 1794) * $signed(input_fmap_69[15:0]) +
	( 15'sd 15912) * $signed(input_fmap_70[15:0]) +
	( 16'sd 23725) * $signed(input_fmap_71[15:0]) +
	( 14'sd 6341) * $signed(input_fmap_72[15:0]) +
	( 12'sd 1835) * $signed(input_fmap_73[15:0]) +
	( 15'sd 14488) * $signed(input_fmap_74[15:0]) +
	( 16'sd 31528) * $signed(input_fmap_75[15:0]) +
	( 16'sd 21558) * $signed(input_fmap_76[15:0]) +
	( 16'sd 24236) * $signed(input_fmap_77[15:0]) +
	( 14'sd 7479) * $signed(input_fmap_78[15:0]) +
	( 16'sd 26331) * $signed(input_fmap_79[15:0]) +
	( 13'sd 2670) * $signed(input_fmap_80[15:0]) +
	( 15'sd 11805) * $signed(input_fmap_81[15:0]) +
	( 15'sd 14200) * $signed(input_fmap_82[15:0]) +
	( 16'sd 16677) * $signed(input_fmap_83[15:0]) +
	( 16'sd 23849) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24549) * $signed(input_fmap_85[15:0]) +
	( 16'sd 27567) * $signed(input_fmap_86[15:0]) +
	( 14'sd 5056) * $signed(input_fmap_87[15:0]) +
	( 16'sd 32670) * $signed(input_fmap_88[15:0]) +
	( 15'sd 8571) * $signed(input_fmap_89[15:0]) +
	( 16'sd 30623) * $signed(input_fmap_90[15:0]) +
	( 14'sd 4998) * $signed(input_fmap_91[15:0]) +
	( 13'sd 2196) * $signed(input_fmap_92[15:0]) +
	( 16'sd 27751) * $signed(input_fmap_93[15:0]) +
	( 16'sd 23580) * $signed(input_fmap_94[15:0]) +
	( 16'sd 16452) * $signed(input_fmap_95[15:0]) +
	( 15'sd 15629) * $signed(input_fmap_96[15:0]) +
	( 16'sd 30482) * $signed(input_fmap_97[15:0]) +
	( 16'sd 22899) * $signed(input_fmap_98[15:0]) +
	( 13'sd 2272) * $signed(input_fmap_99[15:0]) +
	( 16'sd 29293) * $signed(input_fmap_100[15:0]) +
	( 15'sd 8644) * $signed(input_fmap_101[15:0]) +
	( 14'sd 6231) * $signed(input_fmap_102[15:0]) +
	( 11'sd 692) * $signed(input_fmap_103[15:0]) +
	( 11'sd 523) * $signed(input_fmap_104[15:0]) +
	( 14'sd 6533) * $signed(input_fmap_105[15:0]) +
	( 16'sd 24115) * $signed(input_fmap_106[15:0]) +
	( 16'sd 24012) * $signed(input_fmap_107[15:0]) +
	( 14'sd 5897) * $signed(input_fmap_108[15:0]) +
	( 15'sd 15877) * $signed(input_fmap_109[15:0]) +
	( 15'sd 11658) * $signed(input_fmap_110[15:0]) +
	( 14'sd 7735) * $signed(input_fmap_111[15:0]) +
	( 15'sd 9002) * $signed(input_fmap_112[15:0]) +
	( 14'sd 6722) * $signed(input_fmap_113[15:0]) +
	( 16'sd 23433) * $signed(input_fmap_114[15:0]) +
	( 16'sd 25415) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26849) * $signed(input_fmap_116[15:0]) +
	( 16'sd 18237) * $signed(input_fmap_117[15:0]) +
	( 16'sd 23411) * $signed(input_fmap_118[15:0]) +
	( 14'sd 5971) * $signed(input_fmap_119[15:0]) +
	( 11'sd 741) * $signed(input_fmap_120[15:0]) +
	( 14'sd 7823) * $signed(input_fmap_121[15:0]) +
	( 16'sd 20882) * $signed(input_fmap_122[15:0]) +
	( 16'sd 23886) * $signed(input_fmap_123[15:0]) +
	( 16'sd 26749) * $signed(input_fmap_124[15:0]) +
	( 15'sd 10524) * $signed(input_fmap_125[15:0]) +
	( 15'sd 12459) * $signed(input_fmap_126[15:0]) +
	( 16'sd 25069) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 13'sd 2504) * $signed(input_fmap_0[15:0]) +
	( 16'sd 20566) * $signed(input_fmap_1[15:0]) +
	( 15'sd 16233) * $signed(input_fmap_2[15:0]) +
	( 16'sd 22322) * $signed(input_fmap_3[15:0]) +
	( 13'sd 2102) * $signed(input_fmap_4[15:0]) +
	( 16'sd 30803) * $signed(input_fmap_5[15:0]) +
	( 16'sd 27089) * $signed(input_fmap_6[15:0]) +
	( 15'sd 14608) * $signed(input_fmap_7[15:0]) +
	( 16'sd 32491) * $signed(input_fmap_8[15:0]) +
	( 13'sd 2458) * $signed(input_fmap_9[15:0]) +
	( 16'sd 21177) * $signed(input_fmap_10[15:0]) +
	( 14'sd 6850) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20034) * $signed(input_fmap_12[15:0]) +
	( 16'sd 19822) * $signed(input_fmap_13[15:0]) +
	( 14'sd 7346) * $signed(input_fmap_14[15:0]) +
	( 16'sd 31312) * $signed(input_fmap_15[15:0]) +
	( 14'sd 5386) * $signed(input_fmap_16[15:0]) +
	( 15'sd 15888) * $signed(input_fmap_17[15:0]) +
	( 13'sd 2338) * $signed(input_fmap_18[15:0]) +
	( 13'sd 3900) * $signed(input_fmap_19[15:0]) +
	( 16'sd 26897) * $signed(input_fmap_20[15:0]) +
	( 12'sd 2004) * $signed(input_fmap_21[15:0]) +
	( 16'sd 16506) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28545) * $signed(input_fmap_23[15:0]) +
	( 15'sd 10331) * $signed(input_fmap_24[15:0]) +
	( 15'sd 8405) * $signed(input_fmap_25[15:0]) +
	( 15'sd 13385) * $signed(input_fmap_26[15:0]) +
	( 15'sd 12611) * $signed(input_fmap_27[15:0]) +
	( 15'sd 9375) * $signed(input_fmap_28[15:0]) +
	( 13'sd 3901) * $signed(input_fmap_29[15:0]) +
	( 11'sd 611) * $signed(input_fmap_30[15:0]) +
	( 14'sd 7290) * $signed(input_fmap_31[15:0]) +
	( 15'sd 9502) * $signed(input_fmap_32[15:0]) +
	( 16'sd 27699) * $signed(input_fmap_33[15:0]) +
	( 15'sd 15716) * $signed(input_fmap_34[15:0]) +
	( 13'sd 3520) * $signed(input_fmap_35[15:0]) +
	( 13'sd 3999) * $signed(input_fmap_36[15:0]) +
	( 13'sd 3288) * $signed(input_fmap_37[15:0]) +
	( 16'sd 24179) * $signed(input_fmap_38[15:0]) +
	( 16'sd 27582) * $signed(input_fmap_39[15:0]) +
	( 15'sd 8476) * $signed(input_fmap_40[15:0]) +
	( 16'sd 16520) * $signed(input_fmap_41[15:0]) +
	( 15'sd 8919) * $signed(input_fmap_42[15:0]) +
	( 16'sd 19656) * $signed(input_fmap_43[15:0]) +
	( 15'sd 9027) * $signed(input_fmap_44[15:0]) +
	( 16'sd 22134) * $signed(input_fmap_45[15:0]) +
	( 15'sd 15825) * $signed(input_fmap_46[15:0]) +
	( 16'sd 29177) * $signed(input_fmap_47[15:0]) +
	( 15'sd 14570) * $signed(input_fmap_48[15:0]) +
	( 16'sd 20383) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26461) * $signed(input_fmap_50[15:0]) +
	( 15'sd 16195) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3323) * $signed(input_fmap_52[15:0]) +
	( 15'sd 10196) * $signed(input_fmap_53[15:0]) +
	( 16'sd 16865) * $signed(input_fmap_54[15:0]) +
	( 16'sd 19904) * $signed(input_fmap_55[15:0]) +
	( 8'sd 74) * $signed(input_fmap_56[15:0]) +
	( 16'sd 25530) * $signed(input_fmap_57[15:0]) +
	( 16'sd 22077) * $signed(input_fmap_58[15:0]) +
	( 16'sd 26347) * $signed(input_fmap_59[15:0]) +
	( 16'sd 31932) * $signed(input_fmap_60[15:0]) +
	( 14'sd 5633) * $signed(input_fmap_61[15:0]) +
	( 16'sd 20323) * $signed(input_fmap_62[15:0]) +
	( 16'sd 23516) * $signed(input_fmap_63[15:0]) +
	( 15'sd 14811) * $signed(input_fmap_64[15:0]) +
	( 16'sd 16401) * $signed(input_fmap_65[15:0]) +
	( 16'sd 31294) * $signed(input_fmap_66[15:0]) +
	( 14'sd 6366) * $signed(input_fmap_67[15:0]) +
	( 16'sd 27533) * $signed(input_fmap_68[15:0]) +
	( 16'sd 25632) * $signed(input_fmap_69[15:0]) +
	( 13'sd 3029) * $signed(input_fmap_70[15:0]) +
	( 15'sd 10660) * $signed(input_fmap_71[15:0]) +
	( 16'sd 20314) * $signed(input_fmap_72[15:0]) +
	( 15'sd 16368) * $signed(input_fmap_73[15:0]) +
	( 16'sd 30264) * $signed(input_fmap_74[15:0]) +
	( 15'sd 13919) * $signed(input_fmap_75[15:0]) +
	( 15'sd 13338) * $signed(input_fmap_76[15:0]) +
	( 14'sd 6788) * $signed(input_fmap_77[15:0]) +
	( 16'sd 16777) * $signed(input_fmap_78[15:0]) +
	( 16'sd 23025) * $signed(input_fmap_79[15:0]) +
	( 16'sd 23194) * $signed(input_fmap_80[15:0]) +
	( 11'sd 750) * $signed(input_fmap_81[15:0]) +
	( 15'sd 11721) * $signed(input_fmap_82[15:0]) +
	( 15'sd 10802) * $signed(input_fmap_83[15:0]) +
	( 15'sd 14211) * $signed(input_fmap_84[15:0]) +
	( 16'sd 28962) * $signed(input_fmap_85[15:0]) +
	( 12'sd 1080) * $signed(input_fmap_86[15:0]) +
	( 16'sd 21554) * $signed(input_fmap_87[15:0]) +
	( 14'sd 4218) * $signed(input_fmap_88[15:0]) +
	( 16'sd 23549) * $signed(input_fmap_89[15:0]) +
	( 15'sd 15619) * $signed(input_fmap_90[15:0]) +
	( 16'sd 19013) * $signed(input_fmap_91[15:0]) +
	( 14'sd 6142) * $signed(input_fmap_92[15:0]) +
	( 15'sd 16259) * $signed(input_fmap_93[15:0]) +
	( 15'sd 8641) * $signed(input_fmap_94[15:0]) +
	( 16'sd 24675) * $signed(input_fmap_95[15:0]) +
	( 16'sd 23248) * $signed(input_fmap_96[15:0]) +
	( 15'sd 10073) * $signed(input_fmap_97[15:0]) +
	( 16'sd 20672) * $signed(input_fmap_98[15:0]) +
	( 9'sd 239) * $signed(input_fmap_99[15:0]) +
	( 15'sd 11903) * $signed(input_fmap_100[15:0]) +
	( 16'sd 18448) * $signed(input_fmap_101[15:0]) +
	( 13'sd 2292) * $signed(input_fmap_102[15:0]) +
	( 16'sd 21397) * $signed(input_fmap_103[15:0]) +
	( 16'sd 24214) * $signed(input_fmap_104[15:0]) +
	( 16'sd 30892) * $signed(input_fmap_105[15:0]) +
	( 15'sd 11804) * $signed(input_fmap_106[15:0]) +
	( 16'sd 26158) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15117) * $signed(input_fmap_108[15:0]) +
	( 16'sd 30627) * $signed(input_fmap_109[15:0]) +
	( 16'sd 28106) * $signed(input_fmap_110[15:0]) +
	( 16'sd 21372) * $signed(input_fmap_111[15:0]) +
	( 15'sd 13880) * $signed(input_fmap_112[15:0]) +
	( 16'sd 25093) * $signed(input_fmap_113[15:0]) +
	( 13'sd 3332) * $signed(input_fmap_114[15:0]) +
	( 16'sd 28321) * $signed(input_fmap_115[15:0]) +
	( 15'sd 9839) * $signed(input_fmap_116[15:0]) +
	( 14'sd 5667) * $signed(input_fmap_117[15:0]) +
	( 14'sd 7523) * $signed(input_fmap_118[15:0]) +
	( 14'sd 5171) * $signed(input_fmap_119[15:0]) +
	( 12'sd 1908) * $signed(input_fmap_120[15:0]) +
	( 15'sd 11706) * $signed(input_fmap_121[15:0]) +
	( 14'sd 4984) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21253) * $signed(input_fmap_123[15:0]) +
	( 15'sd 15272) * $signed(input_fmap_124[15:0]) +
	( 16'sd 31985) * $signed(input_fmap_125[15:0]) +
	( 15'sd 14115) * $signed(input_fmap_126[15:0]) +
	( 15'sd 10595) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 16'sd 29650) * $signed(input_fmap_0[15:0]) +
	( 16'sd 28275) * $signed(input_fmap_1[15:0]) +
	( 15'sd 10589) * $signed(input_fmap_2[15:0]) +
	( 16'sd 21228) * $signed(input_fmap_3[15:0]) +
	( 15'sd 15667) * $signed(input_fmap_4[15:0]) +
	( 15'sd 12658) * $signed(input_fmap_5[15:0]) +
	( 16'sd 23314) * $signed(input_fmap_6[15:0]) +
	( 16'sd 21322) * $signed(input_fmap_7[15:0]) +
	( 14'sd 6879) * $signed(input_fmap_8[15:0]) +
	( 16'sd 27907) * $signed(input_fmap_9[15:0]) +
	( 15'sd 13049) * $signed(input_fmap_10[15:0]) +
	( 14'sd 6557) * $signed(input_fmap_11[15:0]) +
	( 16'sd 28884) * $signed(input_fmap_12[15:0]) +
	( 16'sd 16930) * $signed(input_fmap_13[15:0]) +
	( 7'sd 43) * $signed(input_fmap_14[15:0]) +
	( 15'sd 10740) * $signed(input_fmap_15[15:0]) +
	( 16'sd 16462) * $signed(input_fmap_16[15:0]) +
	( 16'sd 26637) * $signed(input_fmap_17[15:0]) +
	( 14'sd 7595) * $signed(input_fmap_18[15:0]) +
	( 13'sd 2418) * $signed(input_fmap_19[15:0]) +
	( 14'sd 7363) * $signed(input_fmap_20[15:0]) +
	( 15'sd 10587) * $signed(input_fmap_21[15:0]) +
	( 14'sd 7950) * $signed(input_fmap_22[15:0]) +
	( 16'sd 21767) * $signed(input_fmap_23[15:0]) +
	( 16'sd 26102) * $signed(input_fmap_24[15:0]) +
	( 16'sd 20023) * $signed(input_fmap_25[15:0]) +
	( 16'sd 31974) * $signed(input_fmap_26[15:0]) +
	( 15'sd 8432) * $signed(input_fmap_27[15:0]) +
	( 15'sd 13962) * $signed(input_fmap_28[15:0]) +
	( 16'sd 24357) * $signed(input_fmap_29[15:0]) +
	( 16'sd 23153) * $signed(input_fmap_30[15:0]) +
	( 16'sd 21371) * $signed(input_fmap_31[15:0]) +
	( 16'sd 31949) * $signed(input_fmap_32[15:0]) +
	( 14'sd 5690) * $signed(input_fmap_33[15:0]) +
	( 13'sd 3976) * $signed(input_fmap_34[15:0]) +
	( 15'sd 10126) * $signed(input_fmap_35[15:0]) +
	( 16'sd 27799) * $signed(input_fmap_36[15:0]) +
	( 16'sd 31596) * $signed(input_fmap_37[15:0]) +
	( 15'sd 14848) * $signed(input_fmap_38[15:0]) +
	( 15'sd 13640) * $signed(input_fmap_39[15:0]) +
	( 15'sd 15837) * $signed(input_fmap_40[15:0]) +
	( 16'sd 16667) * $signed(input_fmap_41[15:0]) +
	( 16'sd 29959) * $signed(input_fmap_42[15:0]) +
	( 16'sd 19683) * $signed(input_fmap_43[15:0]) +
	( 16'sd 22396) * $signed(input_fmap_44[15:0]) +
	( 16'sd 31257) * $signed(input_fmap_45[15:0]) +
	( 16'sd 27418) * $signed(input_fmap_46[15:0]) +
	( 16'sd 31006) * $signed(input_fmap_47[15:0]) +
	( 15'sd 14483) * $signed(input_fmap_48[15:0]) +
	( 16'sd 26856) * $signed(input_fmap_49[15:0]) +
	( 16'sd 24555) * $signed(input_fmap_50[15:0]) +
	( 13'sd 3160) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3132) * $signed(input_fmap_52[15:0]) +
	( 16'sd 18171) * $signed(input_fmap_53[15:0]) +
	( 13'sd 2773) * $signed(input_fmap_54[15:0]) +
	( 15'sd 12518) * $signed(input_fmap_55[15:0]) +
	( 16'sd 27059) * $signed(input_fmap_56[15:0]) +
	( 14'sd 5603) * $signed(input_fmap_57[15:0]) +
	( 16'sd 32331) * $signed(input_fmap_58[15:0]) +
	( 16'sd 22583) * $signed(input_fmap_59[15:0]) +
	( 15'sd 11398) * $signed(input_fmap_60[15:0]) +
	( 16'sd 19941) * $signed(input_fmap_61[15:0]) +
	( 15'sd 13116) * $signed(input_fmap_62[15:0]) +
	( 16'sd 31745) * $signed(input_fmap_63[15:0]) +
	( 13'sd 2248) * $signed(input_fmap_64[15:0]) +
	( 15'sd 11335) * $signed(input_fmap_65[15:0]) +
	( 16'sd 27455) * $signed(input_fmap_66[15:0]) +
	( 16'sd 30404) * $signed(input_fmap_67[15:0]) +
	( 15'sd 12719) * $signed(input_fmap_68[15:0]) +
	( 10'sd 454) * $signed(input_fmap_69[15:0]) +
	( 15'sd 12055) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11003) * $signed(input_fmap_71[15:0]) +
	( 16'sd 26182) * $signed(input_fmap_72[15:0]) +
	( 16'sd 23751) * $signed(input_fmap_73[15:0]) +
	( 16'sd 21685) * $signed(input_fmap_74[15:0]) +
	( 15'sd 14449) * $signed(input_fmap_75[15:0]) +
	( 15'sd 10787) * $signed(input_fmap_76[15:0]) +
	( 16'sd 28163) * $signed(input_fmap_77[15:0]) +
	( 16'sd 25600) * $signed(input_fmap_78[15:0]) +
	( 16'sd 17376) * $signed(input_fmap_79[15:0]) +
	( 16'sd 27785) * $signed(input_fmap_80[15:0]) +
	( 16'sd 19314) * $signed(input_fmap_81[15:0]) +
	( 16'sd 27895) * $signed(input_fmap_82[15:0]) +
	( 15'sd 12127) * $signed(input_fmap_83[15:0]) +
	( 16'sd 18410) * $signed(input_fmap_84[15:0]) +
	( 15'sd 11806) * $signed(input_fmap_85[15:0]) +
	( 15'sd 12856) * $signed(input_fmap_86[15:0]) +
	( 15'sd 13379) * $signed(input_fmap_87[15:0]) +
	( 15'sd 13007) * $signed(input_fmap_88[15:0]) +
	( 16'sd 17486) * $signed(input_fmap_89[15:0]) +
	( 16'sd 18029) * $signed(input_fmap_90[15:0]) +
	( 12'sd 1865) * $signed(input_fmap_91[15:0]) +
	( 16'sd 18827) * $signed(input_fmap_92[15:0]) +
	( 15'sd 15555) * $signed(input_fmap_93[15:0]) +
	( 15'sd 9180) * $signed(input_fmap_94[15:0]) +
	( 15'sd 11963) * $signed(input_fmap_95[15:0]) +
	( 14'sd 6937) * $signed(input_fmap_96[15:0]) +
	( 16'sd 19769) * $signed(input_fmap_97[15:0]) +
	( 16'sd 16775) * $signed(input_fmap_98[15:0]) +
	( 16'sd 30657) * $signed(input_fmap_99[15:0]) +
	( 13'sd 2931) * $signed(input_fmap_100[15:0]) +
	( 16'sd 16827) * $signed(input_fmap_101[15:0]) +
	( 15'sd 15569) * $signed(input_fmap_102[15:0]) +
	( 16'sd 20856) * $signed(input_fmap_103[15:0]) +
	( 15'sd 11935) * $signed(input_fmap_104[15:0]) +
	( 15'sd 13279) * $signed(input_fmap_105[15:0]) +
	( 15'sd 10916) * $signed(input_fmap_106[15:0]) +
	( 16'sd 26959) * $signed(input_fmap_107[15:0]) +
	( 10'sd 507) * $signed(input_fmap_108[15:0]) +
	( 12'sd 1529) * $signed(input_fmap_109[15:0]) +
	( 12'sd 1271) * $signed(input_fmap_110[15:0]) +
	( 16'sd 23787) * $signed(input_fmap_111[15:0]) +
	( 16'sd 27339) * $signed(input_fmap_112[15:0]) +
	( 12'sd 1105) * $signed(input_fmap_113[15:0]) +
	( 16'sd 26364) * $signed(input_fmap_114[15:0]) +
	( 15'sd 10280) * $signed(input_fmap_115[15:0]) +
	( 12'sd 1830) * $signed(input_fmap_116[15:0]) +
	( 16'sd 17382) * $signed(input_fmap_117[15:0]) +
	( 14'sd 4858) * $signed(input_fmap_118[15:0]) +
	( 16'sd 17069) * $signed(input_fmap_119[15:0]) +
	( 14'sd 4700) * $signed(input_fmap_120[15:0]) +
	( 16'sd 16434) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9389) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21028) * $signed(input_fmap_123[15:0]) +
	( 16'sd 26567) * $signed(input_fmap_124[15:0]) +
	( 16'sd 23567) * $signed(input_fmap_125[15:0]) +
	( 15'sd 10999) * $signed(input_fmap_126[15:0]) +
	( 13'sd 2449) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 16'sd 22916) * $signed(input_fmap_0[15:0]) +
	( 11'sd 760) * $signed(input_fmap_1[15:0]) +
	( 15'sd 11050) * $signed(input_fmap_2[15:0]) +
	( 15'sd 14022) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30622) * $signed(input_fmap_4[15:0]) +
	( 16'sd 16525) * $signed(input_fmap_5[15:0]) +
	( 16'sd 21874) * $signed(input_fmap_6[15:0]) +
	( 16'sd 28596) * $signed(input_fmap_7[15:0]) +
	( 16'sd 17766) * $signed(input_fmap_8[15:0]) +
	( 15'sd 13282) * $signed(input_fmap_9[15:0]) +
	( 16'sd 31939) * $signed(input_fmap_10[15:0]) +
	( 15'sd 11605) * $signed(input_fmap_11[15:0]) +
	( 16'sd 23127) * $signed(input_fmap_12[15:0]) +
	( 16'sd 21964) * $signed(input_fmap_13[15:0]) +
	( 16'sd 26781) * $signed(input_fmap_14[15:0]) +
	( 14'sd 7510) * $signed(input_fmap_15[15:0]) +
	( 16'sd 24064) * $signed(input_fmap_16[15:0]) +
	( 15'sd 8317) * $signed(input_fmap_17[15:0]) +
	( 15'sd 14636) * $signed(input_fmap_18[15:0]) +
	( 6'sd 26) * $signed(input_fmap_19[15:0]) +
	( 14'sd 5462) * $signed(input_fmap_20[15:0]) +
	( 16'sd 31346) * $signed(input_fmap_21[15:0]) +
	( 16'sd 20663) * $signed(input_fmap_22[15:0]) +
	( 16'sd 22746) * $signed(input_fmap_23[15:0]) +
	( 16'sd 32245) * $signed(input_fmap_24[15:0]) +
	( 12'sd 1664) * $signed(input_fmap_25[15:0]) +
	( 16'sd 16783) * $signed(input_fmap_26[15:0]) +
	( 16'sd 27623) * $signed(input_fmap_27[15:0]) +
	( 16'sd 23495) * $signed(input_fmap_28[15:0]) +
	( 16'sd 23203) * $signed(input_fmap_29[15:0]) +
	( 16'sd 31668) * $signed(input_fmap_30[15:0]) +
	( 15'sd 14502) * $signed(input_fmap_31[15:0]) +
	( 16'sd 27930) * $signed(input_fmap_32[15:0]) +
	( 16'sd 16566) * $signed(input_fmap_33[15:0]) +
	( 15'sd 9507) * $signed(input_fmap_34[15:0]) +
	( 14'sd 7637) * $signed(input_fmap_35[15:0]) +
	( 14'sd 6532) * $signed(input_fmap_36[15:0]) +
	( 16'sd 28613) * $signed(input_fmap_37[15:0]) +
	( 15'sd 10096) * $signed(input_fmap_38[15:0]) +
	( 16'sd 31278) * $signed(input_fmap_39[15:0]) +
	( 16'sd 31544) * $signed(input_fmap_40[15:0]) +
	( 13'sd 3261) * $signed(input_fmap_41[15:0]) +
	( 15'sd 9658) * $signed(input_fmap_42[15:0]) +
	( 16'sd 23726) * $signed(input_fmap_43[15:0]) +
	( 13'sd 2378) * $signed(input_fmap_44[15:0]) +
	( 16'sd 22242) * $signed(input_fmap_45[15:0]) +
	( 16'sd 18591) * $signed(input_fmap_46[15:0]) +
	( 12'sd 1294) * $signed(input_fmap_47[15:0]) +
	( 16'sd 26647) * $signed(input_fmap_48[15:0]) +
	( 14'sd 4380) * $signed(input_fmap_49[15:0]) +
	( 16'sd 20739) * $signed(input_fmap_50[15:0]) +
	( 15'sd 9386) * $signed(input_fmap_51[15:0]) +
	( 16'sd 24659) * $signed(input_fmap_52[15:0]) +
	( 15'sd 12236) * $signed(input_fmap_53[15:0]) +
	( 16'sd 24566) * $signed(input_fmap_54[15:0]) +
	( 14'sd 6335) * $signed(input_fmap_55[15:0]) +
	( 15'sd 8836) * $signed(input_fmap_56[15:0]) +
	( 14'sd 7746) * $signed(input_fmap_57[15:0]) +
	( 16'sd 22702) * $signed(input_fmap_58[15:0]) +
	( 15'sd 14981) * $signed(input_fmap_59[15:0]) +
	( 13'sd 3850) * $signed(input_fmap_60[15:0]) +
	( 15'sd 13820) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29640) * $signed(input_fmap_62[15:0]) +
	( 14'sd 6710) * $signed(input_fmap_63[15:0]) +
	( 13'sd 2863) * $signed(input_fmap_64[15:0]) +
	( 15'sd 16158) * $signed(input_fmap_65[15:0]) +
	( 14'sd 4559) * $signed(input_fmap_66[15:0]) +
	( 16'sd 29844) * $signed(input_fmap_67[15:0]) +
	( 14'sd 5665) * $signed(input_fmap_68[15:0]) +
	( 16'sd 23136) * $signed(input_fmap_69[15:0]) +
	( 15'sd 9081) * $signed(input_fmap_70[15:0]) +
	( 15'sd 12334) * $signed(input_fmap_71[15:0]) +
	( 14'sd 6238) * $signed(input_fmap_72[15:0]) +
	( 15'sd 13376) * $signed(input_fmap_73[15:0]) +
	( 15'sd 11919) * $signed(input_fmap_74[15:0]) +
	( 16'sd 32155) * $signed(input_fmap_75[15:0]) +
	( 14'sd 5072) * $signed(input_fmap_76[15:0]) +
	( 15'sd 14214) * $signed(input_fmap_77[15:0]) +
	( 15'sd 10949) * $signed(input_fmap_78[15:0]) +
	( 13'sd 3943) * $signed(input_fmap_79[15:0]) +
	( 16'sd 28757) * $signed(input_fmap_80[15:0]) +
	( 14'sd 5012) * $signed(input_fmap_81[15:0]) +
	( 16'sd 17330) * $signed(input_fmap_82[15:0]) +
	( 14'sd 6587) * $signed(input_fmap_83[15:0]) +
	( 11'sd 793) * $signed(input_fmap_84[15:0]) +
	( 15'sd 11273) * $signed(input_fmap_85[15:0]) +
	( 16'sd 20806) * $signed(input_fmap_86[15:0]) +
	( 15'sd 11882) * $signed(input_fmap_87[15:0]) +
	( 16'sd 21739) * $signed(input_fmap_88[15:0]) +
	( 15'sd 15317) * $signed(input_fmap_89[15:0]) +
	( 16'sd 31277) * $signed(input_fmap_90[15:0]) +
	( 16'sd 23976) * $signed(input_fmap_91[15:0]) +
	( 14'sd 7247) * $signed(input_fmap_92[15:0]) +
	( 15'sd 14300) * $signed(input_fmap_93[15:0]) +
	( 14'sd 6703) * $signed(input_fmap_94[15:0]) +
	( 16'sd 18752) * $signed(input_fmap_95[15:0]) +
	( 16'sd 20575) * $signed(input_fmap_96[15:0]) +
	( 16'sd 19179) * $signed(input_fmap_97[15:0]) +
	( 15'sd 12165) * $signed(input_fmap_98[15:0]) +
	( 12'sd 1982) * $signed(input_fmap_99[15:0]) +
	( 15'sd 9307) * $signed(input_fmap_100[15:0]) +
	( 14'sd 6990) * $signed(input_fmap_101[15:0]) +
	( 15'sd 9026) * $signed(input_fmap_102[15:0]) +
	( 16'sd 30615) * $signed(input_fmap_103[15:0]) +
	( 16'sd 22397) * $signed(input_fmap_104[15:0]) +
	( 16'sd 19953) * $signed(input_fmap_105[15:0]) +
	( 14'sd 4405) * $signed(input_fmap_106[15:0]) +
	( 15'sd 12793) * $signed(input_fmap_107[15:0]) +
	( 15'sd 12128) * $signed(input_fmap_108[15:0]) +
	( 16'sd 29592) * $signed(input_fmap_109[15:0]) +
	( 15'sd 9472) * $signed(input_fmap_110[15:0]) +
	( 16'sd 30448) * $signed(input_fmap_111[15:0]) +
	( 15'sd 10213) * $signed(input_fmap_112[15:0]) +
	( 16'sd 28375) * $signed(input_fmap_113[15:0]) +
	( 16'sd 30843) * $signed(input_fmap_114[15:0]) +
	( 13'sd 3748) * $signed(input_fmap_115[15:0]) +
	( 16'sd 28163) * $signed(input_fmap_116[15:0]) +
	( 15'sd 8421) * $signed(input_fmap_117[15:0]) +
	( 16'sd 20840) * $signed(input_fmap_118[15:0]) +
	( 16'sd 28086) * $signed(input_fmap_119[15:0]) +
	( 14'sd 8019) * $signed(input_fmap_120[15:0]) +
	( 15'sd 12118) * $signed(input_fmap_121[15:0]) +
	( 15'sd 11926) * $signed(input_fmap_122[15:0]) +
	( 15'sd 10667) * $signed(input_fmap_123[15:0]) +
	( 14'sd 5855) * $signed(input_fmap_124[15:0]) +
	( 16'sd 31962) * $signed(input_fmap_125[15:0]) +
	( 16'sd 27731) * $signed(input_fmap_126[15:0]) +
	( 14'sd 5656) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 13'sd 3654) * $signed(input_fmap_0[15:0]) +
	( 16'sd 30591) * $signed(input_fmap_1[15:0]) +
	( 12'sd 1959) * $signed(input_fmap_2[15:0]) +
	( 15'sd 15128) * $signed(input_fmap_3[15:0]) +
	( 12'sd 1783) * $signed(input_fmap_4[15:0]) +
	( 16'sd 26355) * $signed(input_fmap_5[15:0]) +
	( 15'sd 10427) * $signed(input_fmap_6[15:0]) +
	( 16'sd 27931) * $signed(input_fmap_7[15:0]) +
	( 16'sd 27416) * $signed(input_fmap_8[15:0]) +
	( 14'sd 6063) * $signed(input_fmap_9[15:0]) +
	( 16'sd 30743) * $signed(input_fmap_10[15:0]) +
	( 15'sd 14880) * $signed(input_fmap_11[15:0]) +
	( 16'sd 30927) * $signed(input_fmap_12[15:0]) +
	( 16'sd 23456) * $signed(input_fmap_13[15:0]) +
	( 16'sd 25831) * $signed(input_fmap_14[15:0]) +
	( 16'sd 17134) * $signed(input_fmap_15[15:0]) +
	( 14'sd 5415) * $signed(input_fmap_16[15:0]) +
	( 16'sd 19323) * $signed(input_fmap_17[15:0]) +
	( 15'sd 11026) * $signed(input_fmap_18[15:0]) +
	( 16'sd 18034) * $signed(input_fmap_19[15:0]) +
	( 15'sd 12927) * $signed(input_fmap_20[15:0]) +
	( 13'sd 2064) * $signed(input_fmap_21[15:0]) +
	( 15'sd 8508) * $signed(input_fmap_22[15:0]) +
	( 13'sd 3564) * $signed(input_fmap_23[15:0]) +
	( 14'sd 5604) * $signed(input_fmap_24[15:0]) +
	( 10'sd 333) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22403) * $signed(input_fmap_26[15:0]) +
	( 16'sd 16913) * $signed(input_fmap_27[15:0]) +
	( 14'sd 5048) * $signed(input_fmap_28[15:0]) +
	( 16'sd 30152) * $signed(input_fmap_29[15:0]) +
	( 15'sd 9250) * $signed(input_fmap_30[15:0]) +
	( 16'sd 29515) * $signed(input_fmap_31[15:0]) +
	( 11'sd 582) * $signed(input_fmap_32[15:0]) +
	( 16'sd 28912) * $signed(input_fmap_33[15:0]) +
	( 14'sd 6714) * $signed(input_fmap_34[15:0]) +
	( 16'sd 20564) * $signed(input_fmap_35[15:0]) +
	( 15'sd 13079) * $signed(input_fmap_36[15:0]) +
	( 16'sd 17551) * $signed(input_fmap_37[15:0]) +
	( 16'sd 19386) * $signed(input_fmap_38[15:0]) +
	( 16'sd 21755) * $signed(input_fmap_39[15:0]) +
	( 16'sd 18224) * $signed(input_fmap_40[15:0]) +
	( 16'sd 24148) * $signed(input_fmap_41[15:0]) +
	( 15'sd 15150) * $signed(input_fmap_43[15:0]) +
	( 16'sd 23202) * $signed(input_fmap_44[15:0]) +
	( 11'sd 932) * $signed(input_fmap_45[15:0]) +
	( 14'sd 7156) * $signed(input_fmap_46[15:0]) +
	( 16'sd 27058) * $signed(input_fmap_47[15:0]) +
	( 13'sd 3747) * $signed(input_fmap_48[15:0]) +
	( 15'sd 14500) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22966) * $signed(input_fmap_50[15:0]) +
	( 15'sd 9051) * $signed(input_fmap_51[15:0]) +
	( 16'sd 22149) * $signed(input_fmap_52[15:0]) +
	( 15'sd 8445) * $signed(input_fmap_53[15:0]) +
	( 14'sd 4318) * $signed(input_fmap_54[15:0]) +
	( 16'sd 32605) * $signed(input_fmap_55[15:0]) +
	( 15'sd 15443) * $signed(input_fmap_56[15:0]) +
	( 16'sd 28000) * $signed(input_fmap_57[15:0]) +
	( 14'sd 5315) * $signed(input_fmap_58[15:0]) +
	( 16'sd 17470) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1872) * $signed(input_fmap_60[15:0]) +
	( 15'sd 13120) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3488) * $signed(input_fmap_62[15:0]) +
	( 16'sd 28340) * $signed(input_fmap_63[15:0]) +
	( 16'sd 24820) * $signed(input_fmap_64[15:0]) +
	( 14'sd 7607) * $signed(input_fmap_65[15:0]) +
	( 16'sd 24615) * $signed(input_fmap_66[15:0]) +
	( 16'sd 32423) * $signed(input_fmap_67[15:0]) +
	( 14'sd 4814) * $signed(input_fmap_68[15:0]) +
	( 16'sd 16596) * $signed(input_fmap_69[15:0]) +
	( 16'sd 31954) * $signed(input_fmap_70[15:0]) +
	( 14'sd 5793) * $signed(input_fmap_71[15:0]) +
	( 13'sd 2536) * $signed(input_fmap_72[15:0]) +
	( 14'sd 4546) * $signed(input_fmap_73[15:0]) +
	( 15'sd 8345) * $signed(input_fmap_74[15:0]) +
	( 16'sd 18602) * $signed(input_fmap_75[15:0]) +
	( 15'sd 13379) * $signed(input_fmap_76[15:0]) +
	( 15'sd 14923) * $signed(input_fmap_77[15:0]) +
	( 16'sd 30213) * $signed(input_fmap_78[15:0]) +
	( 16'sd 30776) * $signed(input_fmap_79[15:0]) +
	( 16'sd 25154) * $signed(input_fmap_80[15:0]) +
	( 16'sd 28375) * $signed(input_fmap_81[15:0]) +
	( 14'sd 8156) * $signed(input_fmap_82[15:0]) +
	( 16'sd 23632) * $signed(input_fmap_83[15:0]) +
	( 13'sd 3481) * $signed(input_fmap_84[15:0]) +
	( 16'sd 26224) * $signed(input_fmap_85[15:0]) +
	( 15'sd 10091) * $signed(input_fmap_86[15:0]) +
	( 16'sd 16581) * $signed(input_fmap_87[15:0]) +
	( 13'sd 3315) * $signed(input_fmap_88[15:0]) +
	( 16'sd 23950) * $signed(input_fmap_89[15:0]) +
	( 15'sd 11833) * $signed(input_fmap_90[15:0]) +
	( 14'sd 6802) * $signed(input_fmap_91[15:0]) +
	( 14'sd 4101) * $signed(input_fmap_92[15:0]) +
	( 15'sd 13217) * $signed(input_fmap_93[15:0]) +
	( 16'sd 21727) * $signed(input_fmap_94[15:0]) +
	( 15'sd 12952) * $signed(input_fmap_95[15:0]) +
	( 16'sd 29356) * $signed(input_fmap_96[15:0]) +
	( 16'sd 25481) * $signed(input_fmap_97[15:0]) +
	( 15'sd 13580) * $signed(input_fmap_98[15:0]) +
	( 13'sd 2927) * $signed(input_fmap_99[15:0]) +
	( 14'sd 6315) * $signed(input_fmap_100[15:0]) +
	( 15'sd 16369) * $signed(input_fmap_101[15:0]) +
	( 13'sd 3558) * $signed(input_fmap_102[15:0]) +
	( 15'sd 10387) * $signed(input_fmap_103[15:0]) +
	( 16'sd 23953) * $signed(input_fmap_104[15:0]) +
	( 16'sd 23824) * $signed(input_fmap_105[15:0]) +
	( 16'sd 26737) * $signed(input_fmap_106[15:0]) +
	( 14'sd 6538) * $signed(input_fmap_107[15:0]) +
	( 16'sd 21135) * $signed(input_fmap_108[15:0]) +
	( 15'sd 12857) * $signed(input_fmap_109[15:0]) +
	( 15'sd 10723) * $signed(input_fmap_110[15:0]) +
	( 16'sd 21938) * $signed(input_fmap_111[15:0]) +
	( 13'sd 3300) * $signed(input_fmap_112[15:0]) +
	( 16'sd 23990) * $signed(input_fmap_113[15:0]) +
	( 16'sd 20134) * $signed(input_fmap_114[15:0]) +
	( 15'sd 14176) * $signed(input_fmap_115[15:0]) +
	( 16'sd 25964) * $signed(input_fmap_116[15:0]) +
	( 16'sd 31712) * $signed(input_fmap_117[15:0]) +
	( 14'sd 5815) * $signed(input_fmap_118[15:0]) +
	( 14'sd 6583) * $signed(input_fmap_119[15:0]) +
	( 12'sd 1638) * $signed(input_fmap_120[15:0]) +
	( 16'sd 23463) * $signed(input_fmap_121[15:0]) +
	( 15'sd 13009) * $signed(input_fmap_122[15:0]) +
	( 16'sd 31540) * $signed(input_fmap_123[15:0]) +
	( 16'sd 31478) * $signed(input_fmap_124[15:0]) +
	( 16'sd 17693) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6395) * $signed(input_fmap_126[15:0]) +
	( 16'sd 21359) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 9'sd 156) * $signed(input_fmap_0[15:0]) +
	( 16'sd 20469) * $signed(input_fmap_1[15:0]) +
	( 15'sd 9607) * $signed(input_fmap_2[15:0]) +
	( 15'sd 11364) * $signed(input_fmap_3[15:0]) +
	( 15'sd 13139) * $signed(input_fmap_4[15:0]) +
	( 16'sd 23701) * $signed(input_fmap_5[15:0]) +
	( 16'sd 32187) * $signed(input_fmap_6[15:0]) +
	( 16'sd 18083) * $signed(input_fmap_7[15:0]) +
	( 15'sd 16312) * $signed(input_fmap_8[15:0]) +
	( 16'sd 23578) * $signed(input_fmap_9[15:0]) +
	( 16'sd 20157) * $signed(input_fmap_10[15:0]) +
	( 13'sd 2625) * $signed(input_fmap_11[15:0]) +
	( 14'sd 7441) * $signed(input_fmap_12[15:0]) +
	( 16'sd 30043) * $signed(input_fmap_13[15:0]) +
	( 16'sd 23813) * $signed(input_fmap_14[15:0]) +
	( 11'sd 526) * $signed(input_fmap_15[15:0]) +
	( 16'sd 26294) * $signed(input_fmap_16[15:0]) +
	( 13'sd 2551) * $signed(input_fmap_17[15:0]) +
	( 16'sd 18254) * $signed(input_fmap_18[15:0]) +
	( 15'sd 8950) * $signed(input_fmap_19[15:0]) +
	( 16'sd 29428) * $signed(input_fmap_20[15:0]) +
	( 16'sd 31401) * $signed(input_fmap_21[15:0]) +
	( 13'sd 3967) * $signed(input_fmap_22[15:0]) +
	( 15'sd 12477) * $signed(input_fmap_23[15:0]) +
	( 15'sd 13503) * $signed(input_fmap_24[15:0]) +
	( 16'sd 27914) * $signed(input_fmap_25[15:0]) +
	( 12'sd 1402) * $signed(input_fmap_26[15:0]) +
	( 16'sd 20224) * $signed(input_fmap_27[15:0]) +
	( 15'sd 15189) * $signed(input_fmap_28[15:0]) +
	( 16'sd 18569) * $signed(input_fmap_29[15:0]) +
	( 14'sd 4351) * $signed(input_fmap_30[15:0]) +
	( 14'sd 6124) * $signed(input_fmap_31[15:0]) +
	( 14'sd 5891) * $signed(input_fmap_32[15:0]) +
	( 16'sd 22899) * $signed(input_fmap_33[15:0]) +
	( 16'sd 31976) * $signed(input_fmap_34[15:0]) +
	( 15'sd 9874) * $signed(input_fmap_35[15:0]) +
	( 16'sd 26691) * $signed(input_fmap_36[15:0]) +
	( 16'sd 31151) * $signed(input_fmap_37[15:0]) +
	( 16'sd 28370) * $signed(input_fmap_38[15:0]) +
	( 11'sd 616) * $signed(input_fmap_39[15:0]) +
	( 16'sd 23181) * $signed(input_fmap_40[15:0]) +
	( 15'sd 10326) * $signed(input_fmap_41[15:0]) +
	( 16'sd 26113) * $signed(input_fmap_42[15:0]) +
	( 16'sd 20041) * $signed(input_fmap_43[15:0]) +
	( 13'sd 2680) * $signed(input_fmap_44[15:0]) +
	( 11'sd 698) * $signed(input_fmap_45[15:0]) +
	( 14'sd 4628) * $signed(input_fmap_46[15:0]) +
	( 16'sd 29082) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13817) * $signed(input_fmap_48[15:0]) +
	( 13'sd 3268) * $signed(input_fmap_49[15:0]) +
	( 16'sd 20187) * $signed(input_fmap_50[15:0]) +
	( 16'sd 21983) * $signed(input_fmap_51[15:0]) +
	( 16'sd 23733) * $signed(input_fmap_52[15:0]) +
	( 16'sd 25104) * $signed(input_fmap_53[15:0]) +
	( 14'sd 7316) * $signed(input_fmap_54[15:0]) +
	( 15'sd 14521) * $signed(input_fmap_55[15:0]) +
	( 14'sd 6254) * $signed(input_fmap_56[15:0]) +
	( 16'sd 29419) * $signed(input_fmap_57[15:0]) +
	( 13'sd 2369) * $signed(input_fmap_58[15:0]) +
	( 13'sd 3430) * $signed(input_fmap_59[15:0]) +
	( 14'sd 4257) * $signed(input_fmap_60[15:0]) +
	( 15'sd 8197) * $signed(input_fmap_61[15:0]) +
	( 16'sd 23023) * $signed(input_fmap_62[15:0]) +
	( 16'sd 19997) * $signed(input_fmap_63[15:0]) +
	( 16'sd 22128) * $signed(input_fmap_64[15:0]) +
	( 16'sd 28949) * $signed(input_fmap_65[15:0]) +
	( 16'sd 23365) * $signed(input_fmap_66[15:0]) +
	( 15'sd 13023) * $signed(input_fmap_67[15:0]) +
	( 15'sd 12749) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31438) * $signed(input_fmap_69[15:0]) +
	( 16'sd 30360) * $signed(input_fmap_70[15:0]) +
	( 16'sd 28249) * $signed(input_fmap_71[15:0]) +
	( 16'sd 25871) * $signed(input_fmap_72[15:0]) +
	( 15'sd 10939) * $signed(input_fmap_73[15:0]) +
	( 14'sd 4766) * $signed(input_fmap_74[15:0]) +
	( 16'sd 28373) * $signed(input_fmap_75[15:0]) +
	( 15'sd 14163) * $signed(input_fmap_76[15:0]) +
	( 15'sd 8309) * $signed(input_fmap_77[15:0]) +
	( 16'sd 24293) * $signed(input_fmap_78[15:0]) +
	( 15'sd 12062) * $signed(input_fmap_79[15:0]) +
	( 15'sd 15238) * $signed(input_fmap_80[15:0]) +
	( 16'sd 23317) * $signed(input_fmap_81[15:0]) +
	( 15'sd 11684) * $signed(input_fmap_82[15:0]) +
	( 16'sd 29187) * $signed(input_fmap_83[15:0]) +
	( 16'sd 19010) * $signed(input_fmap_84[15:0]) +
	( 15'sd 10795) * $signed(input_fmap_85[15:0]) +
	( 13'sd 2105) * $signed(input_fmap_86[15:0]) +
	( 16'sd 32421) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6172) * $signed(input_fmap_88[15:0]) +
	( 16'sd 18697) * $signed(input_fmap_89[15:0]) +
	( 16'sd 23204) * $signed(input_fmap_90[15:0]) +
	( 16'sd 20458) * $signed(input_fmap_91[15:0]) +
	( 16'sd 29746) * $signed(input_fmap_92[15:0]) +
	( 14'sd 6728) * $signed(input_fmap_93[15:0]) +
	( 14'sd 4841) * $signed(input_fmap_94[15:0]) +
	( 14'sd 4510) * $signed(input_fmap_95[15:0]) +
	( 14'sd 4936) * $signed(input_fmap_96[15:0]) +
	( 15'sd 15561) * $signed(input_fmap_97[15:0]) +
	( 16'sd 21423) * $signed(input_fmap_98[15:0]) +
	( 15'sd 10710) * $signed(input_fmap_99[15:0]) +
	( 15'sd 14393) * $signed(input_fmap_100[15:0]) +
	( 16'sd 32042) * $signed(input_fmap_101[15:0]) +
	( 16'sd 29725) * $signed(input_fmap_102[15:0]) +
	( 15'sd 13492) * $signed(input_fmap_103[15:0]) +
	( 15'sd 14527) * $signed(input_fmap_104[15:0]) +
	( 14'sd 6164) * $signed(input_fmap_105[15:0]) +
	( 15'sd 10949) * $signed(input_fmap_106[15:0]) +
	( 13'sd 2852) * $signed(input_fmap_107[15:0]) +
	( 16'sd 16385) * $signed(input_fmap_108[15:0]) +
	( 15'sd 16365) * $signed(input_fmap_109[15:0]) +
	( 16'sd 27896) * $signed(input_fmap_110[15:0]) +
	( 16'sd 25005) * $signed(input_fmap_111[15:0]) +
	( 15'sd 10942) * $signed(input_fmap_112[15:0]) +
	( 16'sd 30861) * $signed(input_fmap_113[15:0]) +
	( 14'sd 8040) * $signed(input_fmap_114[15:0]) +
	( 16'sd 31344) * $signed(input_fmap_115[15:0]) +
	( 16'sd 32381) * $signed(input_fmap_116[15:0]) +
	( 16'sd 31257) * $signed(input_fmap_117[15:0]) +
	( 16'sd 19698) * $signed(input_fmap_118[15:0]) +
	( 16'sd 25281) * $signed(input_fmap_119[15:0]) +
	( 14'sd 8153) * $signed(input_fmap_120[15:0]) +
	( 15'sd 16089) * $signed(input_fmap_121[15:0]) +
	( 16'sd 28987) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21209) * $signed(input_fmap_123[15:0]) +
	( 16'sd 24360) * $signed(input_fmap_124[15:0]) +
	( 16'sd 19896) * $signed(input_fmap_125[15:0]) +
	( 16'sd 17506) * $signed(input_fmap_126[15:0]) +
	( 16'sd 25105) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 16'sd 24757) * $signed(input_fmap_0[15:0]) +
	( 15'sd 13148) * $signed(input_fmap_1[15:0]) +
	( 16'sd 17210) * $signed(input_fmap_2[15:0]) +
	( 16'sd 30749) * $signed(input_fmap_3[15:0]) +
	( 14'sd 8146) * $signed(input_fmap_4[15:0]) +
	( 14'sd 7286) * $signed(input_fmap_5[15:0]) +
	( 16'sd 19779) * $signed(input_fmap_6[15:0]) +
	( 16'sd 26855) * $signed(input_fmap_7[15:0]) +
	( 16'sd 26831) * $signed(input_fmap_8[15:0]) +
	( 15'sd 11903) * $signed(input_fmap_9[15:0]) +
	( 16'sd 26109) * $signed(input_fmap_10[15:0]) +
	( 16'sd 21705) * $signed(input_fmap_11[15:0]) +
	( 16'sd 27910) * $signed(input_fmap_12[15:0]) +
	( 16'sd 28288) * $signed(input_fmap_13[15:0]) +
	( 16'sd 27536) * $signed(input_fmap_14[15:0]) +
	( 16'sd 17995) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10412) * $signed(input_fmap_16[15:0]) +
	( 16'sd 21220) * $signed(input_fmap_17[15:0]) +
	( 16'sd 32106) * $signed(input_fmap_18[15:0]) +
	( 16'sd 19880) * $signed(input_fmap_19[15:0]) +
	( 16'sd 30031) * $signed(input_fmap_20[15:0]) +
	( 12'sd 1756) * $signed(input_fmap_21[15:0]) +
	( 12'sd 1733) * $signed(input_fmap_22[15:0]) +
	( 16'sd 30657) * $signed(input_fmap_23[15:0]) +
	( 16'sd 29012) * $signed(input_fmap_24[15:0]) +
	( 16'sd 25972) * $signed(input_fmap_25[15:0]) +
	( 16'sd 19678) * $signed(input_fmap_26[15:0]) +
	( 14'sd 4866) * $signed(input_fmap_27[15:0]) +
	( 16'sd 31179) * $signed(input_fmap_28[15:0]) +
	( 15'sd 14086) * $signed(input_fmap_29[15:0]) +
	( 13'sd 3904) * $signed(input_fmap_30[15:0]) +
	( 14'sd 7447) * $signed(input_fmap_31[15:0]) +
	( 16'sd 16420) * $signed(input_fmap_32[15:0]) +
	( 11'sd 801) * $signed(input_fmap_33[15:0]) +
	( 16'sd 19516) * $signed(input_fmap_34[15:0]) +
	( 15'sd 10013) * $signed(input_fmap_35[15:0]) +
	( 15'sd 14140) * $signed(input_fmap_36[15:0]) +
	( 16'sd 24971) * $signed(input_fmap_37[15:0]) +
	( 14'sd 4907) * $signed(input_fmap_38[15:0]) +
	( 16'sd 30818) * $signed(input_fmap_39[15:0]) +
	( 16'sd 27837) * $signed(input_fmap_40[15:0]) +
	( 16'sd 23388) * $signed(input_fmap_41[15:0]) +
	( 15'sd 9465) * $signed(input_fmap_42[15:0]) +
	( 16'sd 21865) * $signed(input_fmap_43[15:0]) +
	( 16'sd 26379) * $signed(input_fmap_44[15:0]) +
	( 15'sd 9969) * $signed(input_fmap_45[15:0]) +
	( 15'sd 15824) * $signed(input_fmap_46[15:0]) +
	( 11'sd 543) * $signed(input_fmap_47[15:0]) +
	( 16'sd 24728) * $signed(input_fmap_48[15:0]) +
	( 15'sd 8800) * $signed(input_fmap_49[15:0]) +
	( 12'sd 2019) * $signed(input_fmap_50[15:0]) +
	( 16'sd 21049) * $signed(input_fmap_51[15:0]) +
	( 14'sd 5519) * $signed(input_fmap_52[15:0]) +
	( 13'sd 2681) * $signed(input_fmap_53[15:0]) +
	( 14'sd 4467) * $signed(input_fmap_54[15:0]) +
	( 16'sd 22190) * $signed(input_fmap_55[15:0]) +
	( 16'sd 28066) * $signed(input_fmap_56[15:0]) +
	( 15'sd 15992) * $signed(input_fmap_57[15:0]) +
	( 14'sd 7322) * $signed(input_fmap_58[15:0]) +
	( 16'sd 17806) * $signed(input_fmap_59[15:0]) +
	( 13'sd 2126) * $signed(input_fmap_60[15:0]) +
	( 14'sd 6986) * $signed(input_fmap_61[15:0]) +
	( 16'sd 29236) * $signed(input_fmap_62[15:0]) +
	( 16'sd 27108) * $signed(input_fmap_63[15:0]) +
	( 14'sd 4988) * $signed(input_fmap_64[15:0]) +
	( 10'sd 414) * $signed(input_fmap_65[15:0]) +
	( 14'sd 6612) * $signed(input_fmap_66[15:0]) +
	( 16'sd 25455) * $signed(input_fmap_67[15:0]) +
	( 15'sd 11561) * $signed(input_fmap_68[15:0]) +
	( 16'sd 23147) * $signed(input_fmap_69[15:0]) +
	( 14'sd 5361) * $signed(input_fmap_70[15:0]) +
	( 16'sd 27499) * $signed(input_fmap_71[15:0]) +
	( 16'sd 21645) * $signed(input_fmap_72[15:0]) +
	( 16'sd 21783) * $signed(input_fmap_73[15:0]) +
	( 16'sd 28860) * $signed(input_fmap_74[15:0]) +
	( 16'sd 24763) * $signed(input_fmap_75[15:0]) +
	( 15'sd 14770) * $signed(input_fmap_76[15:0]) +
	( 16'sd 17117) * $signed(input_fmap_77[15:0]) +
	( 16'sd 30223) * $signed(input_fmap_78[15:0]) +
	( 16'sd 28060) * $signed(input_fmap_79[15:0]) +
	( 13'sd 3408) * $signed(input_fmap_80[15:0]) +
	( 16'sd 19264) * $signed(input_fmap_81[15:0]) +
	( 16'sd 31497) * $signed(input_fmap_82[15:0]) +
	( 15'sd 11529) * $signed(input_fmap_83[15:0]) +
	( 13'sd 3809) * $signed(input_fmap_84[15:0]) +
	( 16'sd 25169) * $signed(input_fmap_85[15:0]) +
	( 15'sd 16034) * $signed(input_fmap_86[15:0]) +
	( 15'sd 10335) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6138) * $signed(input_fmap_88[15:0]) +
	( 11'sd 752) * $signed(input_fmap_89[15:0]) +
	( 15'sd 9947) * $signed(input_fmap_90[15:0]) +
	( 15'sd 9410) * $signed(input_fmap_91[15:0]) +
	( 16'sd 19240) * $signed(input_fmap_92[15:0]) +
	( 16'sd 17023) * $signed(input_fmap_93[15:0]) +
	( 16'sd 23289) * $signed(input_fmap_94[15:0]) +
	( 16'sd 26878) * $signed(input_fmap_95[15:0]) +
	( 13'sd 3570) * $signed(input_fmap_96[15:0]) +
	( 16'sd 29976) * $signed(input_fmap_97[15:0]) +
	( 15'sd 13111) * $signed(input_fmap_98[15:0]) +
	( 15'sd 11678) * $signed(input_fmap_99[15:0]) +
	( 15'sd 14212) * $signed(input_fmap_100[15:0]) +
	( 16'sd 20766) * $signed(input_fmap_101[15:0]) +
	( 15'sd 12589) * $signed(input_fmap_102[15:0]) +
	( 16'sd 26457) * $signed(input_fmap_103[15:0]) +
	( 16'sd 29135) * $signed(input_fmap_104[15:0]) +
	( 12'sd 1734) * $signed(input_fmap_105[15:0]) +
	( 16'sd 31468) * $signed(input_fmap_106[15:0]) +
	( 15'sd 12892) * $signed(input_fmap_107[15:0]) +
	( 16'sd 29227) * $signed(input_fmap_108[15:0]) +
	( 16'sd 18514) * $signed(input_fmap_109[15:0]) +
	( 16'sd 21639) * $signed(input_fmap_110[15:0]) +
	( 16'sd 21150) * $signed(input_fmap_111[15:0]) +
	( 12'sd 1855) * $signed(input_fmap_112[15:0]) +
	( 13'sd 3176) * $signed(input_fmap_113[15:0]) +
	( 15'sd 14112) * $signed(input_fmap_114[15:0]) +
	( 11'sd 667) * $signed(input_fmap_115[15:0]) +
	( 16'sd 24524) * $signed(input_fmap_116[15:0]) +
	( 16'sd 22586) * $signed(input_fmap_117[15:0]) +
	( 15'sd 11500) * $signed(input_fmap_118[15:0]) +
	( 15'sd 9368) * $signed(input_fmap_119[15:0]) +
	( 14'sd 7360) * $signed(input_fmap_120[15:0]) +
	( 15'sd 12514) * $signed(input_fmap_121[15:0]) +
	( 15'sd 12237) * $signed(input_fmap_122[15:0]) +
	( 15'sd 12158) * $signed(input_fmap_123[15:0]) +
	( 15'sd 11104) * $signed(input_fmap_124[15:0]) +
	( 14'sd 7701) * $signed(input_fmap_125[15:0]) +
	( 14'sd 4148) * $signed(input_fmap_126[15:0]) +
	( 16'sd 19376) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 15'sd 8246) * $signed(input_fmap_0[15:0]) +
	( 15'sd 16125) * $signed(input_fmap_1[15:0]) +
	( 16'sd 20691) * $signed(input_fmap_2[15:0]) +
	( 15'sd 10745) * $signed(input_fmap_3[15:0]) +
	( 14'sd 4339) * $signed(input_fmap_4[15:0]) +
	( 13'sd 2588) * $signed(input_fmap_5[15:0]) +
	( 16'sd 29575) * $signed(input_fmap_6[15:0]) +
	( 14'sd 5191) * $signed(input_fmap_7[15:0]) +
	( 15'sd 12560) * $signed(input_fmap_8[15:0]) +
	( 16'sd 22861) * $signed(input_fmap_9[15:0]) +
	( 16'sd 25703) * $signed(input_fmap_10[15:0]) +
	( 16'sd 28552) * $signed(input_fmap_11[15:0]) +
	( 16'sd 19031) * $signed(input_fmap_12[15:0]) +
	( 16'sd 28380) * $signed(input_fmap_13[15:0]) +
	( 12'sd 1323) * $signed(input_fmap_14[15:0]) +
	( 15'sd 15097) * $signed(input_fmap_15[15:0]) +
	( 16'sd 22914) * $signed(input_fmap_16[15:0]) +
	( 16'sd 24815) * $signed(input_fmap_17[15:0]) +
	( 14'sd 8116) * $signed(input_fmap_18[15:0]) +
	( 16'sd 22607) * $signed(input_fmap_19[15:0]) +
	( 13'sd 2185) * $signed(input_fmap_20[15:0]) +
	( 16'sd 31110) * $signed(input_fmap_21[15:0]) +
	( 15'sd 15365) * $signed(input_fmap_22[15:0]) +
	( 16'sd 29908) * $signed(input_fmap_23[15:0]) +
	( 16'sd 20570) * $signed(input_fmap_24[15:0]) +
	( 15'sd 10015) * $signed(input_fmap_25[15:0]) +
	( 16'sd 20558) * $signed(input_fmap_26[15:0]) +
	( 16'sd 21974) * $signed(input_fmap_27[15:0]) +
	( 14'sd 4295) * $signed(input_fmap_28[15:0]) +
	( 13'sd 2261) * $signed(input_fmap_29[15:0]) +
	( 14'sd 6938) * $signed(input_fmap_30[15:0]) +
	( 16'sd 19116) * $signed(input_fmap_31[15:0]) +
	( 16'sd 24872) * $signed(input_fmap_32[15:0]) +
	( 14'sd 7900) * $signed(input_fmap_33[15:0]) +
	( 12'sd 1445) * $signed(input_fmap_34[15:0]) +
	( 16'sd 22734) * $signed(input_fmap_35[15:0]) +
	( 15'sd 9997) * $signed(input_fmap_36[15:0]) +
	( 16'sd 19411) * $signed(input_fmap_37[15:0]) +
	( 16'sd 16806) * $signed(input_fmap_38[15:0]) +
	( 14'sd 7535) * $signed(input_fmap_39[15:0]) +
	( 16'sd 25470) * $signed(input_fmap_40[15:0]) +
	( 10'sd 355) * $signed(input_fmap_41[15:0]) +
	( 14'sd 4978) * $signed(input_fmap_42[15:0]) +
	( 16'sd 16531) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31131) * $signed(input_fmap_44[15:0]) +
	( 16'sd 28273) * $signed(input_fmap_45[15:0]) +
	( 14'sd 4648) * $signed(input_fmap_46[15:0]) +
	( 15'sd 11991) * $signed(input_fmap_47[15:0]) +
	( 16'sd 19058) * $signed(input_fmap_48[15:0]) +
	( 15'sd 11346) * $signed(input_fmap_49[15:0]) +
	( 16'sd 17065) * $signed(input_fmap_50[15:0]) +
	( 16'sd 27075) * $signed(input_fmap_51[15:0]) +
	( 16'sd 22468) * $signed(input_fmap_52[15:0]) +
	( 16'sd 25877) * $signed(input_fmap_53[15:0]) +
	( 16'sd 16726) * $signed(input_fmap_54[15:0]) +
	( 16'sd 30153) * $signed(input_fmap_55[15:0]) +
	( 16'sd 24390) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17529) * $signed(input_fmap_57[15:0]) +
	( 9'sd 156) * $signed(input_fmap_58[15:0]) +
	( 11'sd 896) * $signed(input_fmap_59[15:0]) +
	( 15'sd 12383) * $signed(input_fmap_60[15:0]) +
	( 16'sd 32211) * $signed(input_fmap_61[15:0]) +
	( 16'sd 19349) * $signed(input_fmap_62[15:0]) +
	( 16'sd 30847) * $signed(input_fmap_63[15:0]) +
	( 12'sd 1415) * $signed(input_fmap_64[15:0]) +
	( 16'sd 22617) * $signed(input_fmap_65[15:0]) +
	( 14'sd 4792) * $signed(input_fmap_66[15:0]) +
	( 16'sd 29645) * $signed(input_fmap_67[15:0]) +
	( 12'sd 1620) * $signed(input_fmap_68[15:0]) +
	( 14'sd 5758) * $signed(input_fmap_69[15:0]) +
	( 14'sd 6969) * $signed(input_fmap_70[15:0]) +
	( 16'sd 17124) * $signed(input_fmap_71[15:0]) +
	( 16'sd 19323) * $signed(input_fmap_72[15:0]) +
	( 16'sd 28870) * $signed(input_fmap_73[15:0]) +
	( 15'sd 14711) * $signed(input_fmap_74[15:0]) +
	( 16'sd 19439) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19435) * $signed(input_fmap_76[15:0]) +
	( 15'sd 10577) * $signed(input_fmap_77[15:0]) +
	( 13'sd 3184) * $signed(input_fmap_78[15:0]) +
	( 16'sd 29192) * $signed(input_fmap_79[15:0]) +
	( 15'sd 8741) * $signed(input_fmap_80[15:0]) +
	( 16'sd 25929) * $signed(input_fmap_81[15:0]) +
	( 15'sd 11190) * $signed(input_fmap_82[15:0]) +
	( 16'sd 27577) * $signed(input_fmap_83[15:0]) +
	( 16'sd 16416) * $signed(input_fmap_84[15:0]) +
	( 12'sd 1076) * $signed(input_fmap_85[15:0]) +
	( 16'sd 19149) * $signed(input_fmap_86[15:0]) +
	( 16'sd 27328) * $signed(input_fmap_87[15:0]) +
	( 16'sd 31865) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5119) * $signed(input_fmap_89[15:0]) +
	( 16'sd 29966) * $signed(input_fmap_90[15:0]) +
	( 14'sd 6603) * $signed(input_fmap_91[15:0]) +
	( 15'sd 8280) * $signed(input_fmap_92[15:0]) +
	( 16'sd 28032) * $signed(input_fmap_93[15:0]) +
	( 14'sd 4287) * $signed(input_fmap_94[15:0]) +
	( 15'sd 16276) * $signed(input_fmap_95[15:0]) +
	( 16'sd 27881) * $signed(input_fmap_96[15:0]) +
	( 16'sd 19369) * $signed(input_fmap_97[15:0]) +
	( 16'sd 27245) * $signed(input_fmap_98[15:0]) +
	( 16'sd 18512) * $signed(input_fmap_99[15:0]) +
	( 15'sd 11148) * $signed(input_fmap_100[15:0]) +
	( 16'sd 25195) * $signed(input_fmap_101[15:0]) +
	( 15'sd 9010) * $signed(input_fmap_102[15:0]) +
	( 16'sd 19408) * $signed(input_fmap_103[15:0]) +
	( 15'sd 14367) * $signed(input_fmap_104[15:0]) +
	( 15'sd 15519) * $signed(input_fmap_105[15:0]) +
	( 14'sd 5634) * $signed(input_fmap_106[15:0]) +
	( 14'sd 7781) * $signed(input_fmap_107[15:0]) +
	( 16'sd 24657) * $signed(input_fmap_108[15:0]) +
	( 16'sd 21017) * $signed(input_fmap_109[15:0]) +
	( 13'sd 3953) * $signed(input_fmap_110[15:0]) +
	( 16'sd 31530) * $signed(input_fmap_111[15:0]) +
	( 14'sd 4380) * $signed(input_fmap_112[15:0]) +
	( 12'sd 1983) * $signed(input_fmap_113[15:0]) +
	( 16'sd 20223) * $signed(input_fmap_114[15:0]) +
	( 12'sd 1502) * $signed(input_fmap_115[15:0]) +
	( 16'sd 19209) * $signed(input_fmap_116[15:0]) +
	( 16'sd 25112) * $signed(input_fmap_117[15:0]) +
	( 11'sd 796) * $signed(input_fmap_118[15:0]) +
	( 15'sd 15555) * $signed(input_fmap_119[15:0]) +
	( 16'sd 31500) * $signed(input_fmap_120[15:0]) +
	( 16'sd 17390) * $signed(input_fmap_121[15:0]) +
	( 16'sd 25474) * $signed(input_fmap_122[15:0]) +
	( 15'sd 13844) * $signed(input_fmap_123[15:0]) +
	( 16'sd 22080) * $signed(input_fmap_124[15:0]) +
	( 16'sd 20837) * $signed(input_fmap_125[15:0]) +
	( 16'sd 18168) * $signed(input_fmap_126[15:0]) +
	( 16'sd 28479) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 16'sd 30045) * $signed(input_fmap_0[15:0]) +
	( 16'sd 26066) * $signed(input_fmap_1[15:0]) +
	( 14'sd 4504) * $signed(input_fmap_2[15:0]) +
	( 14'sd 5262) * $signed(input_fmap_3[15:0]) +
	( 13'sd 2633) * $signed(input_fmap_4[15:0]) +
	( 16'sd 24628) * $signed(input_fmap_5[15:0]) +
	( 14'sd 4673) * $signed(input_fmap_6[15:0]) +
	( 13'sd 2071) * $signed(input_fmap_7[15:0]) +
	( 16'sd 17112) * $signed(input_fmap_8[15:0]) +
	( 15'sd 11290) * $signed(input_fmap_9[15:0]) +
	( 16'sd 21554) * $signed(input_fmap_10[15:0]) +
	( 16'sd 29420) * $signed(input_fmap_11[15:0]) +
	( 10'sd 353) * $signed(input_fmap_12[15:0]) +
	( 16'sd 18596) * $signed(input_fmap_13[15:0]) +
	( 16'sd 24629) * $signed(input_fmap_14[15:0]) +
	( 16'sd 26135) * $signed(input_fmap_15[15:0]) +
	( 14'sd 4907) * $signed(input_fmap_16[15:0]) +
	( 15'sd 10925) * $signed(input_fmap_17[15:0]) +
	( 16'sd 24383) * $signed(input_fmap_18[15:0]) +
	( 14'sd 5225) * $signed(input_fmap_19[15:0]) +
	( 16'sd 31626) * $signed(input_fmap_20[15:0]) +
	( 16'sd 17251) * $signed(input_fmap_21[15:0]) +
	( 15'sd 8991) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24690) * $signed(input_fmap_23[15:0]) +
	( 14'sd 5611) * $signed(input_fmap_24[15:0]) +
	( 10'sd 407) * $signed(input_fmap_25[15:0]) +
	( 15'sd 13908) * $signed(input_fmap_26[15:0]) +
	( 14'sd 4461) * $signed(input_fmap_27[15:0]) +
	( 16'sd 23433) * $signed(input_fmap_28[15:0]) +
	( 14'sd 5555) * $signed(input_fmap_29[15:0]) +
	( 14'sd 5836) * $signed(input_fmap_30[15:0]) +
	( 16'sd 28698) * $signed(input_fmap_31[15:0]) +
	( 13'sd 2643) * $signed(input_fmap_32[15:0]) +
	( 16'sd 17139) * $signed(input_fmap_33[15:0]) +
	( 16'sd 28469) * $signed(input_fmap_34[15:0]) +
	( 13'sd 2332) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2804) * $signed(input_fmap_36[15:0]) +
	( 15'sd 9105) * $signed(input_fmap_37[15:0]) +
	( 14'sd 6932) * $signed(input_fmap_38[15:0]) +
	( 16'sd 17892) * $signed(input_fmap_39[15:0]) +
	( 15'sd 10485) * $signed(input_fmap_40[15:0]) +
	( 16'sd 27024) * $signed(input_fmap_41[15:0]) +
	( 16'sd 26137) * $signed(input_fmap_42[15:0]) +
	( 16'sd 24050) * $signed(input_fmap_43[15:0]) +
	( 15'sd 15424) * $signed(input_fmap_44[15:0]) +
	( 16'sd 24165) * $signed(input_fmap_45[15:0]) +
	( 14'sd 4703) * $signed(input_fmap_46[15:0]) +
	( 15'sd 10606) * $signed(input_fmap_47[15:0]) +
	( 15'sd 8600) * $signed(input_fmap_48[15:0]) +
	( 16'sd 28786) * $signed(input_fmap_49[15:0]) +
	( 14'sd 6584) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15531) * $signed(input_fmap_51[15:0]) +
	( 13'sd 3944) * $signed(input_fmap_52[15:0]) +
	( 15'sd 12687) * $signed(input_fmap_53[15:0]) +
	( 16'sd 29005) * $signed(input_fmap_54[15:0]) +
	( 15'sd 13603) * $signed(input_fmap_55[15:0]) +
	( 16'sd 32400) * $signed(input_fmap_56[15:0]) +
	( 14'sd 7849) * $signed(input_fmap_57[15:0]) +
	( 16'sd 28357) * $signed(input_fmap_58[15:0]) +
	( 15'sd 12699) * $signed(input_fmap_59[15:0]) +
	( 16'sd 18072) * $signed(input_fmap_60[15:0]) +
	( 13'sd 2825) * $signed(input_fmap_61[15:0]) +
	( 15'sd 11943) * $signed(input_fmap_62[15:0]) +
	( 16'sd 26305) * $signed(input_fmap_63[15:0]) +
	( 16'sd 20048) * $signed(input_fmap_64[15:0]) +
	( 16'sd 23263) * $signed(input_fmap_65[15:0]) +
	( 16'sd 22348) * $signed(input_fmap_66[15:0]) +
	( 15'sd 15330) * $signed(input_fmap_67[15:0]) +
	( 15'sd 10792) * $signed(input_fmap_68[15:0]) +
	( 15'sd 11881) * $signed(input_fmap_69[15:0]) +
	( 10'sd 472) * $signed(input_fmap_70[15:0]) +
	( 16'sd 19488) * $signed(input_fmap_71[15:0]) +
	( 14'sd 4463) * $signed(input_fmap_72[15:0]) +
	( 16'sd 31484) * $signed(input_fmap_73[15:0]) +
	( 16'sd 21670) * $signed(input_fmap_74[15:0]) +
	( 16'sd 28767) * $signed(input_fmap_75[15:0]) +
	( 16'sd 17655) * $signed(input_fmap_76[15:0]) +
	( 10'sd 492) * $signed(input_fmap_77[15:0]) +
	( 14'sd 7571) * $signed(input_fmap_78[15:0]) +
	( 15'sd 14496) * $signed(input_fmap_79[15:0]) +
	( 15'sd 12557) * $signed(input_fmap_80[15:0]) +
	( 14'sd 6427) * $signed(input_fmap_81[15:0]) +
	( 14'sd 5096) * $signed(input_fmap_82[15:0]) +
	( 14'sd 4241) * $signed(input_fmap_83[15:0]) +
	( 16'sd 18319) * $signed(input_fmap_84[15:0]) +
	( 16'sd 19230) * $signed(input_fmap_85[15:0]) +
	( 15'sd 10894) * $signed(input_fmap_86[15:0]) +
	( 14'sd 6697) * $signed(input_fmap_87[15:0]) +
	( 15'sd 13951) * $signed(input_fmap_88[15:0]) +
	( 16'sd 19632) * $signed(input_fmap_89[15:0]) +
	( 12'sd 1648) * $signed(input_fmap_90[15:0]) +
	( 14'sd 6251) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25756) * $signed(input_fmap_92[15:0]) +
	( 12'sd 1500) * $signed(input_fmap_93[15:0]) +
	( 15'sd 12362) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25834) * $signed(input_fmap_95[15:0]) +
	( 15'sd 16374) * $signed(input_fmap_96[15:0]) +
	( 14'sd 5360) * $signed(input_fmap_97[15:0]) +
	( 16'sd 19283) * $signed(input_fmap_98[15:0]) +
	( 15'sd 10162) * $signed(input_fmap_99[15:0]) +
	( 14'sd 4139) * $signed(input_fmap_100[15:0]) +
	( 14'sd 7536) * $signed(input_fmap_101[15:0]) +
	( 16'sd 25261) * $signed(input_fmap_102[15:0]) +
	( 16'sd 29150) * $signed(input_fmap_103[15:0]) +
	( 14'sd 5260) * $signed(input_fmap_104[15:0]) +
	( 13'sd 3294) * $signed(input_fmap_105[15:0]) +
	( 15'sd 8438) * $signed(input_fmap_106[15:0]) +
	( 16'sd 31791) * $signed(input_fmap_107[15:0]) +
	( 16'sd 26263) * $signed(input_fmap_108[15:0]) +
	( 16'sd 27382) * $signed(input_fmap_109[15:0]) +
	( 16'sd 25640) * $signed(input_fmap_110[15:0]) +
	( 16'sd 25521) * $signed(input_fmap_111[15:0]) +
	( 16'sd 16885) * $signed(input_fmap_112[15:0]) +
	( 15'sd 9950) * $signed(input_fmap_113[15:0]) +
	( 16'sd 24222) * $signed(input_fmap_114[15:0]) +
	( 14'sd 5985) * $signed(input_fmap_115[15:0]) +
	( 16'sd 16476) * $signed(input_fmap_116[15:0]) +
	( 14'sd 8022) * $signed(input_fmap_117[15:0]) +
	( 14'sd 6828) * $signed(input_fmap_118[15:0]) +
	( 16'sd 26076) * $signed(input_fmap_119[15:0]) +
	( 14'sd 5191) * $signed(input_fmap_120[15:0]) +
	( 16'sd 29372) * $signed(input_fmap_121[15:0]) +
	( 16'sd 30553) * $signed(input_fmap_122[15:0]) +
	( 15'sd 13300) * $signed(input_fmap_123[15:0]) +
	( 15'sd 10290) * $signed(input_fmap_124[15:0]) +
	( 16'sd 18024) * $signed(input_fmap_125[15:0]) +
	( 16'sd 20466) * $signed(input_fmap_126[15:0]) +
	( 16'sd 22886) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 14'sd 4761) * $signed(input_fmap_0[15:0]) +
	( 15'sd 16197) * $signed(input_fmap_1[15:0]) +
	( 15'sd 10201) * $signed(input_fmap_2[15:0]) +
	( 13'sd 2428) * $signed(input_fmap_3[15:0]) +
	( 14'sd 7708) * $signed(input_fmap_4[15:0]) +
	( 15'sd 14969) * $signed(input_fmap_5[15:0]) +
	( 16'sd 23093) * $signed(input_fmap_6[15:0]) +
	( 16'sd 17501) * $signed(input_fmap_7[15:0]) +
	( 16'sd 32592) * $signed(input_fmap_8[15:0]) +
	( 16'sd 22933) * $signed(input_fmap_9[15:0]) +
	( 16'sd 24074) * $signed(input_fmap_10[15:0]) +
	( 15'sd 13820) * $signed(input_fmap_11[15:0]) +
	( 14'sd 7771) * $signed(input_fmap_12[15:0]) +
	( 16'sd 31071) * $signed(input_fmap_13[15:0]) +
	( 16'sd 30065) * $signed(input_fmap_14[15:0]) +
	( 16'sd 26583) * $signed(input_fmap_15[15:0]) +
	( 14'sd 5689) * $signed(input_fmap_16[15:0]) +
	( 16'sd 32466) * $signed(input_fmap_17[15:0]) +
	( 16'sd 17042) * $signed(input_fmap_18[15:0]) +
	( 16'sd 19626) * $signed(input_fmap_19[15:0]) +
	( 16'sd 22937) * $signed(input_fmap_20[15:0]) +
	( 15'sd 13587) * $signed(input_fmap_21[15:0]) +
	( 16'sd 25795) * $signed(input_fmap_22[15:0]) +
	( 16'sd 32488) * $signed(input_fmap_23[15:0]) +
	( 16'sd 19510) * $signed(input_fmap_24[15:0]) +
	( 16'sd 23051) * $signed(input_fmap_25[15:0]) +
	( 16'sd 22582) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1633) * $signed(input_fmap_27[15:0]) +
	( 12'sd 1530) * $signed(input_fmap_28[15:0]) +
	( 15'sd 10235) * $signed(input_fmap_29[15:0]) +
	( 12'sd 1219) * $signed(input_fmap_30[15:0]) +
	( 15'sd 14037) * $signed(input_fmap_31[15:0]) +
	( 16'sd 17597) * $signed(input_fmap_32[15:0]) +
	( 16'sd 31149) * $signed(input_fmap_33[15:0]) +
	( 15'sd 10852) * $signed(input_fmap_34[15:0]) +
	( 16'sd 23852) * $signed(input_fmap_35[15:0]) +
	( 14'sd 6891) * $signed(input_fmap_36[15:0]) +
	( 14'sd 8098) * $signed(input_fmap_37[15:0]) +
	( 16'sd 18269) * $signed(input_fmap_38[15:0]) +
	( 14'sd 6921) * $signed(input_fmap_39[15:0]) +
	( 16'sd 21063) * $signed(input_fmap_40[15:0]) +
	( 15'sd 14193) * $signed(input_fmap_41[15:0]) +
	( 16'sd 28934) * $signed(input_fmap_42[15:0]) +
	( 16'sd 27410) * $signed(input_fmap_43[15:0]) +
	( 16'sd 31412) * $signed(input_fmap_44[15:0]) +
	( 13'sd 3757) * $signed(input_fmap_45[15:0]) +
	( 16'sd 24578) * $signed(input_fmap_46[15:0]) +
	( 16'sd 26498) * $signed(input_fmap_47[15:0]) +
	( 16'sd 25466) * $signed(input_fmap_48[15:0]) +
	( 16'sd 30076) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26327) * $signed(input_fmap_50[15:0]) +
	( 16'sd 30706) * $signed(input_fmap_51[15:0]) +
	( 16'sd 29598) * $signed(input_fmap_52[15:0]) +
	( 14'sd 5745) * $signed(input_fmap_53[15:0]) +
	( 14'sd 7959) * $signed(input_fmap_54[15:0]) +
	( 14'sd 5619) * $signed(input_fmap_55[15:0]) +
	( 16'sd 17348) * $signed(input_fmap_56[15:0]) +
	( 16'sd 25947) * $signed(input_fmap_57[15:0]) +
	( 16'sd 30186) * $signed(input_fmap_58[15:0]) +
	( 16'sd 28168) * $signed(input_fmap_59[15:0]) +
	( 16'sd 25132) * $signed(input_fmap_60[15:0]) +
	( 13'sd 2659) * $signed(input_fmap_61[15:0]) +
	( 15'sd 16108) * $signed(input_fmap_62[15:0]) +
	( 16'sd 29198) * $signed(input_fmap_63[15:0]) +
	( 15'sd 15513) * $signed(input_fmap_64[15:0]) +
	( 16'sd 26314) * $signed(input_fmap_65[15:0]) +
	( 15'sd 13777) * $signed(input_fmap_66[15:0]) +
	( 16'sd 31375) * $signed(input_fmap_67[15:0]) +
	( 14'sd 5746) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31283) * $signed(input_fmap_69[15:0]) +
	( 15'sd 13956) * $signed(input_fmap_70[15:0]) +
	( 13'sd 2364) * $signed(input_fmap_71[15:0]) +
	( 16'sd 19291) * $signed(input_fmap_72[15:0]) +
	( 15'sd 8815) * $signed(input_fmap_73[15:0]) +
	( 16'sd 26311) * $signed(input_fmap_74[15:0]) +
	( 13'sd 3206) * $signed(input_fmap_75[15:0]) +
	( 16'sd 23433) * $signed(input_fmap_76[15:0]) +
	( 16'sd 25087) * $signed(input_fmap_77[15:0]) +
	( 16'sd 32132) * $signed(input_fmap_78[15:0]) +
	( 16'sd 26810) * $signed(input_fmap_79[15:0]) +
	( 13'sd 3767) * $signed(input_fmap_80[15:0]) +
	( 16'sd 26017) * $signed(input_fmap_81[15:0]) +
	( 14'sd 7115) * $signed(input_fmap_82[15:0]) +
	( 15'sd 13739) * $signed(input_fmap_83[15:0]) +
	( 14'sd 4922) * $signed(input_fmap_84[15:0]) +
	( 13'sd 4068) * $signed(input_fmap_85[15:0]) +
	( 16'sd 17583) * $signed(input_fmap_86[15:0]) +
	( 16'sd 16508) * $signed(input_fmap_87[15:0]) +
	( 16'sd 19018) * $signed(input_fmap_88[15:0]) +
	( 15'sd 14063) * $signed(input_fmap_89[15:0]) +
	( 9'sd 191) * $signed(input_fmap_90[15:0]) +
	( 16'sd 18191) * $signed(input_fmap_91[15:0]) +
	( 16'sd 29469) * $signed(input_fmap_92[15:0]) +
	( 15'sd 16047) * $signed(input_fmap_93[15:0]) +
	( 16'sd 26565) * $signed(input_fmap_94[15:0]) +
	( 13'sd 3346) * $signed(input_fmap_95[15:0]) +
	( 15'sd 11652) * $signed(input_fmap_96[15:0]) +
	( 16'sd 23606) * $signed(input_fmap_97[15:0]) +
	( 16'sd 31420) * $signed(input_fmap_98[15:0]) +
	( 13'sd 2989) * $signed(input_fmap_99[15:0]) +
	( 16'sd 20641) * $signed(input_fmap_100[15:0]) +
	( 16'sd 31669) * $signed(input_fmap_101[15:0]) +
	( 16'sd 27755) * $signed(input_fmap_102[15:0]) +
	( 15'sd 9810) * $signed(input_fmap_103[15:0]) +
	( 10'sd 427) * $signed(input_fmap_104[15:0]) +
	( 14'sd 5513) * $signed(input_fmap_105[15:0]) +
	( 16'sd 27123) * $signed(input_fmap_106[15:0]) +
	( 13'sd 3757) * $signed(input_fmap_107[15:0]) +
	( 16'sd 17166) * $signed(input_fmap_108[15:0]) +
	( 16'sd 28974) * $signed(input_fmap_109[15:0]) +
	( 16'sd 20470) * $signed(input_fmap_110[15:0]) +
	( 14'sd 6956) * $signed(input_fmap_111[15:0]) +
	( 16'sd 17645) * $signed(input_fmap_112[15:0]) +
	( 16'sd 20302) * $signed(input_fmap_113[15:0]) +
	( 15'sd 11153) * $signed(input_fmap_114[15:0]) +
	( 12'sd 1633) * $signed(input_fmap_115[15:0]) +
	( 16'sd 32421) * $signed(input_fmap_116[15:0]) +
	( 16'sd 19552) * $signed(input_fmap_117[15:0]) +
	( 14'sd 7935) * $signed(input_fmap_118[15:0]) +
	( 14'sd 8150) * $signed(input_fmap_119[15:0]) +
	( 16'sd 29062) * $signed(input_fmap_120[15:0]) +
	( 16'sd 20635) * $signed(input_fmap_121[15:0]) +
	( 11'sd 720) * $signed(input_fmap_122[15:0]) +
	( 11'sd 629) * $signed(input_fmap_123[15:0]) +
	( 16'sd 26048) * $signed(input_fmap_124[15:0]) +
	( 12'sd 1966) * $signed(input_fmap_125[15:0]) +
	( 14'sd 5974) * $signed(input_fmap_126[15:0]) +
	( 16'sd 28504) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 16'sd 21434) * $signed(input_fmap_0[15:0]) +
	( 16'sd 21279) * $signed(input_fmap_1[15:0]) +
	( 16'sd 31030) * $signed(input_fmap_2[15:0]) +
	( 16'sd 31091) * $signed(input_fmap_3[15:0]) +
	( 15'sd 15183) * $signed(input_fmap_4[15:0]) +
	( 14'sd 4303) * $signed(input_fmap_5[15:0]) +
	( 16'sd 27158) * $signed(input_fmap_6[15:0]) +
	( 15'sd 15321) * $signed(input_fmap_7[15:0]) +
	( 16'sd 22597) * $signed(input_fmap_8[15:0]) +
	( 15'sd 11883) * $signed(input_fmap_9[15:0]) +
	( 16'sd 27992) * $signed(input_fmap_10[15:0]) +
	( 15'sd 12813) * $signed(input_fmap_11[15:0]) +
	( 15'sd 13200) * $signed(input_fmap_12[15:0]) +
	( 16'sd 27080) * $signed(input_fmap_13[15:0]) +
	( 15'sd 14805) * $signed(input_fmap_14[15:0]) +
	( 14'sd 6713) * $signed(input_fmap_15[15:0]) +
	( 13'sd 2781) * $signed(input_fmap_16[15:0]) +
	( 16'sd 27034) * $signed(input_fmap_17[15:0]) +
	( 16'sd 22821) * $signed(input_fmap_18[15:0]) +
	( 15'sd 9526) * $signed(input_fmap_19[15:0]) +
	( 15'sd 10060) * $signed(input_fmap_20[15:0]) +
	( 8'sd 115) * $signed(input_fmap_21[15:0]) +
	( 13'sd 3312) * $signed(input_fmap_22[15:0]) +
	( 15'sd 12363) * $signed(input_fmap_23[15:0]) +
	( 15'sd 14843) * $signed(input_fmap_24[15:0]) +
	( 13'sd 2685) * $signed(input_fmap_25[15:0]) +
	( 16'sd 32228) * $signed(input_fmap_26[15:0]) +
	( 14'sd 5770) * $signed(input_fmap_27[15:0]) +
	( 16'sd 17105) * $signed(input_fmap_28[15:0]) +
	( 16'sd 23798) * $signed(input_fmap_29[15:0]) +
	( 16'sd 31874) * $signed(input_fmap_30[15:0]) +
	( 16'sd 29666) * $signed(input_fmap_31[15:0]) +
	( 14'sd 5389) * $signed(input_fmap_32[15:0]) +
	( 16'sd 22508) * $signed(input_fmap_33[15:0]) +
	( 15'sd 14472) * $signed(input_fmap_34[15:0]) +
	( 16'sd 16939) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2307) * $signed(input_fmap_36[15:0]) +
	( 16'sd 21622) * $signed(input_fmap_37[15:0]) +
	( 13'sd 3215) * $signed(input_fmap_38[15:0]) +
	( 16'sd 23994) * $signed(input_fmap_39[15:0]) +
	( 14'sd 5078) * $signed(input_fmap_40[15:0]) +
	( 13'sd 3405) * $signed(input_fmap_41[15:0]) +
	( 16'sd 31907) * $signed(input_fmap_42[15:0]) +
	( 16'sd 20352) * $signed(input_fmap_43[15:0]) +
	( 13'sd 2878) * $signed(input_fmap_44[15:0]) +
	( 14'sd 6786) * $signed(input_fmap_45[15:0]) +
	( 13'sd 2400) * $signed(input_fmap_46[15:0]) +
	( 16'sd 21153) * $signed(input_fmap_47[15:0]) +
	( 16'sd 21255) * $signed(input_fmap_48[15:0]) +
	( 16'sd 24241) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22552) * $signed(input_fmap_50[15:0]) +
	( 16'sd 21933) * $signed(input_fmap_51[15:0]) +
	( 15'sd 13233) * $signed(input_fmap_52[15:0]) +
	( 16'sd 28662) * $signed(input_fmap_53[15:0]) +
	( 16'sd 19411) * $signed(input_fmap_54[15:0]) +
	( 16'sd 18258) * $signed(input_fmap_55[15:0]) +
	( 14'sd 5511) * $signed(input_fmap_56[15:0]) +
	( 16'sd 19937) * $signed(input_fmap_57[15:0]) +
	( 16'sd 19655) * $signed(input_fmap_58[15:0]) +
	( 16'sd 25738) * $signed(input_fmap_59[15:0]) +
	( 13'sd 2601) * $signed(input_fmap_60[15:0]) +
	( 16'sd 32595) * $signed(input_fmap_61[15:0]) +
	( 16'sd 27349) * $signed(input_fmap_62[15:0]) +
	( 16'sd 17416) * $signed(input_fmap_63[15:0]) +
	( 15'sd 11885) * $signed(input_fmap_64[15:0]) +
	( 16'sd 32272) * $signed(input_fmap_65[15:0]) +
	( 16'sd 25480) * $signed(input_fmap_66[15:0]) +
	( 11'sd 560) * $signed(input_fmap_67[15:0]) +
	( 14'sd 4911) * $signed(input_fmap_68[15:0]) +
	( 16'sd 19825) * $signed(input_fmap_69[15:0]) +
	( 15'sd 8583) * $signed(input_fmap_70[15:0]) +
	( 16'sd 23601) * $signed(input_fmap_71[15:0]) +
	( 13'sd 4081) * $signed(input_fmap_72[15:0]) +
	( 16'sd 26594) * $signed(input_fmap_73[15:0]) +
	( 16'sd 16572) * $signed(input_fmap_74[15:0]) +
	( 14'sd 5679) * $signed(input_fmap_75[15:0]) +
	( 16'sd 28820) * $signed(input_fmap_76[15:0]) +
	( 15'sd 9500) * $signed(input_fmap_77[15:0]) +
	( 16'sd 27766) * $signed(input_fmap_78[15:0]) +
	( 16'sd 20086) * $signed(input_fmap_79[15:0]) +
	( 16'sd 30220) * $signed(input_fmap_80[15:0]) +
	( 16'sd 17736) * $signed(input_fmap_81[15:0]) +
	( 16'sd 25056) * $signed(input_fmap_82[15:0]) +
	( 16'sd 28086) * $signed(input_fmap_83[15:0]) +
	( 15'sd 14562) * $signed(input_fmap_84[15:0]) +
	( 13'sd 3189) * $signed(input_fmap_85[15:0]) +
	( 13'sd 3635) * $signed(input_fmap_86[15:0]) +
	( 15'sd 13861) * $signed(input_fmap_87[15:0]) +
	( 16'sd 29917) * $signed(input_fmap_88[15:0]) +
	( 16'sd 21105) * $signed(input_fmap_89[15:0]) +
	( 14'sd 5634) * $signed(input_fmap_90[15:0]) +
	( 15'sd 14820) * $signed(input_fmap_91[15:0]) +
	( 16'sd 21294) * $signed(input_fmap_92[15:0]) +
	( 16'sd 27867) * $signed(input_fmap_93[15:0]) +
	( 15'sd 13826) * $signed(input_fmap_94[15:0]) +
	( 15'sd 15204) * $signed(input_fmap_95[15:0]) +
	( 15'sd 15581) * $signed(input_fmap_96[15:0]) +
	( 15'sd 9076) * $signed(input_fmap_97[15:0]) +
	( 16'sd 23764) * $signed(input_fmap_98[15:0]) +
	( 15'sd 13021) * $signed(input_fmap_99[15:0]) +
	( 16'sd 25845) * $signed(input_fmap_100[15:0]) +
	( 15'sd 14140) * $signed(input_fmap_101[15:0]) +
	( 16'sd 22182) * $signed(input_fmap_102[15:0]) +
	( 14'sd 6691) * $signed(input_fmap_103[15:0]) +
	( 16'sd 17837) * $signed(input_fmap_104[15:0]) +
	( 13'sd 3230) * $signed(input_fmap_105[15:0]) +
	( 16'sd 32735) * $signed(input_fmap_106[15:0]) +
	( 13'sd 3606) * $signed(input_fmap_107[15:0]) +
	( 15'sd 9540) * $signed(input_fmap_108[15:0]) +
	( 15'sd 13411) * $signed(input_fmap_109[15:0]) +
	( 16'sd 19724) * $signed(input_fmap_110[15:0]) +
	( 14'sd 4799) * $signed(input_fmap_111[15:0]) +
	( 15'sd 13206) * $signed(input_fmap_112[15:0]) +
	( 15'sd 15199) * $signed(input_fmap_113[15:0]) +
	( 15'sd 9308) * $signed(input_fmap_114[15:0]) +
	( 16'sd 23858) * $signed(input_fmap_115[15:0]) +
	( 15'sd 11338) * $signed(input_fmap_116[15:0]) +
	( 12'sd 1972) * $signed(input_fmap_117[15:0]) +
	( 16'sd 18918) * $signed(input_fmap_118[15:0]) +
	( 14'sd 4706) * $signed(input_fmap_119[15:0]) +
	( 16'sd 22122) * $signed(input_fmap_120[15:0]) +
	( 16'sd 24665) * $signed(input_fmap_121[15:0]) +
	( 16'sd 20342) * $signed(input_fmap_122[15:0]) +
	( 16'sd 28963) * $signed(input_fmap_123[15:0]) +
	( 16'sd 28130) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24596) * $signed(input_fmap_125[15:0]) +
	( 16'sd 24810) * $signed(input_fmap_126[15:0]) +
	( 16'sd 31545) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 13'sd 2401) * $signed(input_fmap_0[15:0]) +
	( 16'sd 21437) * $signed(input_fmap_1[15:0]) +
	( 15'sd 13446) * $signed(input_fmap_2[15:0]) +
	( 15'sd 10978) * $signed(input_fmap_3[15:0]) +
	( 16'sd 21632) * $signed(input_fmap_4[15:0]) +
	( 16'sd 27070) * $signed(input_fmap_5[15:0]) +
	( 15'sd 13911) * $signed(input_fmap_6[15:0]) +
	( 16'sd 23459) * $signed(input_fmap_7[15:0]) +
	( 15'sd 8218) * $signed(input_fmap_8[15:0]) +
	( 16'sd 27995) * $signed(input_fmap_9[15:0]) +
	( 16'sd 27533) * $signed(input_fmap_10[15:0]) +
	( 16'sd 23873) * $signed(input_fmap_11[15:0]) +
	( 16'sd 28425) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24517) * $signed(input_fmap_13[15:0]) +
	( 10'sd 495) * $signed(input_fmap_14[15:0]) +
	( 14'sd 6923) * $signed(input_fmap_15[15:0]) +
	( 16'sd 21692) * $signed(input_fmap_16[15:0]) +
	( 16'sd 25117) * $signed(input_fmap_17[15:0]) +
	( 16'sd 21841) * $signed(input_fmap_18[15:0]) +
	( 16'sd 29573) * $signed(input_fmap_19[15:0]) +
	( 15'sd 16221) * $signed(input_fmap_20[15:0]) +
	( 15'sd 10051) * $signed(input_fmap_21[15:0]) +
	( 15'sd 12873) * $signed(input_fmap_22[15:0]) +
	( 15'sd 12915) * $signed(input_fmap_23[15:0]) +
	( 13'sd 3793) * $signed(input_fmap_24[15:0]) +
	( 16'sd 21496) * $signed(input_fmap_25[15:0]) +
	( 15'sd 12357) * $signed(input_fmap_26[15:0]) +
	( 16'sd 26545) * $signed(input_fmap_27[15:0]) +
	( 16'sd 32374) * $signed(input_fmap_28[15:0]) +
	( 15'sd 15356) * $signed(input_fmap_29[15:0]) +
	( 15'sd 15638) * $signed(input_fmap_30[15:0]) +
	( 16'sd 31343) * $signed(input_fmap_31[15:0]) +
	( 16'sd 22138) * $signed(input_fmap_32[15:0]) +
	( 16'sd 18023) * $signed(input_fmap_33[15:0]) +
	( 15'sd 12425) * $signed(input_fmap_34[15:0]) +
	( 15'sd 8683) * $signed(input_fmap_35[15:0]) +
	( 16'sd 29151) * $signed(input_fmap_36[15:0]) +
	( 16'sd 26282) * $signed(input_fmap_37[15:0]) +
	( 16'sd 26692) * $signed(input_fmap_38[15:0]) +
	( 14'sd 7916) * $signed(input_fmap_39[15:0]) +
	( 15'sd 12723) * $signed(input_fmap_40[15:0]) +
	( 10'sd 333) * $signed(input_fmap_41[15:0]) +
	( 15'sd 14781) * $signed(input_fmap_42[15:0]) +
	( 13'sd 2382) * $signed(input_fmap_43[15:0]) +
	( 16'sd 24024) * $signed(input_fmap_44[15:0]) +
	( 15'sd 15105) * $signed(input_fmap_45[15:0]) +
	( 16'sd 21627) * $signed(input_fmap_46[15:0]) +
	( 12'sd 1119) * $signed(input_fmap_47[15:0]) +
	( 15'sd 15889) * $signed(input_fmap_48[15:0]) +
	( 16'sd 19130) * $signed(input_fmap_49[15:0]) +
	( 15'sd 10850) * $signed(input_fmap_50[15:0]) +
	( 15'sd 8887) * $signed(input_fmap_51[15:0]) +
	( 16'sd 28810) * $signed(input_fmap_52[15:0]) +
	( 14'sd 6395) * $signed(input_fmap_53[15:0]) +
	( 15'sd 8845) * $signed(input_fmap_54[15:0]) +
	( 16'sd 26584) * $signed(input_fmap_55[15:0]) +
	( 13'sd 3256) * $signed(input_fmap_56[15:0]) +
	( 15'sd 10699) * $signed(input_fmap_57[15:0]) +
	( 16'sd 29879) * $signed(input_fmap_58[15:0]) +
	( 14'sd 6826) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1975) * $signed(input_fmap_60[15:0]) +
	( 13'sd 2885) * $signed(input_fmap_61[15:0]) +
	( 16'sd 32598) * $signed(input_fmap_62[15:0]) +
	( 16'sd 28010) * $signed(input_fmap_63[15:0]) +
	( 16'sd 19378) * $signed(input_fmap_64[15:0]) +
	( 16'sd 25553) * $signed(input_fmap_65[15:0]) +
	( 16'sd 28687) * $signed(input_fmap_66[15:0]) +
	( 13'sd 3659) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26258) * $signed(input_fmap_68[15:0]) +
	( 16'sd 23205) * $signed(input_fmap_69[15:0]) +
	( 16'sd 26483) * $signed(input_fmap_70[15:0]) +
	( 13'sd 3032) * $signed(input_fmap_71[15:0]) +
	( 13'sd 2708) * $signed(input_fmap_72[15:0]) +
	( 16'sd 28130) * $signed(input_fmap_73[15:0]) +
	( 14'sd 5716) * $signed(input_fmap_74[15:0]) +
	( 14'sd 4889) * $signed(input_fmap_75[15:0]) +
	( 15'sd 15201) * $signed(input_fmap_76[15:0]) +
	( 16'sd 24317) * $signed(input_fmap_77[15:0]) +
	( 14'sd 5050) * $signed(input_fmap_78[15:0]) +
	( 16'sd 30597) * $signed(input_fmap_79[15:0]) +
	( 4'sd 4) * $signed(input_fmap_80[15:0]) +
	( 16'sd 32415) * $signed(input_fmap_81[15:0]) +
	( 15'sd 13580) * $signed(input_fmap_82[15:0]) +
	( 16'sd 24305) * $signed(input_fmap_83[15:0]) +
	( 16'sd 28626) * $signed(input_fmap_84[15:0]) +
	( 14'sd 5017) * $signed(input_fmap_85[15:0]) +
	( 16'sd 18321) * $signed(input_fmap_86[15:0]) +
	( 14'sd 8136) * $signed(input_fmap_87[15:0]) +
	( 14'sd 5822) * $signed(input_fmap_88[15:0]) +
	( 16'sd 32347) * $signed(input_fmap_89[15:0]) +
	( 16'sd 18312) * $signed(input_fmap_90[15:0]) +
	( 16'sd 19856) * $signed(input_fmap_91[15:0]) +
	( 11'sd 934) * $signed(input_fmap_92[15:0]) +
	( 16'sd 20854) * $signed(input_fmap_93[15:0]) +
	( 13'sd 2241) * $signed(input_fmap_94[15:0]) +
	( 14'sd 4803) * $signed(input_fmap_95[15:0]) +
	( 13'sd 2734) * $signed(input_fmap_96[15:0]) +
	( 12'sd 1303) * $signed(input_fmap_97[15:0]) +
	( 16'sd 20764) * $signed(input_fmap_98[15:0]) +
	( 16'sd 29820) * $signed(input_fmap_99[15:0]) +
	( 16'sd 17082) * $signed(input_fmap_100[15:0]) +
	( 16'sd 17456) * $signed(input_fmap_101[15:0]) +
	( 15'sd 8983) * $signed(input_fmap_102[15:0]) +
	( 16'sd 26123) * $signed(input_fmap_103[15:0]) +
	( 16'sd 28141) * $signed(input_fmap_104[15:0]) +
	( 15'sd 8705) * $signed(input_fmap_105[15:0]) +
	( 16'sd 29310) * $signed(input_fmap_106[15:0]) +
	( 16'sd 22279) * $signed(input_fmap_107[15:0]) +
	( 16'sd 18992) * $signed(input_fmap_108[15:0]) +
	( 13'sd 3043) * $signed(input_fmap_109[15:0]) +
	( 16'sd 26060) * $signed(input_fmap_110[15:0]) +
	( 12'sd 1641) * $signed(input_fmap_111[15:0]) +
	( 15'sd 13453) * $signed(input_fmap_112[15:0]) +
	( 16'sd 27290) * $signed(input_fmap_113[15:0]) +
	( 16'sd 18432) * $signed(input_fmap_114[15:0]) +
	( 16'sd 20469) * $signed(input_fmap_115[15:0]) +
	( 14'sd 7357) * $signed(input_fmap_116[15:0]) +
	( 16'sd 31864) * $signed(input_fmap_117[15:0]) +
	( 16'sd 18197) * $signed(input_fmap_118[15:0]) +
	( 16'sd 16883) * $signed(input_fmap_119[15:0]) +
	( 15'sd 8221) * $signed(input_fmap_120[15:0]) +
	( 15'sd 15481) * $signed(input_fmap_121[15:0]) +
	( 12'sd 1997) * $signed(input_fmap_122[15:0]) +
	( 16'sd 18531) * $signed(input_fmap_123[15:0]) +
	( 16'sd 24788) * $signed(input_fmap_124[15:0]) +
	( 16'sd 21810) * $signed(input_fmap_125[15:0]) +
	( 16'sd 24530) * $signed(input_fmap_126[15:0]) +
	( 15'sd 8249) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 16'sd 21207) * $signed(input_fmap_0[15:0]) +
	( 10'sd 349) * $signed(input_fmap_1[15:0]) +
	( 16'sd 17752) * $signed(input_fmap_2[15:0]) +
	( 16'sd 22739) * $signed(input_fmap_3[15:0]) +
	( 15'sd 11938) * $signed(input_fmap_4[15:0]) +
	( 15'sd 9035) * $signed(input_fmap_5[15:0]) +
	( 15'sd 9307) * $signed(input_fmap_6[15:0]) +
	( 16'sd 27037) * $signed(input_fmap_7[15:0]) +
	( 16'sd 21205) * $signed(input_fmap_8[15:0]) +
	( 15'sd 12887) * $signed(input_fmap_9[15:0]) +
	( 16'sd 28741) * $signed(input_fmap_10[15:0]) +
	( 14'sd 4790) * $signed(input_fmap_11[15:0]) +
	( 14'sd 4727) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24756) * $signed(input_fmap_13[15:0]) +
	( 15'sd 15891) * $signed(input_fmap_14[15:0]) +
	( 15'sd 15642) * $signed(input_fmap_15[15:0]) +
	( 16'sd 23395) * $signed(input_fmap_16[15:0]) +
	( 16'sd 28463) * $signed(input_fmap_17[15:0]) +
	( 15'sd 15843) * $signed(input_fmap_18[15:0]) +
	( 16'sd 22975) * $signed(input_fmap_19[15:0]) +
	( 11'sd 747) * $signed(input_fmap_20[15:0]) +
	( 14'sd 7067) * $signed(input_fmap_21[15:0]) +
	( 15'sd 13653) * $signed(input_fmap_22[15:0]) +
	( 15'sd 14299) * $signed(input_fmap_23[15:0]) +
	( 16'sd 30585) * $signed(input_fmap_24[15:0]) +
	( 15'sd 9424) * $signed(input_fmap_25[15:0]) +
	( 16'sd 26346) * $signed(input_fmap_26[15:0]) +
	( 15'sd 13593) * $signed(input_fmap_27[15:0]) +
	( 15'sd 8979) * $signed(input_fmap_28[15:0]) +
	( 14'sd 6495) * $signed(input_fmap_29[15:0]) +
	( 16'sd 31218) * $signed(input_fmap_30[15:0]) +
	( 15'sd 12869) * $signed(input_fmap_31[15:0]) +
	( 16'sd 32189) * $signed(input_fmap_32[15:0]) +
	( 16'sd 21611) * $signed(input_fmap_33[15:0]) +
	( 14'sd 6839) * $signed(input_fmap_34[15:0]) +
	( 15'sd 9835) * $signed(input_fmap_35[15:0]) +
	( 16'sd 19765) * $signed(input_fmap_36[15:0]) +
	( 16'sd 25428) * $signed(input_fmap_37[15:0]) +
	( 16'sd 23869) * $signed(input_fmap_38[15:0]) +
	( 13'sd 2216) * $signed(input_fmap_39[15:0]) +
	( 15'sd 11720) * $signed(input_fmap_40[15:0]) +
	( 16'sd 21134) * $signed(input_fmap_41[15:0]) +
	( 16'sd 22166) * $signed(input_fmap_42[15:0]) +
	( 14'sd 7816) * $signed(input_fmap_43[15:0]) +
	( 13'sd 2601) * $signed(input_fmap_44[15:0]) +
	( 16'sd 28961) * $signed(input_fmap_45[15:0]) +
	( 15'sd 10943) * $signed(input_fmap_46[15:0]) +
	( 14'sd 4953) * $signed(input_fmap_47[15:0]) +
	( 16'sd 24638) * $signed(input_fmap_48[15:0]) +
	( 12'sd 1045) * $signed(input_fmap_49[15:0]) +
	( 15'sd 15067) * $signed(input_fmap_50[15:0]) +
	( 16'sd 20872) * $signed(input_fmap_51[15:0]) +
	( 16'sd 22276) * $signed(input_fmap_52[15:0]) +
	( 15'sd 12358) * $signed(input_fmap_53[15:0]) +
	( 16'sd 29095) * $signed(input_fmap_54[15:0]) +
	( 16'sd 29024) * $signed(input_fmap_55[15:0]) +
	( 15'sd 10237) * $signed(input_fmap_56[15:0]) +
	( 16'sd 29270) * $signed(input_fmap_57[15:0]) +
	( 14'sd 7956) * $signed(input_fmap_58[15:0]) +
	( 16'sd 31200) * $signed(input_fmap_59[15:0]) +
	( 16'sd 27892) * $signed(input_fmap_60[15:0]) +
	( 14'sd 5371) * $signed(input_fmap_61[15:0]) +
	( 15'sd 12506) * $signed(input_fmap_62[15:0]) +
	( 16'sd 23054) * $signed(input_fmap_63[15:0]) +
	( 15'sd 11705) * $signed(input_fmap_64[15:0]) +
	( 14'sd 5021) * $signed(input_fmap_65[15:0]) +
	( 16'sd 26304) * $signed(input_fmap_66[15:0]) +
	( 16'sd 29491) * $signed(input_fmap_67[15:0]) +
	( 14'sd 7098) * $signed(input_fmap_68[15:0]) +
	( 15'sd 8461) * $signed(input_fmap_69[15:0]) +
	( 16'sd 17425) * $signed(input_fmap_70[15:0]) +
	( 16'sd 17470) * $signed(input_fmap_71[15:0]) +
	( 15'sd 9183) * $signed(input_fmap_72[15:0]) +
	( 15'sd 15980) * $signed(input_fmap_73[15:0]) +
	( 16'sd 23740) * $signed(input_fmap_74[15:0]) +
	( 16'sd 25390) * $signed(input_fmap_75[15:0]) +
	( 15'sd 13516) * $signed(input_fmap_76[15:0]) +
	( 16'sd 26894) * $signed(input_fmap_77[15:0]) +
	( 16'sd 26663) * $signed(input_fmap_78[15:0]) +
	( 16'sd 19582) * $signed(input_fmap_79[15:0]) +
	( 16'sd 17791) * $signed(input_fmap_80[15:0]) +
	( 15'sd 8539) * $signed(input_fmap_81[15:0]) +
	( 16'sd 19791) * $signed(input_fmap_82[15:0]) +
	( 16'sd 24202) * $signed(input_fmap_83[15:0]) +
	( 14'sd 7018) * $signed(input_fmap_84[15:0]) +
	( 14'sd 6034) * $signed(input_fmap_85[15:0]) +
	( 12'sd 1976) * $signed(input_fmap_86[15:0]) +
	( 13'sd 3357) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6490) * $signed(input_fmap_88[15:0]) +
	( 15'sd 9745) * $signed(input_fmap_89[15:0]) +
	( 15'sd 12637) * $signed(input_fmap_90[15:0]) +
	( 14'sd 5243) * $signed(input_fmap_91[15:0]) +
	( 15'sd 13890) * $signed(input_fmap_92[15:0]) +
	( 15'sd 10255) * $signed(input_fmap_93[15:0]) +
	( 16'sd 29770) * $signed(input_fmap_94[15:0]) +
	( 15'sd 15987) * $signed(input_fmap_95[15:0]) +
	( 11'sd 938) * $signed(input_fmap_96[15:0]) +
	( 9'sd 145) * $signed(input_fmap_97[15:0]) +
	( 16'sd 20899) * $signed(input_fmap_98[15:0]) +
	( 16'sd 19314) * $signed(input_fmap_99[15:0]) +
	( 16'sd 21454) * $signed(input_fmap_100[15:0]) +
	( 15'sd 15313) * $signed(input_fmap_101[15:0]) +
	( 14'sd 6621) * $signed(input_fmap_102[15:0]) +
	( 16'sd 18426) * $signed(input_fmap_103[15:0]) +
	( 13'sd 2679) * $signed(input_fmap_104[15:0]) +
	( 15'sd 15501) * $signed(input_fmap_105[15:0]) +
	( 14'sd 7569) * $signed(input_fmap_106[15:0]) +
	( 15'sd 11808) * $signed(input_fmap_107[15:0]) +
	( 13'sd 2329) * $signed(input_fmap_108[15:0]) +
	( 16'sd 32375) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22628) * $signed(input_fmap_110[15:0]) +
	( 15'sd 8555) * $signed(input_fmap_111[15:0]) +
	( 15'sd 15760) * $signed(input_fmap_112[15:0]) +
	( 16'sd 23513) * $signed(input_fmap_113[15:0]) +
	( 14'sd 5260) * $signed(input_fmap_114[15:0]) +
	( 13'sd 2673) * $signed(input_fmap_115[15:0]) +
	( 16'sd 30164) * $signed(input_fmap_116[15:0]) +
	( 16'sd 31056) * $signed(input_fmap_117[15:0]) +
	( 16'sd 21356) * $signed(input_fmap_118[15:0]) +
	( 16'sd 17874) * $signed(input_fmap_119[15:0]) +
	( 16'sd 27122) * $signed(input_fmap_120[15:0]) +
	( 16'sd 16791) * $signed(input_fmap_121[15:0]) +
	( 13'sd 2460) * $signed(input_fmap_122[15:0]) +
	( 16'sd 32278) * $signed(input_fmap_123[15:0]) +
	( 15'sd 10283) * $signed(input_fmap_124[15:0]) +
	( 13'sd 2469) * $signed(input_fmap_125[15:0]) +
	( 15'sd 9907) * $signed(input_fmap_126[15:0]) +
	( 16'sd 22218) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 14'sd 7803) * $signed(input_fmap_0[15:0]) +
	( 15'sd 10517) * $signed(input_fmap_1[15:0]) +
	( 16'sd 21127) * $signed(input_fmap_2[15:0]) +
	( 16'sd 23918) * $signed(input_fmap_3[15:0]) +
	( 16'sd 16876) * $signed(input_fmap_4[15:0]) +
	( 14'sd 5725) * $signed(input_fmap_5[15:0]) +
	( 16'sd 26026) * $signed(input_fmap_6[15:0]) +
	( 15'sd 15718) * $signed(input_fmap_7[15:0]) +
	( 14'sd 4717) * $signed(input_fmap_8[15:0]) +
	( 16'sd 24102) * $signed(input_fmap_9[15:0]) +
	( 16'sd 19000) * $signed(input_fmap_10[15:0]) +
	( 16'sd 26280) * $signed(input_fmap_11[15:0]) +
	( 16'sd 24557) * $signed(input_fmap_12[15:0]) +
	( 15'sd 11799) * $signed(input_fmap_13[15:0]) +
	( 14'sd 5054) * $signed(input_fmap_14[15:0]) +
	( 16'sd 31146) * $signed(input_fmap_15[15:0]) +
	( 15'sd 15460) * $signed(input_fmap_16[15:0]) +
	( 16'sd 17135) * $signed(input_fmap_17[15:0]) +
	( 15'sd 14313) * $signed(input_fmap_18[15:0]) +
	( 13'sd 2998) * $signed(input_fmap_19[15:0]) +
	( 16'sd 29694) * $signed(input_fmap_20[15:0]) +
	( 16'sd 26150) * $signed(input_fmap_21[15:0]) +
	( 16'sd 25351) * $signed(input_fmap_22[15:0]) +
	( 16'sd 26840) * $signed(input_fmap_23[15:0]) +
	( 16'sd 31730) * $signed(input_fmap_24[15:0]) +
	( 14'sd 7480) * $signed(input_fmap_25[15:0]) +
	( 14'sd 6909) * $signed(input_fmap_26[15:0]) +
	( 14'sd 6847) * $signed(input_fmap_27[15:0]) +
	( 14'sd 4158) * $signed(input_fmap_28[15:0]) +
	( 15'sd 12117) * $signed(input_fmap_29[15:0]) +
	( 16'sd 18305) * $signed(input_fmap_30[15:0]) +
	( 15'sd 13082) * $signed(input_fmap_31[15:0]) +
	( 16'sd 20104) * $signed(input_fmap_32[15:0]) +
	( 14'sd 6653) * $signed(input_fmap_33[15:0]) +
	( 16'sd 18617) * $signed(input_fmap_34[15:0]) +
	( 16'sd 22507) * $signed(input_fmap_35[15:0]) +
	( 15'sd 13788) * $signed(input_fmap_36[15:0]) +
	( 16'sd 25679) * $signed(input_fmap_37[15:0]) +
	( 15'sd 11904) * $signed(input_fmap_38[15:0]) +
	( 16'sd 17397) * $signed(input_fmap_39[15:0]) +
	( 16'sd 29315) * $signed(input_fmap_40[15:0]) +
	( 15'sd 10679) * $signed(input_fmap_41[15:0]) +
	( 11'sd 719) * $signed(input_fmap_42[15:0]) +
	( 15'sd 9485) * $signed(input_fmap_43[15:0]) +
	( 14'sd 4438) * $signed(input_fmap_44[15:0]) +
	( 15'sd 9564) * $signed(input_fmap_45[15:0]) +
	( 16'sd 21542) * $signed(input_fmap_46[15:0]) +
	( 15'sd 11332) * $signed(input_fmap_47[15:0]) +
	( 16'sd 27604) * $signed(input_fmap_48[15:0]) +
	( 14'sd 7799) * $signed(input_fmap_49[15:0]) +
	( 14'sd 5514) * $signed(input_fmap_50[15:0]) +
	( 15'sd 14378) * $signed(input_fmap_51[15:0]) +
	( 14'sd 8031) * $signed(input_fmap_52[15:0]) +
	( 14'sd 5109) * $signed(input_fmap_53[15:0]) +
	( 16'sd 22124) * $signed(input_fmap_54[15:0]) +
	( 16'sd 19779) * $signed(input_fmap_55[15:0]) +
	( 12'sd 1792) * $signed(input_fmap_56[15:0]) +
	( 15'sd 12569) * $signed(input_fmap_57[15:0]) +
	( 16'sd 32468) * $signed(input_fmap_58[15:0]) +
	( 14'sd 4348) * $signed(input_fmap_59[15:0]) +
	( 16'sd 21352) * $signed(input_fmap_60[15:0]) +
	( 15'sd 12699) * $signed(input_fmap_61[15:0]) +
	( 12'sd 1492) * $signed(input_fmap_62[15:0]) +
	( 16'sd 19467) * $signed(input_fmap_63[15:0]) +
	( 15'sd 14052) * $signed(input_fmap_64[15:0]) +
	( 16'sd 22873) * $signed(input_fmap_65[15:0]) +
	( 14'sd 4735) * $signed(input_fmap_66[15:0]) +
	( 15'sd 12701) * $signed(input_fmap_67[15:0]) +
	( 16'sd 21600) * $signed(input_fmap_68[15:0]) +
	( 13'sd 3447) * $signed(input_fmap_69[15:0]) +
	( 14'sd 8068) * $signed(input_fmap_70[15:0]) +
	( 14'sd 5205) * $signed(input_fmap_71[15:0]) +
	( 16'sd 24743) * $signed(input_fmap_72[15:0]) +
	( 15'sd 9732) * $signed(input_fmap_73[15:0]) +
	( 13'sd 3465) * $signed(input_fmap_74[15:0]) +
	( 16'sd 26308) * $signed(input_fmap_75[15:0]) +
	( 16'sd 21269) * $signed(input_fmap_76[15:0]) +
	( 12'sd 1424) * $signed(input_fmap_77[15:0]) +
	( 16'sd 20165) * $signed(input_fmap_78[15:0]) +
	( 16'sd 23738) * $signed(input_fmap_79[15:0]) +
	( 13'sd 3382) * $signed(input_fmap_80[15:0]) +
	( 16'sd 20198) * $signed(input_fmap_81[15:0]) +
	( 14'sd 7906) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25050) * $signed(input_fmap_83[15:0]) +
	( 13'sd 2353) * $signed(input_fmap_84[15:0]) +
	( 12'sd 1183) * $signed(input_fmap_85[15:0]) +
	( 15'sd 13965) * $signed(input_fmap_86[15:0]) +
	( 16'sd 27329) * $signed(input_fmap_87[15:0]) +
	( 16'sd 21053) * $signed(input_fmap_88[15:0]) +
	( 13'sd 4029) * $signed(input_fmap_89[15:0]) +
	( 16'sd 20614) * $signed(input_fmap_90[15:0]) +
	( 12'sd 1710) * $signed(input_fmap_91[15:0]) +
	( 16'sd 22877) * $signed(input_fmap_92[15:0]) +
	( 15'sd 10592) * $signed(input_fmap_93[15:0]) +
	( 14'sd 6192) * $signed(input_fmap_94[15:0]) +
	( 16'sd 21195) * $signed(input_fmap_95[15:0]) +
	( 16'sd 18786) * $signed(input_fmap_96[15:0]) +
	( 15'sd 9168) * $signed(input_fmap_97[15:0]) +
	( 16'sd 24558) * $signed(input_fmap_98[15:0]) +
	( 12'sd 1792) * $signed(input_fmap_99[15:0]) +
	( 15'sd 13881) * $signed(input_fmap_100[15:0]) +
	( 16'sd 29061) * $signed(input_fmap_101[15:0]) +
	( 16'sd 25371) * $signed(input_fmap_102[15:0]) +
	( 15'sd 14181) * $signed(input_fmap_103[15:0]) +
	( 16'sd 26042) * $signed(input_fmap_104[15:0]) +
	( 16'sd 20221) * $signed(input_fmap_105[15:0]) +
	( 12'sd 1648) * $signed(input_fmap_106[15:0]) +
	( 16'sd 22538) * $signed(input_fmap_107[15:0]) +
	( 16'sd 30105) * $signed(input_fmap_108[15:0]) +
	( 16'sd 17361) * $signed(input_fmap_109[15:0]) +
	( 16'sd 19982) * $signed(input_fmap_110[15:0]) +
	( 15'sd 12123) * $signed(input_fmap_111[15:0]) +
	( 16'sd 24710) * $signed(input_fmap_112[15:0]) +
	( 15'sd 8314) * $signed(input_fmap_113[15:0]) +
	( 13'sd 3295) * $signed(input_fmap_114[15:0]) +
	( 16'sd 26685) * $signed(input_fmap_115[15:0]) +
	( 16'sd 27278) * $signed(input_fmap_116[15:0]) +
	( 15'sd 12852) * $signed(input_fmap_117[15:0]) +
	( 8'sd 103) * $signed(input_fmap_118[15:0]) +
	( 16'sd 21534) * $signed(input_fmap_119[15:0]) +
	( 15'sd 13876) * $signed(input_fmap_120[15:0]) +
	( 13'sd 3749) * $signed(input_fmap_121[15:0]) +
	( 12'sd 1471) * $signed(input_fmap_122[15:0]) +
	( 16'sd 32381) * $signed(input_fmap_123[15:0]) +
	( 13'sd 2750) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24645) * $signed(input_fmap_125[15:0]) +
	( 16'sd 17545) * $signed(input_fmap_126[15:0]) +
	( 14'sd 8000) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 16'sd 24805) * $signed(input_fmap_0[15:0]) +
	( 14'sd 4699) * $signed(input_fmap_1[15:0]) +
	( 16'sd 24134) * $signed(input_fmap_2[15:0]) +
	( 16'sd 32738) * $signed(input_fmap_3[15:0]) +
	( 16'sd 27661) * $signed(input_fmap_4[15:0]) +
	( 16'sd 26615) * $signed(input_fmap_5[15:0]) +
	( 16'sd 30012) * $signed(input_fmap_6[15:0]) +
	( 14'sd 6964) * $signed(input_fmap_7[15:0]) +
	( 14'sd 7121) * $signed(input_fmap_8[15:0]) +
	( 16'sd 18840) * $signed(input_fmap_9[15:0]) +
	( 16'sd 29142) * $signed(input_fmap_10[15:0]) +
	( 16'sd 23465) * $signed(input_fmap_11[15:0]) +
	( 16'sd 20016) * $signed(input_fmap_12[15:0]) +
	( 14'sd 7631) * $signed(input_fmap_13[15:0]) +
	( 14'sd 6584) * $signed(input_fmap_14[15:0]) +
	( 14'sd 5028) * $signed(input_fmap_15[15:0]) +
	( 14'sd 8095) * $signed(input_fmap_16[15:0]) +
	( 15'sd 11436) * $signed(input_fmap_17[15:0]) +
	( 15'sd 10300) * $signed(input_fmap_18[15:0]) +
	( 16'sd 24664) * $signed(input_fmap_19[15:0]) +
	( 16'sd 29996) * $signed(input_fmap_20[15:0]) +
	( 16'sd 25526) * $signed(input_fmap_21[15:0]) +
	( 14'sd 6527) * $signed(input_fmap_22[15:0]) +
	( 16'sd 28776) * $signed(input_fmap_23[15:0]) +
	( 16'sd 29558) * $signed(input_fmap_24[15:0]) +
	( 16'sd 27604) * $signed(input_fmap_25[15:0]) +
	( 14'sd 4522) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2068) * $signed(input_fmap_27[15:0]) +
	( 15'sd 12112) * $signed(input_fmap_28[15:0]) +
	( 15'sd 10034) * $signed(input_fmap_29[15:0]) +
	( 11'sd 817) * $signed(input_fmap_30[15:0]) +
	( 14'sd 7875) * $signed(input_fmap_31[15:0]) +
	( 14'sd 6167) * $signed(input_fmap_32[15:0]) +
	( 14'sd 4142) * $signed(input_fmap_33[15:0]) +
	( 12'sd 1686) * $signed(input_fmap_34[15:0]) +
	( 15'sd 11963) * $signed(input_fmap_35[15:0]) +
	( 16'sd 27741) * $signed(input_fmap_36[15:0]) +
	( 14'sd 6316) * $signed(input_fmap_37[15:0]) +
	( 16'sd 27370) * $signed(input_fmap_38[15:0]) +
	( 16'sd 25209) * $signed(input_fmap_39[15:0]) +
	( 14'sd 7251) * $signed(input_fmap_40[15:0]) +
	( 16'sd 22470) * $signed(input_fmap_41[15:0]) +
	( 13'sd 3808) * $signed(input_fmap_42[15:0]) +
	( 14'sd 7193) * $signed(input_fmap_43[15:0]) +
	( 15'sd 12345) * $signed(input_fmap_44[15:0]) +
	( 16'sd 31493) * $signed(input_fmap_45[15:0]) +
	( 16'sd 27357) * $signed(input_fmap_46[15:0]) +
	( 16'sd 28530) * $signed(input_fmap_47[15:0]) +
	( 15'sd 14416) * $signed(input_fmap_48[15:0]) +
	( 16'sd 28016) * $signed(input_fmap_49[15:0]) +
	( 16'sd 16392) * $signed(input_fmap_50[15:0]) +
	( 15'sd 14934) * $signed(input_fmap_51[15:0]) +
	( 16'sd 21518) * $signed(input_fmap_52[15:0]) +
	( 13'sd 3143) * $signed(input_fmap_53[15:0]) +
	( 15'sd 13171) * $signed(input_fmap_54[15:0]) +
	( 16'sd 30792) * $signed(input_fmap_55[15:0]) +
	( 14'sd 7824) * $signed(input_fmap_56[15:0]) +
	( 16'sd 32274) * $signed(input_fmap_57[15:0]) +
	( 15'sd 15023) * $signed(input_fmap_58[15:0]) +
	( 13'sd 3217) * $signed(input_fmap_59[15:0]) +
	( 14'sd 7050) * $signed(input_fmap_60[15:0]) +
	( 14'sd 5218) * $signed(input_fmap_61[15:0]) +
	( 16'sd 28885) * $signed(input_fmap_62[15:0]) +
	( 16'sd 32492) * $signed(input_fmap_63[15:0]) +
	( 16'sd 21799) * $signed(input_fmap_64[15:0]) +
	( 16'sd 19275) * $signed(input_fmap_65[15:0]) +
	( 16'sd 19368) * $signed(input_fmap_66[15:0]) +
	( 14'sd 5237) * $signed(input_fmap_67[15:0]) +
	( 16'sd 31650) * $signed(input_fmap_68[15:0]) +
	( 14'sd 6964) * $signed(input_fmap_69[15:0]) +
	( 16'sd 25729) * $signed(input_fmap_70[15:0]) +
	( 16'sd 23490) * $signed(input_fmap_71[15:0]) +
	( 15'sd 9768) * $signed(input_fmap_72[15:0]) +
	( 16'sd 31093) * $signed(input_fmap_73[15:0]) +
	( 15'sd 11538) * $signed(input_fmap_74[15:0]) +
	( 16'sd 30793) * $signed(input_fmap_75[15:0]) +
	( 15'sd 9272) * $signed(input_fmap_76[15:0]) +
	( 15'sd 12429) * $signed(input_fmap_77[15:0]) +
	( 13'sd 3141) * $signed(input_fmap_78[15:0]) +
	( 15'sd 14518) * $signed(input_fmap_79[15:0]) +
	( 16'sd 26942) * $signed(input_fmap_80[15:0]) +
	( 14'sd 6075) * $signed(input_fmap_81[15:0]) +
	( 15'sd 9829) * $signed(input_fmap_82[15:0]) +
	( 16'sd 28441) * $signed(input_fmap_83[15:0]) +
	( 15'sd 10402) * $signed(input_fmap_84[15:0]) +
	( 13'sd 2183) * $signed(input_fmap_85[15:0]) +
	( 15'sd 11911) * $signed(input_fmap_86[15:0]) +
	( 15'sd 8512) * $signed(input_fmap_87[15:0]) +
	( 16'sd 26956) * $signed(input_fmap_88[15:0]) +
	( 14'sd 4234) * $signed(input_fmap_89[15:0]) +
	( 16'sd 20435) * $signed(input_fmap_90[15:0]) +
	( 16'sd 22603) * $signed(input_fmap_91[15:0]) +
	( 10'sd 281) * $signed(input_fmap_92[15:0]) +
	( 12'sd 1807) * $signed(input_fmap_93[15:0]) +
	( 16'sd 26771) * $signed(input_fmap_94[15:0]) +
	( 16'sd 21650) * $signed(input_fmap_95[15:0]) +
	( 16'sd 23035) * $signed(input_fmap_96[15:0]) +
	( 14'sd 5551) * $signed(input_fmap_97[15:0]) +
	( 8'sd 103) * $signed(input_fmap_98[15:0]) +
	( 16'sd 18484) * $signed(input_fmap_99[15:0]) +
	( 16'sd 20098) * $signed(input_fmap_100[15:0]) +
	( 16'sd 27390) * $signed(input_fmap_101[15:0]) +
	( 16'sd 28538) * $signed(input_fmap_102[15:0]) +
	( 14'sd 5241) * $signed(input_fmap_103[15:0]) +
	( 16'sd 32650) * $signed(input_fmap_104[15:0]) +
	( 16'sd 31897) * $signed(input_fmap_105[15:0]) +
	( 16'sd 24251) * $signed(input_fmap_106[15:0]) +
	( 14'sd 7086) * $signed(input_fmap_107[15:0]) +
	( 14'sd 6330) * $signed(input_fmap_108[15:0]) +
	( 15'sd 16336) * $signed(input_fmap_109[15:0]) +
	( 16'sd 23349) * $signed(input_fmap_110[15:0]) +
	( 16'sd 27927) * $signed(input_fmap_111[15:0]) +
	( 15'sd 10812) * $signed(input_fmap_112[15:0]) +
	( 14'sd 5229) * $signed(input_fmap_113[15:0]) +
	( 15'sd 10333) * $signed(input_fmap_114[15:0]) +
	( 15'sd 16229) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15152) * $signed(input_fmap_116[15:0]) +
	( 13'sd 2234) * $signed(input_fmap_117[15:0]) +
	( 6'sd 16) * $signed(input_fmap_118[15:0]) +
	( 14'sd 4703) * $signed(input_fmap_119[15:0]) +
	( 16'sd 24291) * $signed(input_fmap_120[15:0]) +
	( 15'sd 13872) * $signed(input_fmap_121[15:0]) +
	( 15'sd 14665) * $signed(input_fmap_122[15:0]) +
	( 11'sd 973) * $signed(input_fmap_123[15:0]) +
	( 15'sd 13329) * $signed(input_fmap_124[15:0]) +
	( 16'sd 18599) * $signed(input_fmap_125[15:0]) +
	( 16'sd 32386) * $signed(input_fmap_126[15:0]) +
	( 16'sd 32121) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 16'sd 26528) * $signed(input_fmap_0[15:0]) +
	( 13'sd 3406) * $signed(input_fmap_1[15:0]) +
	( 16'sd 26541) * $signed(input_fmap_2[15:0]) +
	( 7'sd 45) * $signed(input_fmap_3[15:0]) +
	( 16'sd 18652) * $signed(input_fmap_4[15:0]) +
	( 14'sd 4779) * $signed(input_fmap_5[15:0]) +
	( 16'sd 16458) * $signed(input_fmap_6[15:0]) +
	( 16'sd 23490) * $signed(input_fmap_7[15:0]) +
	( 15'sd 12512) * $signed(input_fmap_8[15:0]) +
	( 16'sd 29653) * $signed(input_fmap_9[15:0]) +
	( 15'sd 13957) * $signed(input_fmap_10[15:0]) +
	( 16'sd 18650) * $signed(input_fmap_11[15:0]) +
	( 16'sd 25861) * $signed(input_fmap_12[15:0]) +
	( 16'sd 22494) * $signed(input_fmap_13[15:0]) +
	( 16'sd 23630) * $signed(input_fmap_14[15:0]) +
	( 6'sd 22) * $signed(input_fmap_15[15:0]) +
	( 13'sd 3391) * $signed(input_fmap_16[15:0]) +
	( 16'sd 24904) * $signed(input_fmap_17[15:0]) +
	( 15'sd 10103) * $signed(input_fmap_18[15:0]) +
	( 16'sd 27052) * $signed(input_fmap_19[15:0]) +
	( 12'sd 1883) * $signed(input_fmap_20[15:0]) +
	( 16'sd 30599) * $signed(input_fmap_21[15:0]) +
	( 16'sd 32764) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24526) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17562) * $signed(input_fmap_24[15:0]) +
	( 16'sd 23763) * $signed(input_fmap_25[15:0]) +
	( 16'sd 17218) * $signed(input_fmap_26[15:0]) +
	( 15'sd 8724) * $signed(input_fmap_27[15:0]) +
	( 15'sd 12149) * $signed(input_fmap_28[15:0]) +
	( 14'sd 8015) * $signed(input_fmap_29[15:0]) +
	( 16'sd 29500) * $signed(input_fmap_30[15:0]) +
	( 16'sd 22389) * $signed(input_fmap_31[15:0]) +
	( 16'sd 26436) * $signed(input_fmap_32[15:0]) +
	( 14'sd 5687) * $signed(input_fmap_33[15:0]) +
	( 15'sd 9773) * $signed(input_fmap_34[15:0]) +
	( 15'sd 10573) * $signed(input_fmap_35[15:0]) +
	( 14'sd 7613) * $signed(input_fmap_36[15:0]) +
	( 11'sd 694) * $signed(input_fmap_37[15:0]) +
	( 14'sd 7204) * $signed(input_fmap_38[15:0]) +
	( 15'sd 15741) * $signed(input_fmap_39[15:0]) +
	( 16'sd 30945) * $signed(input_fmap_40[15:0]) +
	( 15'sd 14227) * $signed(input_fmap_41[15:0]) +
	( 15'sd 15921) * $signed(input_fmap_42[15:0]) +
	( 16'sd 22155) * $signed(input_fmap_43[15:0]) +
	( 16'sd 18324) * $signed(input_fmap_44[15:0]) +
	( 6'sd 19) * $signed(input_fmap_45[15:0]) +
	( 11'sd 882) * $signed(input_fmap_46[15:0]) +
	( 16'sd 24571) * $signed(input_fmap_47[15:0]) +
	( 16'sd 25654) * $signed(input_fmap_48[15:0]) +
	( 15'sd 10848) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26611) * $signed(input_fmap_50[15:0]) +
	( 8'sd 104) * $signed(input_fmap_51[15:0]) +
	( 16'sd 29087) * $signed(input_fmap_52[15:0]) +
	( 13'sd 2711) * $signed(input_fmap_53[15:0]) +
	( 16'sd 22504) * $signed(input_fmap_54[15:0]) +
	( 16'sd 28215) * $signed(input_fmap_55[15:0]) +
	( 16'sd 27645) * $signed(input_fmap_56[15:0]) +
	( 15'sd 11518) * $signed(input_fmap_57[15:0]) +
	( 13'sd 3167) * $signed(input_fmap_58[15:0]) +
	( 15'sd 11549) * $signed(input_fmap_59[15:0]) +
	( 14'sd 4108) * $signed(input_fmap_60[15:0]) +
	( 16'sd 22246) * $signed(input_fmap_61[15:0]) +
	( 13'sd 2355) * $signed(input_fmap_62[15:0]) +
	( 15'sd 13162) * $signed(input_fmap_63[15:0]) +
	( 16'sd 23241) * $signed(input_fmap_64[15:0]) +
	( 13'sd 3734) * $signed(input_fmap_65[15:0]) +
	( 16'sd 32626) * $signed(input_fmap_66[15:0]) +
	( 16'sd 21830) * $signed(input_fmap_67[15:0]) +
	( 15'sd 12708) * $signed(input_fmap_68[15:0]) +
	( 14'sd 6890) * $signed(input_fmap_69[15:0]) +
	( 15'sd 12714) * $signed(input_fmap_70[15:0]) +
	( 16'sd 26983) * $signed(input_fmap_71[15:0]) +
	( 15'sd 15337) * $signed(input_fmap_72[15:0]) +
	( 14'sd 5603) * $signed(input_fmap_73[15:0]) +
	( 13'sd 2259) * $signed(input_fmap_74[15:0]) +
	( 16'sd 17860) * $signed(input_fmap_75[15:0]) +
	( 16'sd 19544) * $signed(input_fmap_76[15:0]) +
	( 16'sd 19753) * $signed(input_fmap_77[15:0]) +
	( 16'sd 27460) * $signed(input_fmap_78[15:0]) +
	( 13'sd 2107) * $signed(input_fmap_79[15:0]) +
	( 15'sd 15466) * $signed(input_fmap_80[15:0]) +
	( 16'sd 31944) * $signed(input_fmap_81[15:0]) +
	( 11'sd 885) * $signed(input_fmap_82[15:0]) +
	( 15'sd 8253) * $signed(input_fmap_83[15:0]) +
	( 15'sd 12817) * $signed(input_fmap_84[15:0]) +
	( 16'sd 26140) * $signed(input_fmap_85[15:0]) +
	( 16'sd 25337) * $signed(input_fmap_86[15:0]) +
	( 15'sd 15779) * $signed(input_fmap_87[15:0]) +
	( 15'sd 11369) * $signed(input_fmap_88[15:0]) +
	( 16'sd 30034) * $signed(input_fmap_89[15:0]) +
	( 15'sd 14713) * $signed(input_fmap_90[15:0]) +
	( 15'sd 14868) * $signed(input_fmap_91[15:0]) +
	( 16'sd 25347) * $signed(input_fmap_92[15:0]) +
	( 16'sd 21663) * $signed(input_fmap_93[15:0]) +
	( 16'sd 29271) * $signed(input_fmap_94[15:0]) +
	( 16'sd 24413) * $signed(input_fmap_95[15:0]) +
	( 10'sd 294) * $signed(input_fmap_96[15:0]) +
	( 16'sd 30979) * $signed(input_fmap_97[15:0]) +
	( 16'sd 16942) * $signed(input_fmap_98[15:0]) +
	( 15'sd 13941) * $signed(input_fmap_99[15:0]) +
	( 15'sd 16231) * $signed(input_fmap_100[15:0]) +
	( 16'sd 21250) * $signed(input_fmap_101[15:0]) +
	( 15'sd 13280) * $signed(input_fmap_102[15:0]) +
	( 14'sd 4786) * $signed(input_fmap_103[15:0]) +
	( 15'sd 8399) * $signed(input_fmap_104[15:0]) +
	( 16'sd 32028) * $signed(input_fmap_105[15:0]) +
	( 16'sd 25633) * $signed(input_fmap_106[15:0]) +
	( 11'sd 664) * $signed(input_fmap_107[15:0]) +
	( 16'sd 21537) * $signed(input_fmap_108[15:0]) +
	( 16'sd 22490) * $signed(input_fmap_109[15:0]) +
	( 15'sd 9039) * $signed(input_fmap_110[15:0]) +
	( 16'sd 18661) * $signed(input_fmap_111[15:0]) +
	( 16'sd 21214) * $signed(input_fmap_112[15:0]) +
	( 16'sd 25763) * $signed(input_fmap_113[15:0]) +
	( 16'sd 19926) * $signed(input_fmap_114[15:0]) +
	( 16'sd 30279) * $signed(input_fmap_115[15:0]) +
	( 16'sd 18138) * $signed(input_fmap_116[15:0]) +
	( 13'sd 2777) * $signed(input_fmap_117[15:0]) +
	( 15'sd 9538) * $signed(input_fmap_118[15:0]) +
	( 16'sd 25861) * $signed(input_fmap_119[15:0]) +
	( 14'sd 7094) * $signed(input_fmap_120[15:0]) +
	( 16'sd 25459) * $signed(input_fmap_121[15:0]) +
	( 12'sd 1946) * $signed(input_fmap_122[15:0]) +
	( 15'sd 16304) * $signed(input_fmap_123[15:0]) +
	( 16'sd 24962) * $signed(input_fmap_124[15:0]) +
	( 15'sd 8574) * $signed(input_fmap_125[15:0]) +
	( 16'sd 26862) * $signed(input_fmap_126[15:0]) +
	( 16'sd 27181) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 15'sd 12516) * $signed(input_fmap_0[15:0]) +
	( 12'sd 1092) * $signed(input_fmap_1[15:0]) +
	( 16'sd 17307) * $signed(input_fmap_2[15:0]) +
	( 11'sd 776) * $signed(input_fmap_3[15:0]) +
	( 16'sd 25956) * $signed(input_fmap_4[15:0]) +
	( 13'sd 2745) * $signed(input_fmap_5[15:0]) +
	( 15'sd 14986) * $signed(input_fmap_6[15:0]) +
	( 16'sd 27860) * $signed(input_fmap_7[15:0]) +
	( 16'sd 19089) * $signed(input_fmap_8[15:0]) +
	( 14'sd 4229) * $signed(input_fmap_9[15:0]) +
	( 16'sd 29267) * $signed(input_fmap_10[15:0]) +
	( 14'sd 5513) * $signed(input_fmap_11[15:0]) +
	( 14'sd 5499) * $signed(input_fmap_12[15:0]) +
	( 15'sd 15356) * $signed(input_fmap_13[15:0]) +
	( 14'sd 5298) * $signed(input_fmap_14[15:0]) +
	( 16'sd 27525) * $signed(input_fmap_15[15:0]) +
	( 16'sd 31683) * $signed(input_fmap_16[15:0]) +
	( 14'sd 4176) * $signed(input_fmap_17[15:0]) +
	( 16'sd 24742) * $signed(input_fmap_18[15:0]) +
	( 16'sd 19140) * $signed(input_fmap_19[15:0]) +
	( 15'sd 8868) * $signed(input_fmap_20[15:0]) +
	( 15'sd 10339) * $signed(input_fmap_21[15:0]) +
	( 15'sd 12476) * $signed(input_fmap_22[15:0]) +
	( 16'sd 24827) * $signed(input_fmap_23[15:0]) +
	( 16'sd 32434) * $signed(input_fmap_24[15:0]) +
	( 10'sd 432) * $signed(input_fmap_25[15:0]) +
	( 12'sd 2020) * $signed(input_fmap_26[15:0]) +
	( 14'sd 6326) * $signed(input_fmap_27[15:0]) +
	( 15'sd 8698) * $signed(input_fmap_28[15:0]) +
	( 14'sd 6764) * $signed(input_fmap_29[15:0]) +
	( 11'sd 656) * $signed(input_fmap_30[15:0]) +
	( 15'sd 13941) * $signed(input_fmap_31[15:0]) +
	( 14'sd 7411) * $signed(input_fmap_32[15:0]) +
	( 15'sd 8323) * $signed(input_fmap_33[15:0]) +
	( 14'sd 5099) * $signed(input_fmap_34[15:0]) +
	( 16'sd 25147) * $signed(input_fmap_35[15:0]) +
	( 16'sd 20317) * $signed(input_fmap_36[15:0]) +
	( 15'sd 11012) * $signed(input_fmap_37[15:0]) +
	( 15'sd 11488) * $signed(input_fmap_38[15:0]) +
	( 16'sd 21102) * $signed(input_fmap_39[15:0]) +
	( 16'sd 27099) * $signed(input_fmap_40[15:0]) +
	( 9'sd 187) * $signed(input_fmap_41[15:0]) +
	( 16'sd 26125) * $signed(input_fmap_42[15:0]) +
	( 15'sd 10139) * $signed(input_fmap_43[15:0]) +
	( 16'sd 23279) * $signed(input_fmap_44[15:0]) +
	( 16'sd 22422) * $signed(input_fmap_45[15:0]) +
	( 15'sd 15081) * $signed(input_fmap_46[15:0]) +
	( 16'sd 19574) * $signed(input_fmap_47[15:0]) +
	( 14'sd 5415) * $signed(input_fmap_48[15:0]) +
	( 15'sd 10427) * $signed(input_fmap_49[15:0]) +
	( 15'sd 15445) * $signed(input_fmap_50[15:0]) +
	( 16'sd 25600) * $signed(input_fmap_51[15:0]) +
	( 15'sd 16189) * $signed(input_fmap_52[15:0]) +
	( 14'sd 6899) * $signed(input_fmap_53[15:0]) +
	( 16'sd 25312) * $signed(input_fmap_54[15:0]) +
	( 16'sd 16430) * $signed(input_fmap_55[15:0]) +
	( 15'sd 10363) * $signed(input_fmap_56[15:0]) +
	( 16'sd 19582) * $signed(input_fmap_57[15:0]) +
	( 15'sd 12126) * $signed(input_fmap_58[15:0]) +
	( 16'sd 20427) * $signed(input_fmap_59[15:0]) +
	( 16'sd 18141) * $signed(input_fmap_60[15:0]) +
	( 16'sd 27348) * $signed(input_fmap_61[15:0]) +
	( 16'sd 26277) * $signed(input_fmap_62[15:0]) +
	( 16'sd 28110) * $signed(input_fmap_63[15:0]) +
	( 12'sd 1357) * $signed(input_fmap_64[15:0]) +
	( 16'sd 22880) * $signed(input_fmap_65[15:0]) +
	( 11'sd 748) * $signed(input_fmap_66[15:0]) +
	( 15'sd 8788) * $signed(input_fmap_67[15:0]) +
	( 14'sd 4538) * $signed(input_fmap_68[15:0]) +
	( 16'sd 30923) * $signed(input_fmap_69[15:0]) +
	( 16'sd 30864) * $signed(input_fmap_70[15:0]) +
	( 16'sd 22305) * $signed(input_fmap_71[15:0]) +
	( 15'sd 14768) * $signed(input_fmap_72[15:0]) +
	( 15'sd 9393) * $signed(input_fmap_73[15:0]) +
	( 16'sd 23223) * $signed(input_fmap_74[15:0]) +
	( 16'sd 29968) * $signed(input_fmap_75[15:0]) +
	( 16'sd 31132) * $signed(input_fmap_76[15:0]) +
	( 16'sd 17533) * $signed(input_fmap_77[15:0]) +
	( 16'sd 29880) * $signed(input_fmap_78[15:0]) +
	( 16'sd 28567) * $signed(input_fmap_79[15:0]) +
	( 15'sd 13323) * $signed(input_fmap_80[15:0]) +
	( 16'sd 29493) * $signed(input_fmap_81[15:0]) +
	( 15'sd 15085) * $signed(input_fmap_82[15:0]) +
	( 16'sd 19182) * $signed(input_fmap_83[15:0]) +
	( 16'sd 24842) * $signed(input_fmap_84[15:0]) +
	( 13'sd 3796) * $signed(input_fmap_85[15:0]) +
	( 16'sd 30391) * $signed(input_fmap_86[15:0]) +
	( 15'sd 11824) * $signed(input_fmap_87[15:0]) +
	( 15'sd 11435) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5939) * $signed(input_fmap_89[15:0]) +
	( 16'sd 31384) * $signed(input_fmap_90[15:0]) +
	( 16'sd 25384) * $signed(input_fmap_91[15:0]) +
	( 16'sd 21614) * $signed(input_fmap_92[15:0]) +
	( 16'sd 20907) * $signed(input_fmap_93[15:0]) +
	( 16'sd 29439) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25385) * $signed(input_fmap_95[15:0]) +
	( 16'sd 17437) * $signed(input_fmap_96[15:0]) +
	( 16'sd 30346) * $signed(input_fmap_97[15:0]) +
	( 14'sd 8015) * $signed(input_fmap_98[15:0]) +
	( 16'sd 24757) * $signed(input_fmap_99[15:0]) +
	( 16'sd 24630) * $signed(input_fmap_100[15:0]) +
	( 16'sd 24836) * $signed(input_fmap_101[15:0]) +
	( 15'sd 10387) * $signed(input_fmap_102[15:0]) +
	( 16'sd 31173) * $signed(input_fmap_103[15:0]) +
	( 14'sd 4529) * $signed(input_fmap_104[15:0]) +
	( 16'sd 19751) * $signed(input_fmap_105[15:0]) +
	( 15'sd 8463) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27001) * $signed(input_fmap_107[15:0]) +
	( 14'sd 5049) * $signed(input_fmap_108[15:0]) +
	( 16'sd 24217) * $signed(input_fmap_109[15:0]) +
	( 15'sd 14442) * $signed(input_fmap_110[15:0]) +
	( 10'sd 352) * $signed(input_fmap_111[15:0]) +
	( 12'sd 1963) * $signed(input_fmap_112[15:0]) +
	( 15'sd 10620) * $signed(input_fmap_113[15:0]) +
	( 15'sd 9481) * $signed(input_fmap_114[15:0]) +
	( 14'sd 4339) * $signed(input_fmap_115[15:0]) +
	( 13'sd 3056) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27057) * $signed(input_fmap_117[15:0]) +
	( 15'sd 13125) * $signed(input_fmap_118[15:0]) +
	( 15'sd 11314) * $signed(input_fmap_119[15:0]) +
	( 16'sd 21345) * $signed(input_fmap_120[15:0]) +
	( 16'sd 17119) * $signed(input_fmap_121[15:0]) +
	( 15'sd 10491) * $signed(input_fmap_122[15:0]) +
	( 16'sd 22421) * $signed(input_fmap_123[15:0]) +
	( 16'sd 21642) * $signed(input_fmap_124[15:0]) +
	( 14'sd 6644) * $signed(input_fmap_125[15:0]) +
	( 15'sd 13690) * $signed(input_fmap_126[15:0]) +
	( 15'sd 11417) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 15'sd 10681) * $signed(input_fmap_0[15:0]) +
	( 14'sd 7077) * $signed(input_fmap_1[15:0]) +
	( 16'sd 29407) * $signed(input_fmap_2[15:0]) +
	( 15'sd 11848) * $signed(input_fmap_3[15:0]) +
	( 16'sd 21136) * $signed(input_fmap_4[15:0]) +
	( 15'sd 9173) * $signed(input_fmap_5[15:0]) +
	( 16'sd 22693) * $signed(input_fmap_6[15:0]) +
	( 16'sd 21494) * $signed(input_fmap_7[15:0]) +
	( 16'sd 30180) * $signed(input_fmap_8[15:0]) +
	( 15'sd 12839) * $signed(input_fmap_9[15:0]) +
	( 16'sd 22437) * $signed(input_fmap_10[15:0]) +
	( 16'sd 22444) * $signed(input_fmap_11[15:0]) +
	( 15'sd 8392) * $signed(input_fmap_12[15:0]) +
	( 16'sd 24420) * $signed(input_fmap_13[15:0]) +
	( 15'sd 11642) * $signed(input_fmap_14[15:0]) +
	( 16'sd 24237) * $signed(input_fmap_15[15:0]) +
	( 15'sd 9229) * $signed(input_fmap_16[15:0]) +
	( 16'sd 22017) * $signed(input_fmap_17[15:0]) +
	( 13'sd 3855) * $signed(input_fmap_18[15:0]) +
	( 15'sd 9716) * $signed(input_fmap_19[15:0]) +
	( 16'sd 17553) * $signed(input_fmap_20[15:0]) +
	( 16'sd 28612) * $signed(input_fmap_21[15:0]) +
	( 15'sd 15155) * $signed(input_fmap_22[15:0]) +
	( 16'sd 26022) * $signed(input_fmap_23[15:0]) +
	( 11'sd 588) * $signed(input_fmap_24[15:0]) +
	( 14'sd 6577) * $signed(input_fmap_25[15:0]) +
	( 15'sd 10882) * $signed(input_fmap_26[15:0]) +
	( 16'sd 29600) * $signed(input_fmap_27[15:0]) +
	( 16'sd 20705) * $signed(input_fmap_28[15:0]) +
	( 14'sd 4855) * $signed(input_fmap_29[15:0]) +
	( 16'sd 23912) * $signed(input_fmap_30[15:0]) +
	( 16'sd 21492) * $signed(input_fmap_31[15:0]) +
	( 15'sd 11951) * $signed(input_fmap_32[15:0]) +
	( 13'sd 3820) * $signed(input_fmap_33[15:0]) +
	( 16'sd 22639) * $signed(input_fmap_34[15:0]) +
	( 16'sd 21040) * $signed(input_fmap_35[15:0]) +
	( 14'sd 6761) * $signed(input_fmap_36[15:0]) +
	( 14'sd 5090) * $signed(input_fmap_37[15:0]) +
	( 16'sd 19398) * $signed(input_fmap_38[15:0]) +
	( 15'sd 10289) * $signed(input_fmap_39[15:0]) +
	( 13'sd 2272) * $signed(input_fmap_40[15:0]) +
	( 16'sd 23037) * $signed(input_fmap_41[15:0]) +
	( 16'sd 32602) * $signed(input_fmap_42[15:0]) +
	( 16'sd 19403) * $signed(input_fmap_43[15:0]) +
	( 15'sd 10018) * $signed(input_fmap_44[15:0]) +
	( 15'sd 9185) * $signed(input_fmap_45[15:0]) +
	( 16'sd 24063) * $signed(input_fmap_46[15:0]) +
	( 15'sd 12228) * $signed(input_fmap_47[15:0]) +
	( 16'sd 20347) * $signed(input_fmap_48[15:0]) +
	( 16'sd 23648) * $signed(input_fmap_49[15:0]) +
	( 16'sd 16930) * $signed(input_fmap_50[15:0]) +
	( 15'sd 15121) * $signed(input_fmap_51[15:0]) +
	( 16'sd 31366) * $signed(input_fmap_52[15:0]) +
	( 16'sd 27425) * $signed(input_fmap_53[15:0]) +
	( 10'sd 404) * $signed(input_fmap_54[15:0]) +
	( 16'sd 17678) * $signed(input_fmap_55[15:0]) +
	( 15'sd 9948) * $signed(input_fmap_56[15:0]) +
	( 15'sd 8315) * $signed(input_fmap_57[15:0]) +
	( 16'sd 31398) * $signed(input_fmap_58[15:0]) +
	( 12'sd 1182) * $signed(input_fmap_59[15:0]) +
	( 16'sd 29545) * $signed(input_fmap_60[15:0]) +
	( 15'sd 10092) * $signed(input_fmap_61[15:0]) +
	( 15'sd 12341) * $signed(input_fmap_62[15:0]) +
	( 15'sd 12570) * $signed(input_fmap_63[15:0]) +
	( 16'sd 25730) * $signed(input_fmap_64[15:0]) +
	( 14'sd 4338) * $signed(input_fmap_65[15:0]) +
	( 15'sd 14121) * $signed(input_fmap_66[15:0]) +
	( 16'sd 22480) * $signed(input_fmap_67[15:0]) +
	( 15'sd 14193) * $signed(input_fmap_68[15:0]) +
	( 15'sd 8744) * $signed(input_fmap_69[15:0]) +
	( 16'sd 27613) * $signed(input_fmap_70[15:0]) +
	( 14'sd 7473) * $signed(input_fmap_71[15:0]) +
	( 16'sd 16433) * $signed(input_fmap_72[15:0]) +
	( 16'sd 26932) * $signed(input_fmap_73[15:0]) +
	( 15'sd 13342) * $signed(input_fmap_74[15:0]) +
	( 15'sd 10114) * $signed(input_fmap_75[15:0]) +
	( 15'sd 11368) * $signed(input_fmap_76[15:0]) +
	( 16'sd 21572) * $signed(input_fmap_77[15:0]) +
	( 16'sd 18249) * $signed(input_fmap_78[15:0]) +
	( 16'sd 18111) * $signed(input_fmap_79[15:0]) +
	( 14'sd 6956) * $signed(input_fmap_80[15:0]) +
	( 14'sd 5403) * $signed(input_fmap_81[15:0]) +
	( 16'sd 22041) * $signed(input_fmap_82[15:0]) +
	( 15'sd 9654) * $signed(input_fmap_83[15:0]) +
	( 16'sd 18209) * $signed(input_fmap_84[15:0]) +
	( 16'sd 27150) * $signed(input_fmap_85[15:0]) +
	( 14'sd 4147) * $signed(input_fmap_86[15:0]) +
	( 15'sd 13331) * $signed(input_fmap_87[15:0]) +
	( 16'sd 23725) * $signed(input_fmap_88[15:0]) +
	( 16'sd 24211) * $signed(input_fmap_89[15:0]) +
	( 16'sd 17611) * $signed(input_fmap_90[15:0]) +
	( 16'sd 23675) * $signed(input_fmap_91[15:0]) +
	( 16'sd 21146) * $signed(input_fmap_92[15:0]) +
	( 16'sd 23547) * $signed(input_fmap_93[15:0]) +
	( 14'sd 4865) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25082) * $signed(input_fmap_95[15:0]) +
	( 13'sd 4033) * $signed(input_fmap_96[15:0]) +
	( 13'sd 3595) * $signed(input_fmap_97[15:0]) +
	( 16'sd 29516) * $signed(input_fmap_98[15:0]) +
	( 15'sd 16174) * $signed(input_fmap_99[15:0]) +
	( 16'sd 22750) * $signed(input_fmap_100[15:0]) +
	( 16'sd 21789) * $signed(input_fmap_101[15:0]) +
	( 16'sd 25880) * $signed(input_fmap_102[15:0]) +
	( 16'sd 18205) * $signed(input_fmap_103[15:0]) +
	( 14'sd 7971) * $signed(input_fmap_104[15:0]) +
	( 16'sd 29712) * $signed(input_fmap_105[15:0]) +
	( 16'sd 21649) * $signed(input_fmap_106[15:0]) +
	( 15'sd 15163) * $signed(input_fmap_107[15:0]) +
	( 15'sd 10447) * $signed(input_fmap_108[15:0]) +
	( 15'sd 10533) * $signed(input_fmap_109[15:0]) +
	( 12'sd 1933) * $signed(input_fmap_110[15:0]) +
	( 14'sd 7961) * $signed(input_fmap_111[15:0]) +
	( 15'sd 11619) * $signed(input_fmap_112[15:0]) +
	( 16'sd 25898) * $signed(input_fmap_113[15:0]) +
	( 15'sd 14147) * $signed(input_fmap_114[15:0]) +
	( 15'sd 15287) * $signed(input_fmap_115[15:0]) +
	( 16'sd 19590) * $signed(input_fmap_116[15:0]) +
	( 16'sd 25421) * $signed(input_fmap_117[15:0]) +
	( 16'sd 32120) * $signed(input_fmap_118[15:0]) +
	( 16'sd 30399) * $signed(input_fmap_119[15:0]) +
	( 16'sd 23144) * $signed(input_fmap_120[15:0]) +
	( 16'sd 24935) * $signed(input_fmap_121[15:0]) +
	( 16'sd 25163) * $signed(input_fmap_122[15:0]) +
	( 16'sd 17543) * $signed(input_fmap_123[15:0]) +
	( 16'sd 32594) * $signed(input_fmap_124[15:0]) +
	( 13'sd 3892) * $signed(input_fmap_125[15:0]) +
	( 16'sd 27076) * $signed(input_fmap_126[15:0]) +
	( 15'sd 12799) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 14'sd 4696) * $signed(input_fmap_0[15:0]) +
	( 16'sd 31118) * $signed(input_fmap_1[15:0]) +
	( 16'sd 25260) * $signed(input_fmap_2[15:0]) +
	( 15'sd 9939) * $signed(input_fmap_3[15:0]) +
	( 13'sd 3546) * $signed(input_fmap_4[15:0]) +
	( 16'sd 21016) * $signed(input_fmap_5[15:0]) +
	( 15'sd 8823) * $signed(input_fmap_6[15:0]) +
	( 16'sd 30371) * $signed(input_fmap_7[15:0]) +
	( 13'sd 3217) * $signed(input_fmap_8[15:0]) +
	( 15'sd 10082) * $signed(input_fmap_9[15:0]) +
	( 16'sd 30292) * $signed(input_fmap_10[15:0]) +
	( 15'sd 14987) * $signed(input_fmap_11[15:0]) +
	( 16'sd 31857) * $signed(input_fmap_12[15:0]) +
	( 14'sd 7564) * $signed(input_fmap_13[15:0]) +
	( 16'sd 26798) * $signed(input_fmap_14[15:0]) +
	( 16'sd 25057) * $signed(input_fmap_15[15:0]) +
	( 15'sd 11812) * $signed(input_fmap_16[15:0]) +
	( 16'sd 30997) * $signed(input_fmap_17[15:0]) +
	( 16'sd 27407) * $signed(input_fmap_18[15:0]) +
	( 13'sd 3136) * $signed(input_fmap_19[15:0]) +
	( 16'sd 28994) * $signed(input_fmap_20[15:0]) +
	( 15'sd 8366) * $signed(input_fmap_21[15:0]) +
	( 14'sd 7209) * $signed(input_fmap_22[15:0]) +
	( 15'sd 9397) * $signed(input_fmap_23[15:0]) +
	( 15'sd 14108) * $signed(input_fmap_24[15:0]) +
	( 15'sd 14051) * $signed(input_fmap_25[15:0]) +
	( 16'sd 28231) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1803) * $signed(input_fmap_27[15:0]) +
	( 13'sd 3074) * $signed(input_fmap_28[15:0]) +
	( 16'sd 22647) * $signed(input_fmap_29[15:0]) +
	( 13'sd 4016) * $signed(input_fmap_30[15:0]) +
	( 15'sd 10941) * $signed(input_fmap_31[15:0]) +
	( 16'sd 25666) * $signed(input_fmap_32[15:0]) +
	( 16'sd 17108) * $signed(input_fmap_33[15:0]) +
	( 15'sd 14564) * $signed(input_fmap_34[15:0]) +
	( 15'sd 10428) * $signed(input_fmap_35[15:0]) +
	( 15'sd 11902) * $signed(input_fmap_36[15:0]) +
	( 14'sd 7431) * $signed(input_fmap_37[15:0]) +
	( 16'sd 17282) * $signed(input_fmap_38[15:0]) +
	( 15'sd 14225) * $signed(input_fmap_39[15:0]) +
	( 16'sd 17048) * $signed(input_fmap_40[15:0]) +
	( 16'sd 32408) * $signed(input_fmap_41[15:0]) +
	( 16'sd 17042) * $signed(input_fmap_42[15:0]) +
	( 14'sd 5511) * $signed(input_fmap_43[15:0]) +
	( 16'sd 29868) * $signed(input_fmap_44[15:0]) +
	( 16'sd 24761) * $signed(input_fmap_45[15:0]) +
	( 16'sd 23126) * $signed(input_fmap_46[15:0]) +
	( 15'sd 12420) * $signed(input_fmap_47[15:0]) +
	( 14'sd 6526) * $signed(input_fmap_48[15:0]) +
	( 14'sd 7764) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22721) * $signed(input_fmap_50[15:0]) +
	( 15'sd 14042) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19377) * $signed(input_fmap_52[15:0]) +
	( 15'sd 13737) * $signed(input_fmap_53[15:0]) +
	( 13'sd 2866) * $signed(input_fmap_54[15:0]) +
	( 15'sd 13288) * $signed(input_fmap_55[15:0]) +
	( 16'sd 19826) * $signed(input_fmap_56[15:0]) +
	( 16'sd 21994) * $signed(input_fmap_57[15:0]) +
	( 13'sd 3489) * $signed(input_fmap_58[15:0]) +
	( 16'sd 22366) * $signed(input_fmap_59[15:0]) +
	( 15'sd 8646) * $signed(input_fmap_60[15:0]) +
	( 15'sd 14647) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3239) * $signed(input_fmap_62[15:0]) +
	( 16'sd 18028) * $signed(input_fmap_63[15:0]) +
	( 14'sd 6601) * $signed(input_fmap_64[15:0]) +
	( 16'sd 25015) * $signed(input_fmap_65[15:0]) +
	( 15'sd 14240) * $signed(input_fmap_66[15:0]) +
	( 16'sd 31319) * $signed(input_fmap_67[15:0]) +
	( 10'sd 462) * $signed(input_fmap_68[15:0]) +
	( 16'sd 22769) * $signed(input_fmap_69[15:0]) +
	( 15'sd 14045) * $signed(input_fmap_70[15:0]) +
	( 16'sd 28479) * $signed(input_fmap_71[15:0]) +
	( 12'sd 1691) * $signed(input_fmap_72[15:0]) +
	( 16'sd 28178) * $signed(input_fmap_73[15:0]) +
	( 16'sd 23582) * $signed(input_fmap_74[15:0]) +
	( 14'sd 5984) * $signed(input_fmap_75[15:0]) +
	( 16'sd 20224) * $signed(input_fmap_76[15:0]) +
	( 16'sd 29578) * $signed(input_fmap_77[15:0]) +
	( 14'sd 6962) * $signed(input_fmap_78[15:0]) +
	( 16'sd 28491) * $signed(input_fmap_79[15:0]) +
	( 16'sd 20798) * $signed(input_fmap_80[15:0]) +
	( 15'sd 16378) * $signed(input_fmap_81[15:0]) +
	( 15'sd 10742) * $signed(input_fmap_82[15:0]) +
	( 16'sd 24739) * $signed(input_fmap_83[15:0]) +
	( 16'sd 26272) * $signed(input_fmap_84[15:0]) +
	( 14'sd 6073) * $signed(input_fmap_85[15:0]) +
	( 16'sd 22945) * $signed(input_fmap_86[15:0]) +
	( 15'sd 9621) * $signed(input_fmap_87[15:0]) +
	( 16'sd 31879) * $signed(input_fmap_88[15:0]) +
	( 16'sd 28865) * $signed(input_fmap_89[15:0]) +
	( 16'sd 32390) * $signed(input_fmap_90[15:0]) +
	( 16'sd 20116) * $signed(input_fmap_91[15:0]) +
	( 14'sd 8164) * $signed(input_fmap_92[15:0]) +
	( 12'sd 2003) * $signed(input_fmap_93[15:0]) +
	( 15'sd 10544) * $signed(input_fmap_94[15:0]) +
	( 16'sd 17537) * $signed(input_fmap_95[15:0]) +
	( 16'sd 23083) * $signed(input_fmap_96[15:0]) +
	( 14'sd 4898) * $signed(input_fmap_97[15:0]) +
	( 14'sd 5293) * $signed(input_fmap_98[15:0]) +
	( 16'sd 21691) * $signed(input_fmap_99[15:0]) +
	( 16'sd 20739) * $signed(input_fmap_100[15:0]) +
	( 15'sd 10032) * $signed(input_fmap_101[15:0]) +
	( 16'sd 26590) * $signed(input_fmap_102[15:0]) +
	( 16'sd 17010) * $signed(input_fmap_103[15:0]) +
	( 15'sd 10441) * $signed(input_fmap_104[15:0]) +
	( 15'sd 12318) * $signed(input_fmap_105[15:0]) +
	( 15'sd 9311) * $signed(input_fmap_106[15:0]) +
	( 16'sd 27702) * $signed(input_fmap_107[15:0]) +
	( 13'sd 2722) * $signed(input_fmap_108[15:0]) +
	( 13'sd 3422) * $signed(input_fmap_109[15:0]) +
	( 15'sd 12418) * $signed(input_fmap_110[15:0]) +
	( 16'sd 17915) * $signed(input_fmap_111[15:0]) +
	( 8'sd 114) * $signed(input_fmap_112[15:0]) +
	( 16'sd 31762) * $signed(input_fmap_113[15:0]) +
	( 14'sd 5466) * $signed(input_fmap_114[15:0]) +
	( 14'sd 4675) * $signed(input_fmap_115[15:0]) +
	( 16'sd 20729) * $signed(input_fmap_116[15:0]) +
	( 15'sd 13932) * $signed(input_fmap_117[15:0]) +
	( 16'sd 29594) * $signed(input_fmap_118[15:0]) +
	( 14'sd 6822) * $signed(input_fmap_119[15:0]) +
	( 16'sd 21437) * $signed(input_fmap_120[15:0]) +
	( 15'sd 10734) * $signed(input_fmap_121[15:0]) +
	( 15'sd 9568) * $signed(input_fmap_122[15:0]) +
	( 16'sd 23604) * $signed(input_fmap_123[15:0]) +
	( 15'sd 15628) * $signed(input_fmap_124[15:0]) +
	( 12'sd 1928) * $signed(input_fmap_125[15:0]) +
	( 15'sd 14533) * $signed(input_fmap_126[15:0]) +
	( 14'sd 6545) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 16'sd 30288) * $signed(input_fmap_0[15:0]) +
	( 16'sd 31488) * $signed(input_fmap_1[15:0]) +
	( 16'sd 18701) * $signed(input_fmap_2[15:0]) +
	( 16'sd 31465) * $signed(input_fmap_3[15:0]) +
	( 13'sd 2813) * $signed(input_fmap_4[15:0]) +
	( 16'sd 30490) * $signed(input_fmap_5[15:0]) +
	( 12'sd 1582) * $signed(input_fmap_6[15:0]) +
	( 16'sd 18664) * $signed(input_fmap_7[15:0]) +
	( 14'sd 7178) * $signed(input_fmap_8[15:0]) +
	( 15'sd 9799) * $signed(input_fmap_9[15:0]) +
	( 16'sd 28184) * $signed(input_fmap_10[15:0]) +
	( 16'sd 30500) * $signed(input_fmap_11[15:0]) +
	( 16'sd 29525) * $signed(input_fmap_12[15:0]) +
	( 15'sd 11434) * $signed(input_fmap_13[15:0]) +
	( 16'sd 24843) * $signed(input_fmap_14[15:0]) +
	( 14'sd 4800) * $signed(input_fmap_15[15:0]) +
	( 14'sd 5631) * $signed(input_fmap_16[15:0]) +
	( 13'sd 3183) * $signed(input_fmap_17[15:0]) +
	( 16'sd 16978) * $signed(input_fmap_18[15:0]) +
	( 16'sd 32383) * $signed(input_fmap_19[15:0]) +
	( 14'sd 4349) * $signed(input_fmap_20[15:0]) +
	( 16'sd 19476) * $signed(input_fmap_21[15:0]) +
	( 16'sd 29806) * $signed(input_fmap_22[15:0]) +
	( 14'sd 7094) * $signed(input_fmap_23[15:0]) +
	( 16'sd 17988) * $signed(input_fmap_24[15:0]) +
	( 16'sd 21433) * $signed(input_fmap_25[15:0]) +
	( 16'sd 29584) * $signed(input_fmap_26[15:0]) +
	( 16'sd 28301) * $signed(input_fmap_27[15:0]) +
	( 16'sd 21509) * $signed(input_fmap_28[15:0]) +
	( 15'sd 13876) * $signed(input_fmap_29[15:0]) +
	( 16'sd 24019) * $signed(input_fmap_30[15:0]) +
	( 16'sd 21658) * $signed(input_fmap_31[15:0]) +
	( 16'sd 18163) * $signed(input_fmap_32[15:0]) +
	( 16'sd 26102) * $signed(input_fmap_33[15:0]) +
	( 16'sd 21113) * $signed(input_fmap_34[15:0]) +
	( 15'sd 9969) * $signed(input_fmap_35[15:0]) +
	( 16'sd 21940) * $signed(input_fmap_36[15:0]) +
	( 15'sd 15787) * $signed(input_fmap_37[15:0]) +
	( 11'sd 797) * $signed(input_fmap_38[15:0]) +
	( 16'sd 19138) * $signed(input_fmap_39[15:0]) +
	( 16'sd 22609) * $signed(input_fmap_40[15:0]) +
	( 14'sd 6476) * $signed(input_fmap_41[15:0]) +
	( 16'sd 21897) * $signed(input_fmap_42[15:0]) +
	( 15'sd 14635) * $signed(input_fmap_43[15:0]) +
	( 15'sd 15317) * $signed(input_fmap_44[15:0]) +
	( 12'sd 1633) * $signed(input_fmap_45[15:0]) +
	( 16'sd 19083) * $signed(input_fmap_46[15:0]) +
	( 14'sd 7382) * $signed(input_fmap_47[15:0]) +
	( 16'sd 25505) * $signed(input_fmap_48[15:0]) +
	( 15'sd 15382) * $signed(input_fmap_49[15:0]) +
	( 15'sd 12869) * $signed(input_fmap_50[15:0]) +
	( 16'sd 18961) * $signed(input_fmap_51[15:0]) +
	( 16'sd 22736) * $signed(input_fmap_52[15:0]) +
	( 15'sd 9502) * $signed(input_fmap_53[15:0]) +
	( 16'sd 17580) * $signed(input_fmap_54[15:0]) +
	( 16'sd 19917) * $signed(input_fmap_55[15:0]) +
	( 15'sd 13045) * $signed(input_fmap_56[15:0]) +
	( 16'sd 30850) * $signed(input_fmap_57[15:0]) +
	( 12'sd 1353) * $signed(input_fmap_58[15:0]) +
	( 15'sd 10194) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1872) * $signed(input_fmap_60[15:0]) +
	( 15'sd 13985) * $signed(input_fmap_61[15:0]) +
	( 16'sd 31182) * $signed(input_fmap_62[15:0]) +
	( 11'sd 718) * $signed(input_fmap_63[15:0]) +
	( 13'sd 2239) * $signed(input_fmap_64[15:0]) +
	( 16'sd 28436) * $signed(input_fmap_65[15:0]) +
	( 16'sd 24375) * $signed(input_fmap_66[15:0]) +
	( 15'sd 12115) * $signed(input_fmap_67[15:0]) +
	( 16'sd 21946) * $signed(input_fmap_68[15:0]) +
	( 16'sd 24165) * $signed(input_fmap_69[15:0]) +
	( 16'sd 17032) * $signed(input_fmap_70[15:0]) +
	( 16'sd 23551) * $signed(input_fmap_71[15:0]) +
	( 15'sd 15222) * $signed(input_fmap_72[15:0]) +
	( 14'sd 5731) * $signed(input_fmap_73[15:0]) +
	( 15'sd 14446) * $signed(input_fmap_74[15:0]) +
	( 14'sd 5487) * $signed(input_fmap_75[15:0]) +
	( 15'sd 15516) * $signed(input_fmap_76[15:0]) +
	( 11'sd 894) * $signed(input_fmap_77[15:0]) +
	( 12'sd 1252) * $signed(input_fmap_78[15:0]) +
	( 16'sd 17855) * $signed(input_fmap_79[15:0]) +
	( 12'sd 1205) * $signed(input_fmap_80[15:0]) +
	( 16'sd 30919) * $signed(input_fmap_81[15:0]) +
	( 16'sd 23352) * $signed(input_fmap_82[15:0]) +
	( 10'sd 332) * $signed(input_fmap_83[15:0]) +
	( 15'sd 14800) * $signed(input_fmap_84[15:0]) +
	( 16'sd 24611) * $signed(input_fmap_85[15:0]) +
	( 12'sd 1286) * $signed(input_fmap_86[15:0]) +
	( 16'sd 21370) * $signed(input_fmap_87[15:0]) +
	( 16'sd 31633) * $signed(input_fmap_88[15:0]) +
	( 16'sd 16435) * $signed(input_fmap_89[15:0]) +
	( 12'sd 1440) * $signed(input_fmap_90[15:0]) +
	( 15'sd 9639) * $signed(input_fmap_91[15:0]) +
	( 14'sd 6854) * $signed(input_fmap_92[15:0]) +
	( 12'sd 1092) * $signed(input_fmap_93[15:0]) +
	( 13'sd 2436) * $signed(input_fmap_94[15:0]) +
	( 16'sd 18188) * $signed(input_fmap_95[15:0]) +
	( 13'sd 2288) * $signed(input_fmap_96[15:0]) +
	( 16'sd 20348) * $signed(input_fmap_97[15:0]) +
	( 16'sd 24732) * $signed(input_fmap_98[15:0]) +
	( 16'sd 17410) * $signed(input_fmap_99[15:0]) +
	( 14'sd 4699) * $signed(input_fmap_100[15:0]) +
	( 11'sd 722) * $signed(input_fmap_101[15:0]) +
	( 14'sd 7925) * $signed(input_fmap_102[15:0]) +
	( 16'sd 25182) * $signed(input_fmap_103[15:0]) +
	( 16'sd 24299) * $signed(input_fmap_104[15:0]) +
	( 15'sd 11227) * $signed(input_fmap_105[15:0]) +
	( 16'sd 28458) * $signed(input_fmap_106[15:0]) +
	( 16'sd 29685) * $signed(input_fmap_107[15:0]) +
	( 12'sd 1248) * $signed(input_fmap_108[15:0]) +
	( 15'sd 16185) * $signed(input_fmap_109[15:0]) +
	( 16'sd 26009) * $signed(input_fmap_110[15:0]) +
	( 14'sd 4174) * $signed(input_fmap_111[15:0]) +
	( 14'sd 6561) * $signed(input_fmap_112[15:0]) +
	( 16'sd 20304) * $signed(input_fmap_113[15:0]) +
	( 13'sd 2449) * $signed(input_fmap_114[15:0]) +
	( 15'sd 14997) * $signed(input_fmap_115[15:0]) +
	( 15'sd 16147) * $signed(input_fmap_116[15:0]) +
	( 15'sd 9567) * $signed(input_fmap_117[15:0]) +
	( 16'sd 30793) * $signed(input_fmap_118[15:0]) +
	( 16'sd 23451) * $signed(input_fmap_119[15:0]) +
	( 15'sd 15834) * $signed(input_fmap_120[15:0]) +
	( 16'sd 24788) * $signed(input_fmap_121[15:0]) +
	( 14'sd 4173) * $signed(input_fmap_122[15:0]) +
	( 16'sd 24289) * $signed(input_fmap_123[15:0]) +
	( 16'sd 21675) * $signed(input_fmap_124[15:0]) +
	( 16'sd 28149) * $signed(input_fmap_125[15:0]) +
	( 15'sd 15788) * $signed(input_fmap_126[15:0]) +
	( 15'sd 11496) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 13'sd 2428) * $signed(input_fmap_0[15:0]) +
	( 16'sd 27164) * $signed(input_fmap_1[15:0]) +
	( 11'sd 859) * $signed(input_fmap_2[15:0]) +
	( 16'sd 24347) * $signed(input_fmap_3[15:0]) +
	( 16'sd 25425) * $signed(input_fmap_4[15:0]) +
	( 15'sd 12812) * $signed(input_fmap_5[15:0]) +
	( 12'sd 1399) * $signed(input_fmap_6[15:0]) +
	( 13'sd 2560) * $signed(input_fmap_7[15:0]) +
	( 10'sd 486) * $signed(input_fmap_8[15:0]) +
	( 15'sd 13164) * $signed(input_fmap_9[15:0]) +
	( 14'sd 4708) * $signed(input_fmap_10[15:0]) +
	( 15'sd 16256) * $signed(input_fmap_11[15:0]) +
	( 16'sd 22746) * $signed(input_fmap_12[15:0]) +
	( 14'sd 6362) * $signed(input_fmap_13[15:0]) +
	( 16'sd 20368) * $signed(input_fmap_14[15:0]) +
	( 16'sd 17269) * $signed(input_fmap_15[15:0]) +
	( 15'sd 11413) * $signed(input_fmap_16[15:0]) +
	( 16'sd 21278) * $signed(input_fmap_17[15:0]) +
	( 16'sd 16473) * $signed(input_fmap_18[15:0]) +
	( 15'sd 11777) * $signed(input_fmap_19[15:0]) +
	( 15'sd 16336) * $signed(input_fmap_20[15:0]) +
	( 16'sd 18751) * $signed(input_fmap_21[15:0]) +
	( 15'sd 13459) * $signed(input_fmap_22[15:0]) +
	( 15'sd 13547) * $signed(input_fmap_23[15:0]) +
	( 9'sd 163) * $signed(input_fmap_24[15:0]) +
	( 16'sd 16539) * $signed(input_fmap_25[15:0]) +
	( 15'sd 14790) * $signed(input_fmap_26[15:0]) +
	( 16'sd 31071) * $signed(input_fmap_27[15:0]) +
	( 16'sd 23693) * $signed(input_fmap_28[15:0]) +
	( 13'sd 4022) * $signed(input_fmap_29[15:0]) +
	( 16'sd 25058) * $signed(input_fmap_30[15:0]) +
	( 16'sd 20815) * $signed(input_fmap_31[15:0]) +
	( 16'sd 24600) * $signed(input_fmap_32[15:0]) +
	( 16'sd 24000) * $signed(input_fmap_33[15:0]) +
	( 16'sd 24500) * $signed(input_fmap_34[15:0]) +
	( 16'sd 20450) * $signed(input_fmap_35[15:0]) +
	( 16'sd 25241) * $signed(input_fmap_36[15:0]) +
	( 15'sd 14305) * $signed(input_fmap_37[15:0]) +
	( 16'sd 20166) * $signed(input_fmap_38[15:0]) +
	( 16'sd 23675) * $signed(input_fmap_39[15:0]) +
	( 16'sd 26637) * $signed(input_fmap_40[15:0]) +
	( 13'sd 2086) * $signed(input_fmap_41[15:0]) +
	( 15'sd 10545) * $signed(input_fmap_42[15:0]) +
	( 16'sd 21939) * $signed(input_fmap_43[15:0]) +
	( 15'sd 10440) * $signed(input_fmap_44[15:0]) +
	( 16'sd 18480) * $signed(input_fmap_45[15:0]) +
	( 14'sd 5735) * $signed(input_fmap_46[15:0]) +
	( 16'sd 22109) * $signed(input_fmap_47[15:0]) +
	( 15'sd 12743) * $signed(input_fmap_48[15:0]) +
	( 15'sd 14172) * $signed(input_fmap_49[15:0]) +
	( 16'sd 17059) * $signed(input_fmap_50[15:0]) +
	( 10'sd 290) * $signed(input_fmap_51[15:0]) +
	( 12'sd 1223) * $signed(input_fmap_52[15:0]) +
	( 16'sd 24302) * $signed(input_fmap_53[15:0]) +
	( 14'sd 4862) * $signed(input_fmap_54[15:0]) +
	( 16'sd 26024) * $signed(input_fmap_55[15:0]) +
	( 16'sd 25179) * $signed(input_fmap_56[15:0]) +
	( 11'sd 1004) * $signed(input_fmap_57[15:0]) +
	( 15'sd 9017) * $signed(input_fmap_58[15:0]) +
	( 15'sd 15869) * $signed(input_fmap_59[15:0]) +
	( 16'sd 20816) * $signed(input_fmap_60[15:0]) +
	( 15'sd 9030) * $signed(input_fmap_61[15:0]) +
	( 13'sd 3565) * $signed(input_fmap_62[15:0]) +
	( 15'sd 12849) * $signed(input_fmap_63[15:0]) +
	( 16'sd 31765) * $signed(input_fmap_64[15:0]) +
	( 16'sd 26090) * $signed(input_fmap_65[15:0]) +
	( 14'sd 7171) * $signed(input_fmap_66[15:0]) +
	( 16'sd 16648) * $signed(input_fmap_67[15:0]) +
	( 16'sd 18087) * $signed(input_fmap_68[15:0]) +
	( 16'sd 23653) * $signed(input_fmap_69[15:0]) +
	( 16'sd 20506) * $signed(input_fmap_70[15:0]) +
	( 15'sd 14107) * $signed(input_fmap_71[15:0]) +
	( 15'sd 15969) * $signed(input_fmap_72[15:0]) +
	( 16'sd 19087) * $signed(input_fmap_73[15:0]) +
	( 16'sd 16932) * $signed(input_fmap_74[15:0]) +
	( 16'sd 16907) * $signed(input_fmap_75[15:0]) +
	( 16'sd 21782) * $signed(input_fmap_76[15:0]) +
	( 12'sd 1046) * $signed(input_fmap_77[15:0]) +
	( 15'sd 11485) * $signed(input_fmap_78[15:0]) +
	( 16'sd 23137) * $signed(input_fmap_79[15:0]) +
	( 15'sd 14140) * $signed(input_fmap_80[15:0]) +
	( 15'sd 10232) * $signed(input_fmap_81[15:0]) +
	( 15'sd 12923) * $signed(input_fmap_82[15:0]) +
	( 15'sd 15819) * $signed(input_fmap_83[15:0]) +
	( 16'sd 31572) * $signed(input_fmap_84[15:0]) +
	( 15'sd 15031) * $signed(input_fmap_85[15:0]) +
	( 15'sd 16332) * $signed(input_fmap_86[15:0]) +
	( 16'sd 20582) * $signed(input_fmap_87[15:0]) +
	( 16'sd 22352) * $signed(input_fmap_88[15:0]) +
	( 13'sd 2155) * $signed(input_fmap_89[15:0]) +
	( 16'sd 29081) * $signed(input_fmap_90[15:0]) +
	( 16'sd 21772) * $signed(input_fmap_91[15:0]) +
	( 16'sd 26027) * $signed(input_fmap_92[15:0]) +
	( 13'sd 3423) * $signed(input_fmap_93[15:0]) +
	( 16'sd 32202) * $signed(input_fmap_94[15:0]) +
	( 16'sd 20645) * $signed(input_fmap_95[15:0]) +
	( 16'sd 32709) * $signed(input_fmap_96[15:0]) +
	( 16'sd 18504) * $signed(input_fmap_97[15:0]) +
	( 16'sd 31910) * $signed(input_fmap_98[15:0]) +
	( 16'sd 17893) * $signed(input_fmap_99[15:0]) +
	( 16'sd 29773) * $signed(input_fmap_100[15:0]) +
	( 16'sd 17561) * $signed(input_fmap_101[15:0]) +
	( 14'sd 6380) * $signed(input_fmap_102[15:0]) +
	( 16'sd 16552) * $signed(input_fmap_103[15:0]) +
	( 16'sd 26550) * $signed(input_fmap_104[15:0]) +
	( 16'sd 20610) * $signed(input_fmap_105[15:0]) +
	( 16'sd 23329) * $signed(input_fmap_106[15:0]) +
	( 16'sd 31928) * $signed(input_fmap_107[15:0]) +
	( 15'sd 14425) * $signed(input_fmap_108[15:0]) +
	( 14'sd 6705) * $signed(input_fmap_109[15:0]) +
	( 16'sd 23855) * $signed(input_fmap_110[15:0]) +
	( 15'sd 10658) * $signed(input_fmap_111[15:0]) +
	( 16'sd 26368) * $signed(input_fmap_112[15:0]) +
	( 11'sd 624) * $signed(input_fmap_113[15:0]) +
	( 16'sd 20505) * $signed(input_fmap_114[15:0]) +
	( 15'sd 10449) * $signed(input_fmap_115[15:0]) +
	( 16'sd 27211) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27072) * $signed(input_fmap_117[15:0]) +
	( 15'sd 16177) * $signed(input_fmap_118[15:0]) +
	( 15'sd 16189) * $signed(input_fmap_119[15:0]) +
	( 15'sd 15085) * $signed(input_fmap_120[15:0]) +
	( 15'sd 12115) * $signed(input_fmap_121[15:0]) +
	( 15'sd 8702) * $signed(input_fmap_122[15:0]) +
	( 16'sd 22180) * $signed(input_fmap_123[15:0]) +
	( 15'sd 12054) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24700) * $signed(input_fmap_125[15:0]) +
	( 16'sd 20325) * $signed(input_fmap_126[15:0]) +
	( 15'sd 11795) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 15'sd 12967) * $signed(input_fmap_0[15:0]) +
	( 15'sd 9351) * $signed(input_fmap_1[15:0]) +
	( 15'sd 14619) * $signed(input_fmap_2[15:0]) +
	( 16'sd 20143) * $signed(input_fmap_3[15:0]) +
	( 16'sd 25630) * $signed(input_fmap_4[15:0]) +
	( 16'sd 27085) * $signed(input_fmap_5[15:0]) +
	( 13'sd 3509) * $signed(input_fmap_6[15:0]) +
	( 16'sd 25918) * $signed(input_fmap_7[15:0]) +
	( 16'sd 17928) * $signed(input_fmap_8[15:0]) +
	( 15'sd 14328) * $signed(input_fmap_9[15:0]) +
	( 15'sd 10454) * $signed(input_fmap_10[15:0]) +
	( 16'sd 18873) * $signed(input_fmap_11[15:0]) +
	( 15'sd 10991) * $signed(input_fmap_12[15:0]) +
	( 13'sd 3466) * $signed(input_fmap_13[15:0]) +
	( 16'sd 16846) * $signed(input_fmap_14[15:0]) +
	( 14'sd 6999) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10686) * $signed(input_fmap_16[15:0]) +
	( 16'sd 29632) * $signed(input_fmap_17[15:0]) +
	( 14'sd 5907) * $signed(input_fmap_18[15:0]) +
	( 16'sd 21730) * $signed(input_fmap_19[15:0]) +
	( 15'sd 13238) * $signed(input_fmap_20[15:0]) +
	( 16'sd 18094) * $signed(input_fmap_21[15:0]) +
	( 16'sd 21108) * $signed(input_fmap_22[15:0]) +
	( 13'sd 3259) * $signed(input_fmap_23[15:0]) +
	( 15'sd 12145) * $signed(input_fmap_24[15:0]) +
	( 15'sd 15361) * $signed(input_fmap_25[15:0]) +
	( 14'sd 6836) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2584) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24356) * $signed(input_fmap_28[15:0]) +
	( 16'sd 18723) * $signed(input_fmap_29[15:0]) +
	( 16'sd 27578) * $signed(input_fmap_30[15:0]) +
	( 9'sd 131) * $signed(input_fmap_31[15:0]) +
	( 15'sd 14884) * $signed(input_fmap_32[15:0]) +
	( 14'sd 7907) * $signed(input_fmap_33[15:0]) +
	( 16'sd 17887) * $signed(input_fmap_34[15:0]) +
	( 16'sd 27935) * $signed(input_fmap_35[15:0]) +
	( 16'sd 31562) * $signed(input_fmap_36[15:0]) +
	( 16'sd 27723) * $signed(input_fmap_37[15:0]) +
	( 16'sd 29379) * $signed(input_fmap_38[15:0]) +
	( 13'sd 3699) * $signed(input_fmap_39[15:0]) +
	( 14'sd 4455) * $signed(input_fmap_40[15:0]) +
	( 14'sd 6698) * $signed(input_fmap_41[15:0]) +
	( 16'sd 20461) * $signed(input_fmap_42[15:0]) +
	( 16'sd 26341) * $signed(input_fmap_43[15:0]) +
	( 11'sd 988) * $signed(input_fmap_44[15:0]) +
	( 16'sd 30035) * $signed(input_fmap_45[15:0]) +
	( 16'sd 20473) * $signed(input_fmap_46[15:0]) +
	( 16'sd 16701) * $signed(input_fmap_47[15:0]) +
	( 15'sd 12475) * $signed(input_fmap_48[15:0]) +
	( 16'sd 31546) * $signed(input_fmap_49[15:0]) +
	( 16'sd 32529) * $signed(input_fmap_50[15:0]) +
	( 15'sd 10319) * $signed(input_fmap_51[15:0]) +
	( 15'sd 13318) * $signed(input_fmap_52[15:0]) +
	( 13'sd 3169) * $signed(input_fmap_53[15:0]) +
	( 16'sd 30652) * $signed(input_fmap_54[15:0]) +
	( 16'sd 32453) * $signed(input_fmap_55[15:0]) +
	( 16'sd 17736) * $signed(input_fmap_56[15:0]) +
	( 14'sd 6637) * $signed(input_fmap_57[15:0]) +
	( 16'sd 24549) * $signed(input_fmap_58[15:0]) +
	( 16'sd 21982) * $signed(input_fmap_59[15:0]) +
	( 15'sd 14170) * $signed(input_fmap_60[15:0]) +
	( 16'sd 27316) * $signed(input_fmap_61[15:0]) +
	( 15'sd 10564) * $signed(input_fmap_62[15:0]) +
	( 14'sd 5925) * $signed(input_fmap_63[15:0]) +
	( 16'sd 23686) * $signed(input_fmap_64[15:0]) +
	( 16'sd 26944) * $signed(input_fmap_65[15:0]) +
	( 16'sd 31007) * $signed(input_fmap_66[15:0]) +
	( 15'sd 15427) * $signed(input_fmap_67[15:0]) +
	( 16'sd 30066) * $signed(input_fmap_68[15:0]) +
	( 15'sd 14789) * $signed(input_fmap_69[15:0]) +
	( 15'sd 11934) * $signed(input_fmap_70[15:0]) +
	( 14'sd 7542) * $signed(input_fmap_71[15:0]) +
	( 16'sd 32551) * $signed(input_fmap_72[15:0]) +
	( 15'sd 13718) * $signed(input_fmap_73[15:0]) +
	( 16'sd 31472) * $signed(input_fmap_74[15:0]) +
	( 15'sd 15531) * $signed(input_fmap_75[15:0]) +
	( 15'sd 11894) * $signed(input_fmap_76[15:0]) +
	( 16'sd 27562) * $signed(input_fmap_77[15:0]) +
	( 14'sd 6096) * $signed(input_fmap_78[15:0]) +
	( 14'sd 4644) * $signed(input_fmap_79[15:0]) +
	( 15'sd 11487) * $signed(input_fmap_80[15:0]) +
	( 12'sd 1083) * $signed(input_fmap_81[15:0]) +
	( 15'sd 14830) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25908) * $signed(input_fmap_83[15:0]) +
	( 11'sd 957) * $signed(input_fmap_84[15:0]) +
	( 16'sd 31959) * $signed(input_fmap_85[15:0]) +
	( 16'sd 29779) * $signed(input_fmap_86[15:0]) +
	( 14'sd 7074) * $signed(input_fmap_87[15:0]) +
	( 15'sd 9900) * $signed(input_fmap_88[15:0]) +
	( 14'sd 4528) * $signed(input_fmap_89[15:0]) +
	( 15'sd 8431) * $signed(input_fmap_90[15:0]) +
	( 16'sd 31963) * $signed(input_fmap_91[15:0]) +
	( 16'sd 32001) * $signed(input_fmap_92[15:0]) +
	( 12'sd 1311) * $signed(input_fmap_93[15:0]) +
	( 16'sd 21158) * $signed(input_fmap_94[15:0]) +
	( 15'sd 14761) * $signed(input_fmap_95[15:0]) +
	( 16'sd 26999) * $signed(input_fmap_96[15:0]) +
	( 12'sd 1911) * $signed(input_fmap_97[15:0]) +
	( 12'sd 1268) * $signed(input_fmap_98[15:0]) +
	( 16'sd 18377) * $signed(input_fmap_99[15:0]) +
	( 15'sd 15412) * $signed(input_fmap_100[15:0]) +
	( 16'sd 17587) * $signed(input_fmap_101[15:0]) +
	( 15'sd 10222) * $signed(input_fmap_102[15:0]) +
	( 15'sd 10323) * $signed(input_fmap_103[15:0]) +
	( 15'sd 12716) * $signed(input_fmap_104[15:0]) +
	( 16'sd 32680) * $signed(input_fmap_105[15:0]) +
	( 13'sd 3486) * $signed(input_fmap_106[15:0]) +
	( 14'sd 4859) * $signed(input_fmap_107[15:0]) +
	( 15'sd 11076) * $signed(input_fmap_108[15:0]) +
	( 10'sd 355) * $signed(input_fmap_109[15:0]) +
	( 12'sd 2047) * $signed(input_fmap_110[15:0]) +
	( 16'sd 24524) * $signed(input_fmap_111[15:0]) +
	( 16'sd 20031) * $signed(input_fmap_112[15:0]) +
	( 14'sd 8147) * $signed(input_fmap_113[15:0]) +
	( 16'sd 31099) * $signed(input_fmap_114[15:0]) +
	( 14'sd 7086) * $signed(input_fmap_115[15:0]) +
	( 14'sd 7914) * $signed(input_fmap_116[15:0]) +
	( 15'sd 13448) * $signed(input_fmap_117[15:0]) +
	( 14'sd 5203) * $signed(input_fmap_118[15:0]) +
	( 16'sd 20036) * $signed(input_fmap_119[15:0]) +
	( 16'sd 28964) * $signed(input_fmap_120[15:0]) +
	( 15'sd 10993) * $signed(input_fmap_121[15:0]) +
	( 16'sd 17747) * $signed(input_fmap_122[15:0]) +
	( 16'sd 27604) * $signed(input_fmap_123[15:0]) +
	( 14'sd 5047) * $signed(input_fmap_124[15:0]) +
	( 14'sd 6783) * $signed(input_fmap_125[15:0]) +
	( 14'sd 7368) * $signed(input_fmap_126[15:0]) +
	( 16'sd 30908) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 16'sd 17632) * $signed(input_fmap_0[15:0]) +
	( 16'sd 25388) * $signed(input_fmap_1[15:0]) +
	( 16'sd 22417) * $signed(input_fmap_2[15:0]) +
	( 16'sd 17055) * $signed(input_fmap_3[15:0]) +
	( 16'sd 23780) * $signed(input_fmap_4[15:0]) +
	( 10'sd 472) * $signed(input_fmap_5[15:0]) +
	( 16'sd 28521) * $signed(input_fmap_6[15:0]) +
	( 16'sd 21108) * $signed(input_fmap_7[15:0]) +
	( 14'sd 7838) * $signed(input_fmap_8[15:0]) +
	( 15'sd 8658) * $signed(input_fmap_9[15:0]) +
	( 15'sd 10961) * $signed(input_fmap_10[15:0]) +
	( 15'sd 8860) * $signed(input_fmap_11[15:0]) +
	( 16'sd 27023) * $signed(input_fmap_12[15:0]) +
	( 16'sd 21096) * $signed(input_fmap_13[15:0]) +
	( 16'sd 25688) * $signed(input_fmap_14[15:0]) +
	( 16'sd 29386) * $signed(input_fmap_15[15:0]) +
	( 16'sd 16467) * $signed(input_fmap_16[15:0]) +
	( 16'sd 20647) * $signed(input_fmap_17[15:0]) +
	( 12'sd 2004) * $signed(input_fmap_18[15:0]) +
	( 16'sd 31274) * $signed(input_fmap_19[15:0]) +
	( 15'sd 9897) * $signed(input_fmap_20[15:0]) +
	( 13'sd 4000) * $signed(input_fmap_21[15:0]) +
	( 10'sd 363) * $signed(input_fmap_22[15:0]) +
	( 16'sd 18769) * $signed(input_fmap_23[15:0]) +
	( 16'sd 31715) * $signed(input_fmap_24[15:0]) +
	( 15'sd 9002) * $signed(input_fmap_25[15:0]) +
	( 12'sd 1721) * $signed(input_fmap_26[15:0]) +
	( 14'sd 4277) * $signed(input_fmap_27[15:0]) +
	( 16'sd 23432) * $signed(input_fmap_28[15:0]) +
	( 16'sd 17171) * $signed(input_fmap_29[15:0]) +
	( 13'sd 3072) * $signed(input_fmap_30[15:0]) +
	( 15'sd 14524) * $signed(input_fmap_31[15:0]) +
	( 11'sd 725) * $signed(input_fmap_32[15:0]) +
	( 10'sd 370) * $signed(input_fmap_33[15:0]) +
	( 16'sd 22837) * $signed(input_fmap_34[15:0]) +
	( 15'sd 12045) * $signed(input_fmap_35[15:0]) +
	( 16'sd 23968) * $signed(input_fmap_36[15:0]) +
	( 12'sd 1081) * $signed(input_fmap_37[15:0]) +
	( 15'sd 11881) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24352) * $signed(input_fmap_39[15:0]) +
	( 13'sd 3260) * $signed(input_fmap_40[15:0]) +
	( 16'sd 29299) * $signed(input_fmap_41[15:0]) +
	( 16'sd 21984) * $signed(input_fmap_42[15:0]) +
	( 15'sd 9024) * $signed(input_fmap_43[15:0]) +
	( 15'sd 13005) * $signed(input_fmap_44[15:0]) +
	( 16'sd 31760) * $signed(input_fmap_45[15:0]) +
	( 16'sd 32262) * $signed(input_fmap_46[15:0]) +
	( 15'sd 11839) * $signed(input_fmap_47[15:0]) +
	( 15'sd 15787) * $signed(input_fmap_48[15:0]) +
	( 16'sd 28751) * $signed(input_fmap_49[15:0]) +
	( 15'sd 11405) * $signed(input_fmap_50[15:0]) +
	( 12'sd 1515) * $signed(input_fmap_51[15:0]) +
	( 15'sd 15454) * $signed(input_fmap_52[15:0]) +
	( 16'sd 27079) * $signed(input_fmap_53[15:0]) +
	( 15'sd 16159) * $signed(input_fmap_54[15:0]) +
	( 14'sd 5623) * $signed(input_fmap_55[15:0]) +
	( 14'sd 7381) * $signed(input_fmap_56[15:0]) +
	( 16'sd 18580) * $signed(input_fmap_57[15:0]) +
	( 15'sd 8636) * $signed(input_fmap_58[15:0]) +
	( 16'sd 25556) * $signed(input_fmap_59[15:0]) +
	( 16'sd 23845) * $signed(input_fmap_60[15:0]) +
	( 11'sd 628) * $signed(input_fmap_61[15:0]) +
	( 14'sd 5981) * $signed(input_fmap_62[15:0]) +
	( 16'sd 20251) * $signed(input_fmap_63[15:0]) +
	( 16'sd 22729) * $signed(input_fmap_64[15:0]) +
	( 15'sd 14111) * $signed(input_fmap_65[15:0]) +
	( 16'sd 29514) * $signed(input_fmap_66[15:0]) +
	( 16'sd 16784) * $signed(input_fmap_67[15:0]) +
	( 16'sd 17518) * $signed(input_fmap_68[15:0]) +
	( 16'sd 22445) * $signed(input_fmap_69[15:0]) +
	( 15'sd 13967) * $signed(input_fmap_70[15:0]) +
	( 13'sd 3219) * $signed(input_fmap_71[15:0]) +
	( 14'sd 6732) * $signed(input_fmap_72[15:0]) +
	( 16'sd 30123) * $signed(input_fmap_73[15:0]) +
	( 12'sd 1600) * $signed(input_fmap_74[15:0]) +
	( 14'sd 4703) * $signed(input_fmap_75[15:0]) +
	( 15'sd 12067) * $signed(input_fmap_76[15:0]) +
	( 14'sd 6748) * $signed(input_fmap_77[15:0]) +
	( 16'sd 23642) * $signed(input_fmap_78[15:0]) +
	( 15'sd 16339) * $signed(input_fmap_79[15:0]) +
	( 16'sd 29019) * $signed(input_fmap_80[15:0]) +
	( 16'sd 21592) * $signed(input_fmap_81[15:0]) +
	( 14'sd 7639) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25191) * $signed(input_fmap_83[15:0]) +
	( 16'sd 21736) * $signed(input_fmap_84[15:0]) +
	( 16'sd 30852) * $signed(input_fmap_85[15:0]) +
	( 14'sd 6622) * $signed(input_fmap_86[15:0]) +
	( 16'sd 29587) * $signed(input_fmap_87[15:0]) +
	( 16'sd 31251) * $signed(input_fmap_88[15:0]) +
	( 16'sd 21966) * $signed(input_fmap_89[15:0]) +
	( 16'sd 31303) * $signed(input_fmap_90[15:0]) +
	( 15'sd 13479) * $signed(input_fmap_91[15:0]) +
	( 16'sd 30816) * $signed(input_fmap_92[15:0]) +
	( 16'sd 17398) * $signed(input_fmap_93[15:0]) +
	( 15'sd 15301) * $signed(input_fmap_94[15:0]) +
	( 16'sd 22633) * $signed(input_fmap_95[15:0]) +
	( 16'sd 17156) * $signed(input_fmap_96[15:0]) +
	( 16'sd 24706) * $signed(input_fmap_97[15:0]) +
	( 15'sd 9454) * $signed(input_fmap_98[15:0]) +
	( 16'sd 22373) * $signed(input_fmap_99[15:0]) +
	( 15'sd 13638) * $signed(input_fmap_100[15:0]) +
	( 15'sd 11613) * $signed(input_fmap_101[15:0]) +
	( 13'sd 3626) * $signed(input_fmap_102[15:0]) +
	( 16'sd 30102) * $signed(input_fmap_103[15:0]) +
	( 16'sd 21722) * $signed(input_fmap_104[15:0]) +
	( 15'sd 11334) * $signed(input_fmap_105[15:0]) +
	( 16'sd 19447) * $signed(input_fmap_106[15:0]) +
	( 14'sd 7435) * $signed(input_fmap_107[15:0]) +
	( 15'sd 8355) * $signed(input_fmap_108[15:0]) +
	( 16'sd 19522) * $signed(input_fmap_109[15:0]) +
	( 15'sd 14957) * $signed(input_fmap_110[15:0]) +
	( 16'sd 28251) * $signed(input_fmap_111[15:0]) +
	( 15'sd 8223) * $signed(input_fmap_112[15:0]) +
	( 16'sd 18544) * $signed(input_fmap_113[15:0]) +
	( 16'sd 22730) * $signed(input_fmap_114[15:0]) +
	( 16'sd 23708) * $signed(input_fmap_115[15:0]) +
	( 15'sd 8890) * $signed(input_fmap_116[15:0]) +
	( 13'sd 3804) * $signed(input_fmap_117[15:0]) +
	( 14'sd 8083) * $signed(input_fmap_118[15:0]) +
	( 16'sd 18823) * $signed(input_fmap_119[15:0]) +
	( 16'sd 20446) * $signed(input_fmap_120[15:0]) +
	( 15'sd 11980) * $signed(input_fmap_121[15:0]) +
	( 16'sd 17722) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21097) * $signed(input_fmap_123[15:0]) +
	( 16'sd 26331) * $signed(input_fmap_124[15:0]) +
	( 16'sd 22899) * $signed(input_fmap_125[15:0]) +
	( 16'sd 32581) * $signed(input_fmap_126[15:0]) +
	( 15'sd 14929) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 16'sd 17628) * $signed(input_fmap_0[15:0]) +
	( 16'sd 26791) * $signed(input_fmap_1[15:0]) +
	( 15'sd 9730) * $signed(input_fmap_2[15:0]) +
	( 16'sd 28218) * $signed(input_fmap_3[15:0]) +
	( 12'sd 1442) * $signed(input_fmap_4[15:0]) +
	( 16'sd 27671) * $signed(input_fmap_5[15:0]) +
	( 16'sd 19015) * $signed(input_fmap_6[15:0]) +
	( 16'sd 25513) * $signed(input_fmap_7[15:0]) +
	( 15'sd 13325) * $signed(input_fmap_8[15:0]) +
	( 16'sd 19741) * $signed(input_fmap_9[15:0]) +
	( 16'sd 30595) * $signed(input_fmap_10[15:0]) +
	( 16'sd 20571) * $signed(input_fmap_11[15:0]) +
	( 14'sd 6214) * $signed(input_fmap_12[15:0]) +
	( 16'sd 26738) * $signed(input_fmap_13[15:0]) +
	( 12'sd 1046) * $signed(input_fmap_14[15:0]) +
	( 16'sd 32121) * $signed(input_fmap_15[15:0]) +
	( 14'sd 5050) * $signed(input_fmap_16[15:0]) +
	( 15'sd 12749) * $signed(input_fmap_17[15:0]) +
	( 16'sd 25027) * $signed(input_fmap_18[15:0]) +
	( 16'sd 24303) * $signed(input_fmap_19[15:0]) +
	( 13'sd 3357) * $signed(input_fmap_20[15:0]) +
	( 15'sd 14340) * $signed(input_fmap_21[15:0]) +
	( 15'sd 14385) * $signed(input_fmap_22[15:0]) +
	( 15'sd 14388) * $signed(input_fmap_23[15:0]) +
	( 14'sd 6783) * $signed(input_fmap_24[15:0]) +
	( 16'sd 25713) * $signed(input_fmap_25[15:0]) +
	( 13'sd 3750) * $signed(input_fmap_26[15:0]) +
	( 14'sd 5715) * $signed(input_fmap_27[15:0]) +
	( 16'sd 20757) * $signed(input_fmap_28[15:0]) +
	( 14'sd 4330) * $signed(input_fmap_29[15:0]) +
	( 14'sd 7215) * $signed(input_fmap_30[15:0]) +
	( 14'sd 5553) * $signed(input_fmap_31[15:0]) +
	( 9'sd 222) * $signed(input_fmap_32[15:0]) +
	( 16'sd 18857) * $signed(input_fmap_33[15:0]) +
	( 14'sd 7338) * $signed(input_fmap_34[15:0]) +
	( 16'sd 31033) * $signed(input_fmap_35[15:0]) +
	( 12'sd 1867) * $signed(input_fmap_36[15:0]) +
	( 16'sd 25801) * $signed(input_fmap_37[15:0]) +
	( 13'sd 2377) * $signed(input_fmap_38[15:0]) +
	( 16'sd 25357) * $signed(input_fmap_39[15:0]) +
	( 11'sd 636) * $signed(input_fmap_40[15:0]) +
	( 16'sd 29226) * $signed(input_fmap_41[15:0]) +
	( 16'sd 28646) * $signed(input_fmap_42[15:0]) +
	( 16'sd 24818) * $signed(input_fmap_43[15:0]) +
	( 16'sd 17855) * $signed(input_fmap_44[15:0]) +
	( 14'sd 7099) * $signed(input_fmap_45[15:0]) +
	( 16'sd 22878) * $signed(input_fmap_46[15:0]) +
	( 14'sd 4613) * $signed(input_fmap_47[15:0]) +
	( 16'sd 22603) * $signed(input_fmap_48[15:0]) +
	( 16'sd 31225) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22642) * $signed(input_fmap_50[15:0]) +
	( 11'sd 646) * $signed(input_fmap_51[15:0]) +
	( 14'sd 7531) * $signed(input_fmap_52[15:0]) +
	( 16'sd 30489) * $signed(input_fmap_53[15:0]) +
	( 13'sd 3132) * $signed(input_fmap_54[15:0]) +
	( 14'sd 8128) * $signed(input_fmap_55[15:0]) +
	( 15'sd 15380) * $signed(input_fmap_56[15:0]) +
	( 11'sd 1018) * $signed(input_fmap_57[15:0]) +
	( 16'sd 17899) * $signed(input_fmap_58[15:0]) +
	( 16'sd 20323) * $signed(input_fmap_59[15:0]) +
	( 16'sd 31282) * $signed(input_fmap_60[15:0]) +
	( 16'sd 29416) * $signed(input_fmap_61[15:0]) +
	( 15'sd 15347) * $signed(input_fmap_62[15:0]) +
	( 16'sd 32103) * $signed(input_fmap_63[15:0]) +
	( 15'sd 10306) * $signed(input_fmap_64[15:0]) +
	( 14'sd 7927) * $signed(input_fmap_65[15:0]) +
	( 16'sd 23930) * $signed(input_fmap_66[15:0]) +
	( 16'sd 20113) * $signed(input_fmap_67[15:0]) +
	( 16'sd 16872) * $signed(input_fmap_68[15:0]) +
	( 16'sd 26010) * $signed(input_fmap_69[15:0]) +
	( 14'sd 5521) * $signed(input_fmap_70[15:0]) +
	( 16'sd 29535) * $signed(input_fmap_71[15:0]) +
	( 16'sd 23387) * $signed(input_fmap_72[15:0]) +
	( 16'sd 27791) * $signed(input_fmap_73[15:0]) +
	( 13'sd 2184) * $signed(input_fmap_74[15:0]) +
	( 15'sd 14689) * $signed(input_fmap_75[15:0]) +
	( 16'sd 22103) * $signed(input_fmap_76[15:0]) +
	( 15'sd 13677) * $signed(input_fmap_77[15:0]) +
	( 14'sd 7187) * $signed(input_fmap_78[15:0]) +
	( 12'sd 1716) * $signed(input_fmap_79[15:0]) +
	( 13'sd 2221) * $signed(input_fmap_80[15:0]) +
	( 16'sd 20690) * $signed(input_fmap_81[15:0]) +
	( 15'sd 13218) * $signed(input_fmap_82[15:0]) +
	( 12'sd 1254) * $signed(input_fmap_83[15:0]) +
	( 14'sd 5266) * $signed(input_fmap_84[15:0]) +
	( 16'sd 21615) * $signed(input_fmap_85[15:0]) +
	( 16'sd 31021) * $signed(input_fmap_86[15:0]) +
	( 15'sd 14139) * $signed(input_fmap_87[15:0]) +
	( 16'sd 25966) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5487) * $signed(input_fmap_89[15:0]) +
	( 14'sd 5592) * $signed(input_fmap_90[15:0]) +
	( 14'sd 4629) * $signed(input_fmap_91[15:0]) +
	( 14'sd 7777) * $signed(input_fmap_92[15:0]) +
	( 16'sd 29414) * $signed(input_fmap_93[15:0]) +
	( 14'sd 6669) * $signed(input_fmap_94[15:0]) +
	( 16'sd 20829) * $signed(input_fmap_95[15:0]) +
	( 15'sd 8301) * $signed(input_fmap_96[15:0]) +
	( 13'sd 2282) * $signed(input_fmap_97[15:0]) +
	( 16'sd 20480) * $signed(input_fmap_98[15:0]) +
	( 14'sd 5226) * $signed(input_fmap_99[15:0]) +
	( 16'sd 23802) * $signed(input_fmap_100[15:0]) +
	( 15'sd 9670) * $signed(input_fmap_101[15:0]) +
	( 16'sd 23628) * $signed(input_fmap_102[15:0]) +
	( 16'sd 29293) * $signed(input_fmap_103[15:0]) +
	( 15'sd 15509) * $signed(input_fmap_104[15:0]) +
	( 10'sd 380) * $signed(input_fmap_105[15:0]) +
	( 16'sd 32049) * $signed(input_fmap_106[15:0]) +
	( 14'sd 4356) * $signed(input_fmap_107[15:0]) +
	( 14'sd 7438) * $signed(input_fmap_108[15:0]) +
	( 16'sd 17239) * $signed(input_fmap_109[15:0]) +
	( 16'sd 30210) * $signed(input_fmap_110[15:0]) +
	( 16'sd 28885) * $signed(input_fmap_111[15:0]) +
	( 16'sd 31964) * $signed(input_fmap_112[15:0]) +
	( 15'sd 12778) * $signed(input_fmap_113[15:0]) +
	( 13'sd 3658) * $signed(input_fmap_114[15:0]) +
	( 15'sd 9556) * $signed(input_fmap_115[15:0]) +
	( 15'sd 13592) * $signed(input_fmap_116[15:0]) +
	( 16'sd 32492) * $signed(input_fmap_117[15:0]) +
	( 16'sd 22497) * $signed(input_fmap_118[15:0]) +
	( 16'sd 29062) * $signed(input_fmap_119[15:0]) +
	( 16'sd 24054) * $signed(input_fmap_120[15:0]) +
	( 16'sd 31034) * $signed(input_fmap_121[15:0]) +
	( 16'sd 21019) * $signed(input_fmap_122[15:0]) +
	( 11'sd 821) * $signed(input_fmap_123[15:0]) +
	( 16'sd 20485) * $signed(input_fmap_124[15:0]) +
	( 16'sd 28015) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6469) * $signed(input_fmap_126[15:0]) +
	( 15'sd 15486) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 14'sd 4793) * $signed(input_fmap_0[15:0]) +
	( 13'sd 2672) * $signed(input_fmap_1[15:0]) +
	( 16'sd 20015) * $signed(input_fmap_2[15:0]) +
	( 16'sd 22447) * $signed(input_fmap_3[15:0]) +
	( 16'sd 30861) * $signed(input_fmap_4[15:0]) +
	( 16'sd 20762) * $signed(input_fmap_5[15:0]) +
	( 16'sd 22166) * $signed(input_fmap_6[15:0]) +
	( 16'sd 25464) * $signed(input_fmap_7[15:0]) +
	( 16'sd 25398) * $signed(input_fmap_8[15:0]) +
	( 16'sd 22014) * $signed(input_fmap_9[15:0]) +
	( 15'sd 14714) * $signed(input_fmap_10[15:0]) +
	( 15'sd 15377) * $signed(input_fmap_11[15:0]) +
	( 16'sd 25133) * $signed(input_fmap_12[15:0]) +
	( 15'sd 14042) * $signed(input_fmap_13[15:0]) +
	( 13'sd 2966) * $signed(input_fmap_14[15:0]) +
	( 16'sd 32763) * $signed(input_fmap_15[15:0]) +
	( 16'sd 19825) * $signed(input_fmap_16[15:0]) +
	( 16'sd 20284) * $signed(input_fmap_17[15:0]) +
	( 16'sd 25892) * $signed(input_fmap_18[15:0]) +
	( 15'sd 12610) * $signed(input_fmap_19[15:0]) +
	( 16'sd 21670) * $signed(input_fmap_20[15:0]) +
	( 14'sd 4294) * $signed(input_fmap_21[15:0]) +
	( 16'sd 18465) * $signed(input_fmap_22[15:0]) +
	( 16'sd 25537) * $signed(input_fmap_23[15:0]) +
	( 16'sd 21918) * $signed(input_fmap_24[15:0]) +
	( 16'sd 20831) * $signed(input_fmap_25[15:0]) +
	( 16'sd 19522) * $signed(input_fmap_26[15:0]) +
	( 15'sd 10290) * $signed(input_fmap_27[15:0]) +
	( 16'sd 25163) * $signed(input_fmap_28[15:0]) +
	( 15'sd 12471) * $signed(input_fmap_29[15:0]) +
	( 16'sd 30522) * $signed(input_fmap_30[15:0]) +
	( 15'sd 13686) * $signed(input_fmap_31[15:0]) +
	( 15'sd 10816) * $signed(input_fmap_32[15:0]) +
	( 15'sd 15090) * $signed(input_fmap_33[15:0]) +
	( 16'sd 31240) * $signed(input_fmap_34[15:0]) +
	( 15'sd 12499) * $signed(input_fmap_35[15:0]) +
	( 10'sd 298) * $signed(input_fmap_36[15:0]) +
	( 16'sd 32640) * $signed(input_fmap_37[15:0]) +
	( 14'sd 7218) * $signed(input_fmap_38[15:0]) +
	( 16'sd 29860) * $signed(input_fmap_39[15:0]) +
	( 16'sd 31232) * $signed(input_fmap_40[15:0]) +
	( 16'sd 27881) * $signed(input_fmap_41[15:0]) +
	( 16'sd 26367) * $signed(input_fmap_42[15:0]) +
	( 16'sd 20758) * $signed(input_fmap_43[15:0]) +
	( 16'sd 19379) * $signed(input_fmap_44[15:0]) +
	( 16'sd 18964) * $signed(input_fmap_45[15:0]) +
	( 15'sd 10916) * $signed(input_fmap_46[15:0]) +
	( 16'sd 24957) * $signed(input_fmap_47[15:0]) +
	( 15'sd 10063) * $signed(input_fmap_48[15:0]) +
	( 16'sd 23209) * $signed(input_fmap_49[15:0]) +
	( 13'sd 3385) * $signed(input_fmap_50[15:0]) +
	( 15'sd 14515) * $signed(input_fmap_51[15:0]) +
	( 16'sd 22735) * $signed(input_fmap_52[15:0]) +
	( 15'sd 8556) * $signed(input_fmap_53[15:0]) +
	( 13'sd 3489) * $signed(input_fmap_54[15:0]) +
	( 16'sd 32423) * $signed(input_fmap_55[15:0]) +
	( 15'sd 12327) * $signed(input_fmap_56[15:0]) +
	( 15'sd 11318) * $signed(input_fmap_57[15:0]) +
	( 16'sd 22747) * $signed(input_fmap_58[15:0]) +
	( 16'sd 19051) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1802) * $signed(input_fmap_60[15:0]) +
	( 15'sd 11993) * $signed(input_fmap_61[15:0]) +
	( 16'sd 24833) * $signed(input_fmap_62[15:0]) +
	( 11'sd 877) * $signed(input_fmap_63[15:0]) +
	( 16'sd 24089) * $signed(input_fmap_64[15:0]) +
	( 16'sd 20243) * $signed(input_fmap_65[15:0]) +
	( 16'sd 18139) * $signed(input_fmap_66[15:0]) +
	( 15'sd 10350) * $signed(input_fmap_67[15:0]) +
	( 16'sd 20568) * $signed(input_fmap_68[15:0]) +
	( 16'sd 21003) * $signed(input_fmap_69[15:0]) +
	( 15'sd 11177) * $signed(input_fmap_70[15:0]) +
	( 15'sd 14106) * $signed(input_fmap_71[15:0]) +
	( 15'sd 11348) * $signed(input_fmap_72[15:0]) +
	( 15'sd 8748) * $signed(input_fmap_73[15:0]) +
	( 16'sd 18826) * $signed(input_fmap_74[15:0]) +
	( 16'sd 28096) * $signed(input_fmap_75[15:0]) +
	( 13'sd 2706) * $signed(input_fmap_76[15:0]) +
	( 16'sd 18788) * $signed(input_fmap_77[15:0]) +
	( 16'sd 31313) * $signed(input_fmap_78[15:0]) +
	( 13'sd 2567) * $signed(input_fmap_79[15:0]) +
	( 16'sd 31918) * $signed(input_fmap_80[15:0]) +
	( 15'sd 13773) * $signed(input_fmap_81[15:0]) +
	( 16'sd 32013) * $signed(input_fmap_82[15:0]) +
	( 16'sd 30299) * $signed(input_fmap_83[15:0]) +
	( 15'sd 9957) * $signed(input_fmap_84[15:0]) +
	( 15'sd 12325) * $signed(input_fmap_85[15:0]) +
	( 16'sd 22697) * $signed(input_fmap_86[15:0]) +
	( 16'sd 19631) * $signed(input_fmap_87[15:0]) +
	( 14'sd 6244) * $signed(input_fmap_88[15:0]) +
	( 16'sd 19581) * $signed(input_fmap_89[15:0]) +
	( 16'sd 25807) * $signed(input_fmap_90[15:0]) +
	( 16'sd 31090) * $signed(input_fmap_91[15:0]) +
	( 16'sd 17612) * $signed(input_fmap_92[15:0]) +
	( 15'sd 11693) * $signed(input_fmap_93[15:0]) +
	( 16'sd 19404) * $signed(input_fmap_94[15:0]) +
	( 16'sd 30017) * $signed(input_fmap_95[15:0]) +
	( 16'sd 23423) * $signed(input_fmap_96[15:0]) +
	( 14'sd 6496) * $signed(input_fmap_97[15:0]) +
	( 16'sd 16473) * $signed(input_fmap_98[15:0]) +
	( 15'sd 12100) * $signed(input_fmap_99[15:0]) +
	( 15'sd 8560) * $signed(input_fmap_100[15:0]) +
	( 11'sd 521) * $signed(input_fmap_101[15:0]) +
	( 16'sd 25417) * $signed(input_fmap_102[15:0]) +
	( 13'sd 2926) * $signed(input_fmap_103[15:0]) +
	( 16'sd 18362) * $signed(input_fmap_104[15:0]) +
	( 16'sd 19159) * $signed(input_fmap_105[15:0]) +
	( 16'sd 31243) * $signed(input_fmap_106[15:0]) +
	( 15'sd 11857) * $signed(input_fmap_107[15:0]) +
	( 16'sd 22644) * $signed(input_fmap_108[15:0]) +
	( 16'sd 25658) * $signed(input_fmap_109[15:0]) +
	( 16'sd 31425) * $signed(input_fmap_110[15:0]) +
	( 16'sd 19410) * $signed(input_fmap_111[15:0]) +
	( 16'sd 32420) * $signed(input_fmap_112[15:0]) +
	( 15'sd 15883) * $signed(input_fmap_113[15:0]) +
	( 16'sd 19123) * $signed(input_fmap_114[15:0]) +
	( 16'sd 18598) * $signed(input_fmap_115[15:0]) +
	( 16'sd 23818) * $signed(input_fmap_116[15:0]) +
	( 13'sd 2773) * $signed(input_fmap_117[15:0]) +
	( 15'sd 15937) * $signed(input_fmap_118[15:0]) +
	( 15'sd 14519) * $signed(input_fmap_119[15:0]) +
	( 10'sd 386) * $signed(input_fmap_120[15:0]) +
	( 14'sd 8035) * $signed(input_fmap_121[15:0]) +
	( 15'sd 12693) * $signed(input_fmap_122[15:0]) +
	( 15'sd 11697) * $signed(input_fmap_123[15:0]) +
	( 16'sd 25674) * $signed(input_fmap_124[15:0]) +
	( 13'sd 2928) * $signed(input_fmap_125[15:0]) +
	( 14'sd 4286) * $signed(input_fmap_126[15:0]) +
	( 16'sd 26993) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 16'sd 28119) * $signed(input_fmap_0[15:0]) +
	( 16'sd 29348) * $signed(input_fmap_1[15:0]) +
	( 14'sd 6654) * $signed(input_fmap_2[15:0]) +
	( 15'sd 13385) * $signed(input_fmap_3[15:0]) +
	( 16'sd 29368) * $signed(input_fmap_4[15:0]) +
	( 14'sd 8016) * $signed(input_fmap_5[15:0]) +
	( 16'sd 32011) * $signed(input_fmap_6[15:0]) +
	( 16'sd 22809) * $signed(input_fmap_7[15:0]) +
	( 15'sd 11177) * $signed(input_fmap_8[15:0]) +
	( 16'sd 16971) * $signed(input_fmap_9[15:0]) +
	( 12'sd 1881) * $signed(input_fmap_10[15:0]) +
	( 16'sd 18844) * $signed(input_fmap_11[15:0]) +
	( 16'sd 21177) * $signed(input_fmap_12[15:0]) +
	( 16'sd 28425) * $signed(input_fmap_13[15:0]) +
	( 14'sd 7657) * $signed(input_fmap_14[15:0]) +
	( 16'sd 27868) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10279) * $signed(input_fmap_16[15:0]) +
	( 12'sd 2000) * $signed(input_fmap_17[15:0]) +
	( 16'sd 17896) * $signed(input_fmap_18[15:0]) +
	( 16'sd 24659) * $signed(input_fmap_19[15:0]) +
	( 16'sd 21678) * $signed(input_fmap_20[15:0]) +
	( 16'sd 29294) * $signed(input_fmap_21[15:0]) +
	( 16'sd 30949) * $signed(input_fmap_22[15:0]) +
	( 15'sd 10230) * $signed(input_fmap_23[15:0]) +
	( 14'sd 5757) * $signed(input_fmap_24[15:0]) +
	( 14'sd 5988) * $signed(input_fmap_25[15:0]) +
	( 15'sd 12855) * $signed(input_fmap_26[15:0]) +
	( 12'sd 1751) * $signed(input_fmap_27[15:0]) +
	( 16'sd 31073) * $signed(input_fmap_28[15:0]) +
	( 14'sd 4632) * $signed(input_fmap_29[15:0]) +
	( 16'sd 23936) * $signed(input_fmap_30[15:0]) +
	( 16'sd 27146) * $signed(input_fmap_31[15:0]) +
	( 16'sd 24154) * $signed(input_fmap_32[15:0]) +
	( 16'sd 31054) * $signed(input_fmap_33[15:0]) +
	( 14'sd 4732) * $signed(input_fmap_34[15:0]) +
	( 15'sd 13536) * $signed(input_fmap_35[15:0]) +
	( 16'sd 21296) * $signed(input_fmap_36[15:0]) +
	( 15'sd 12690) * $signed(input_fmap_37[15:0]) +
	( 14'sd 7463) * $signed(input_fmap_38[15:0]) +
	( 14'sd 5633) * $signed(input_fmap_39[15:0]) +
	( 16'sd 30708) * $signed(input_fmap_40[15:0]) +
	( 16'sd 23489) * $signed(input_fmap_41[15:0]) +
	( 16'sd 18007) * $signed(input_fmap_42[15:0]) +
	( 16'sd 31890) * $signed(input_fmap_43[15:0]) +
	( 11'sd 833) * $signed(input_fmap_44[15:0]) +
	( 15'sd 15611) * $signed(input_fmap_45[15:0]) +
	( 15'sd 11730) * $signed(input_fmap_46[15:0]) +
	( 16'sd 23804) * $signed(input_fmap_47[15:0]) +
	( 16'sd 21722) * $signed(input_fmap_48[15:0]) +
	( 15'sd 14455) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26085) * $signed(input_fmap_50[15:0]) +
	( 16'sd 16802) * $signed(input_fmap_51[15:0]) +
	( 15'sd 8257) * $signed(input_fmap_52[15:0]) +
	( 14'sd 6326) * $signed(input_fmap_53[15:0]) +
	( 15'sd 8472) * $signed(input_fmap_54[15:0]) +
	( 16'sd 23166) * $signed(input_fmap_55[15:0]) +
	( 16'sd 23759) * $signed(input_fmap_56[15:0]) +
	( 15'sd 9956) * $signed(input_fmap_57[15:0]) +
	( 10'sd 450) * $signed(input_fmap_58[15:0]) +
	( 16'sd 18267) * $signed(input_fmap_59[15:0]) +
	( 16'sd 30588) * $signed(input_fmap_60[15:0]) +
	( 15'sd 15829) * $signed(input_fmap_61[15:0]) +
	( 14'sd 7855) * $signed(input_fmap_62[15:0]) +
	( 15'sd 8455) * $signed(input_fmap_63[15:0]) +
	( 16'sd 26985) * $signed(input_fmap_64[15:0]) +
	( 16'sd 26094) * $signed(input_fmap_65[15:0]) +
	( 15'sd 13948) * $signed(input_fmap_66[15:0]) +
	( 16'sd 27605) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26502) * $signed(input_fmap_68[15:0]) +
	( 15'sd 13057) * $signed(input_fmap_69[15:0]) +
	( 14'sd 4346) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11456) * $signed(input_fmap_71[15:0]) +
	( 15'sd 12127) * $signed(input_fmap_72[15:0]) +
	( 7'sd 36) * $signed(input_fmap_73[15:0]) +
	( 12'sd 1521) * $signed(input_fmap_74[15:0]) +
	( 13'sd 2282) * $signed(input_fmap_75[15:0]) +
	( 13'sd 2716) * $signed(input_fmap_76[15:0]) +
	( 16'sd 21118) * $signed(input_fmap_77[15:0]) +
	( 13'sd 3188) * $signed(input_fmap_78[15:0]) +
	( 16'sd 25515) * $signed(input_fmap_79[15:0]) +
	( 13'sd 2896) * $signed(input_fmap_80[15:0]) +
	( 16'sd 21357) * $signed(input_fmap_81[15:0]) +
	( 14'sd 7962) * $signed(input_fmap_82[15:0]) +
	( 16'sd 22709) * $signed(input_fmap_83[15:0]) +
	( 14'sd 5799) * $signed(input_fmap_84[15:0]) +
	( 15'sd 11143) * $signed(input_fmap_85[15:0]) +
	( 11'sd 825) * $signed(input_fmap_86[15:0]) +
	( 16'sd 16747) * $signed(input_fmap_87[15:0]) +
	( 16'sd 23735) * $signed(input_fmap_88[15:0]) +
	( 16'sd 29088) * $signed(input_fmap_89[15:0]) +
	( 15'sd 11148) * $signed(input_fmap_90[15:0]) +
	( 15'sd 9360) * $signed(input_fmap_91[15:0]) +
	( 13'sd 3629) * $signed(input_fmap_92[15:0]) +
	( 16'sd 30268) * $signed(input_fmap_93[15:0]) +
	( 14'sd 8101) * $signed(input_fmap_94[15:0]) +
	( 16'sd 21469) * $signed(input_fmap_95[15:0]) +
	( 16'sd 18446) * $signed(input_fmap_96[15:0]) +
	( 16'sd 17074) * $signed(input_fmap_97[15:0]) +
	( 16'sd 24937) * $signed(input_fmap_98[15:0]) +
	( 15'sd 8545) * $signed(input_fmap_99[15:0]) +
	( 16'sd 26349) * $signed(input_fmap_100[15:0]) +
	( 14'sd 6424) * $signed(input_fmap_101[15:0]) +
	( 14'sd 4442) * $signed(input_fmap_102[15:0]) +
	( 16'sd 31019) * $signed(input_fmap_103[15:0]) +
	( 12'sd 1818) * $signed(input_fmap_104[15:0]) +
	( 15'sd 15425) * $signed(input_fmap_105[15:0]) +
	( 12'sd 1087) * $signed(input_fmap_106[15:0]) +
	( 16'sd 26772) * $signed(input_fmap_107[15:0]) +
	( 16'sd 23772) * $signed(input_fmap_108[15:0]) +
	( 13'sd 3296) * $signed(input_fmap_109[15:0]) +
	( 16'sd 31201) * $signed(input_fmap_110[15:0]) +
	( 13'sd 4039) * $signed(input_fmap_111[15:0]) +
	( 15'sd 13275) * $signed(input_fmap_112[15:0]) +
	( 16'sd 20303) * $signed(input_fmap_113[15:0]) +
	( 14'sd 4133) * $signed(input_fmap_114[15:0]) +
	( 15'sd 9330) * $signed(input_fmap_115[15:0]) +
	( 16'sd 19923) * $signed(input_fmap_116[15:0]) +
	( 15'sd 12810) * $signed(input_fmap_117[15:0]) +
	( 16'sd 26962) * $signed(input_fmap_118[15:0]) +
	( 15'sd 11631) * $signed(input_fmap_119[15:0]) +
	( 15'sd 8493) * $signed(input_fmap_120[15:0]) +
	( 16'sd 28597) * $signed(input_fmap_121[15:0]) +
	( 16'sd 18933) * $signed(input_fmap_122[15:0]) +
	( 13'sd 3585) * $signed(input_fmap_123[15:0]) +
	( 11'sd 650) * $signed(input_fmap_124[15:0]) +
	( 14'sd 4394) * $signed(input_fmap_125[15:0]) +
	( 15'sd 13266) * $signed(input_fmap_126[15:0]) +
	( 14'sd 6020) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 16'sd 28042) * $signed(input_fmap_0[15:0]) +
	( 13'sd 3728) * $signed(input_fmap_1[15:0]) +
	( 14'sd 5218) * $signed(input_fmap_2[15:0]) +
	( 13'sd 2793) * $signed(input_fmap_3[15:0]) +
	( 16'sd 32064) * $signed(input_fmap_4[15:0]) +
	( 12'sd 1056) * $signed(input_fmap_5[15:0]) +
	( 14'sd 4865) * $signed(input_fmap_6[15:0]) +
	( 16'sd 18526) * $signed(input_fmap_7[15:0]) +
	( 16'sd 25854) * $signed(input_fmap_8[15:0]) +
	( 16'sd 26894) * $signed(input_fmap_9[15:0]) +
	( 15'sd 11026) * $signed(input_fmap_10[15:0]) +
	( 16'sd 23035) * $signed(input_fmap_11[15:0]) +
	( 14'sd 6547) * $signed(input_fmap_12[15:0]) +
	( 16'sd 22445) * $signed(input_fmap_13[15:0]) +
	( 15'sd 15623) * $signed(input_fmap_14[15:0]) +
	( 16'sd 27569) * $signed(input_fmap_15[15:0]) +
	( 15'sd 15920) * $signed(input_fmap_16[15:0]) +
	( 13'sd 3551) * $signed(input_fmap_17[15:0]) +
	( 9'sd 208) * $signed(input_fmap_18[15:0]) +
	( 15'sd 14431) * $signed(input_fmap_19[15:0]) +
	( 15'sd 13847) * $signed(input_fmap_20[15:0]) +
	( 16'sd 19833) * $signed(input_fmap_21[15:0]) +
	( 13'sd 3437) * $signed(input_fmap_22[15:0]) +
	( 15'sd 13584) * $signed(input_fmap_23[15:0]) +
	( 10'sd 386) * $signed(input_fmap_24[15:0]) +
	( 16'sd 29868) * $signed(input_fmap_25[15:0]) +
	( 16'sd 25878) * $signed(input_fmap_26[15:0]) +
	( 15'sd 8362) * $signed(input_fmap_27[15:0]) +
	( 15'sd 8727) * $signed(input_fmap_28[15:0]) +
	( 15'sd 12932) * $signed(input_fmap_29[15:0]) +
	( 15'sd 12495) * $signed(input_fmap_30[15:0]) +
	( 16'sd 24485) * $signed(input_fmap_31[15:0]) +
	( 16'sd 17221) * $signed(input_fmap_32[15:0]) +
	( 14'sd 7132) * $signed(input_fmap_33[15:0]) +
	( 15'sd 9028) * $signed(input_fmap_34[15:0]) +
	( 16'sd 22881) * $signed(input_fmap_35[15:0]) +
	( 16'sd 21596) * $signed(input_fmap_36[15:0]) +
	( 12'sd 1920) * $signed(input_fmap_37[15:0]) +
	( 16'sd 25818) * $signed(input_fmap_38[15:0]) +
	( 16'sd 32520) * $signed(input_fmap_39[15:0]) +
	( 16'sd 21350) * $signed(input_fmap_40[15:0]) +
	( 16'sd 16909) * $signed(input_fmap_41[15:0]) +
	( 16'sd 22734) * $signed(input_fmap_42[15:0]) +
	( 16'sd 31914) * $signed(input_fmap_43[15:0]) +
	( 16'sd 17782) * $signed(input_fmap_44[15:0]) +
	( 12'sd 1410) * $signed(input_fmap_45[15:0]) +
	( 16'sd 21164) * $signed(input_fmap_46[15:0]) +
	( 16'sd 32732) * $signed(input_fmap_47[15:0]) +
	( 16'sd 23400) * $signed(input_fmap_48[15:0]) +
	( 15'sd 11577) * $signed(input_fmap_49[15:0]) +
	( 16'sd 20574) * $signed(input_fmap_50[15:0]) +
	( 15'sd 11660) * $signed(input_fmap_51[15:0]) +
	( 15'sd 12904) * $signed(input_fmap_52[15:0]) +
	( 15'sd 13574) * $signed(input_fmap_53[15:0]) +
	( 16'sd 19909) * $signed(input_fmap_54[15:0]) +
	( 16'sd 21012) * $signed(input_fmap_55[15:0]) +
	( 14'sd 4285) * $signed(input_fmap_56[15:0]) +
	( 16'sd 17378) * $signed(input_fmap_57[15:0]) +
	( 15'sd 14948) * $signed(input_fmap_58[15:0]) +
	( 10'sd 342) * $signed(input_fmap_59[15:0]) +
	( 14'sd 5450) * $signed(input_fmap_60[15:0]) +
	( 16'sd 16423) * $signed(input_fmap_61[15:0]) +
	( 16'sd 30670) * $signed(input_fmap_62[15:0]) +
	( 11'sd 1010) * $signed(input_fmap_63[15:0]) +
	( 16'sd 26891) * $signed(input_fmap_64[15:0]) +
	( 16'sd 24185) * $signed(input_fmap_65[15:0]) +
	( 16'sd 27114) * $signed(input_fmap_66[15:0]) +
	( 16'sd 28212) * $signed(input_fmap_67[15:0]) +
	( 14'sd 5535) * $signed(input_fmap_68[15:0]) +
	( 14'sd 4415) * $signed(input_fmap_69[15:0]) +
	( 16'sd 17533) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31828) * $signed(input_fmap_71[15:0]) +
	( 16'sd 18938) * $signed(input_fmap_72[15:0]) +
	( 13'sd 3072) * $signed(input_fmap_73[15:0]) +
	( 16'sd 32695) * $signed(input_fmap_74[15:0]) +
	( 15'sd 10148) * $signed(input_fmap_75[15:0]) +
	( 15'sd 16372) * $signed(input_fmap_76[15:0]) +
	( 16'sd 24598) * $signed(input_fmap_77[15:0]) +
	( 16'sd 31203) * $signed(input_fmap_78[15:0]) +
	( 15'sd 13087) * $signed(input_fmap_79[15:0]) +
	( 15'sd 9319) * $signed(input_fmap_80[15:0]) +
	( 16'sd 19646) * $signed(input_fmap_81[15:0]) +
	( 11'sd 610) * $signed(input_fmap_82[15:0]) +
	( 13'sd 2189) * $signed(input_fmap_83[15:0]) +
	( 13'sd 3706) * $signed(input_fmap_84[15:0]) +
	( 16'sd 27885) * $signed(input_fmap_85[15:0]) +
	( 16'sd 30087) * $signed(input_fmap_86[15:0]) +
	( 14'sd 7738) * $signed(input_fmap_87[15:0]) +
	( 16'sd 28872) * $signed(input_fmap_88[15:0]) +
	( 13'sd 3492) * $signed(input_fmap_89[15:0]) +
	( 15'sd 16291) * $signed(input_fmap_90[15:0]) +
	( 15'sd 13799) * $signed(input_fmap_91[15:0]) +
	( 15'sd 16090) * $signed(input_fmap_92[15:0]) +
	( 15'sd 15169) * $signed(input_fmap_93[15:0]) +
	( 16'sd 30179) * $signed(input_fmap_94[15:0]) +
	( 16'sd 23054) * $signed(input_fmap_95[15:0]) +
	( 14'sd 5546) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27422) * $signed(input_fmap_97[15:0]) +
	( 14'sd 5470) * $signed(input_fmap_98[15:0]) +
	( 14'sd 7583) * $signed(input_fmap_99[15:0]) +
	( 11'sd 636) * $signed(input_fmap_100[15:0]) +
	( 16'sd 32379) * $signed(input_fmap_101[15:0]) +
	( 11'sd 601) * $signed(input_fmap_102[15:0]) +
	( 16'sd 29688) * $signed(input_fmap_103[15:0]) +
	( 16'sd 20276) * $signed(input_fmap_104[15:0]) +
	( 16'sd 21125) * $signed(input_fmap_105[15:0]) +
	( 14'sd 8038) * $signed(input_fmap_106[15:0]) +
	( 12'sd 1397) * $signed(input_fmap_107[15:0]) +
	( 16'sd 17080) * $signed(input_fmap_108[15:0]) +
	( 16'sd 24350) * $signed(input_fmap_109[15:0]) +
	( 16'sd 21687) * $signed(input_fmap_110[15:0]) +
	( 16'sd 24810) * $signed(input_fmap_111[15:0]) +
	( 16'sd 29322) * $signed(input_fmap_112[15:0]) +
	( 14'sd 7475) * $signed(input_fmap_113[15:0]) +
	( 10'sd 401) * $signed(input_fmap_114[15:0]) +
	( 16'sd 21643) * $signed(input_fmap_115[15:0]) +
	( 16'sd 18798) * $signed(input_fmap_116[15:0]) +
	( 15'sd 8790) * $signed(input_fmap_117[15:0]) +
	( 13'sd 3435) * $signed(input_fmap_118[15:0]) +
	( 15'sd 10079) * $signed(input_fmap_119[15:0]) +
	( 16'sd 32621) * $signed(input_fmap_120[15:0]) +
	( 15'sd 10794) * $signed(input_fmap_121[15:0]) +
	( 15'sd 16100) * $signed(input_fmap_122[15:0]) +
	( 16'sd 22653) * $signed(input_fmap_123[15:0]) +
	( 15'sd 13159) * $signed(input_fmap_124[15:0]) +
	( 16'sd 19948) * $signed(input_fmap_125[15:0]) +
	( 14'sd 5642) * $signed(input_fmap_126[15:0]) +
	( 16'sd 29979) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 16'sd 30588) * $signed(input_fmap_0[15:0]) +
	( 13'sd 3779) * $signed(input_fmap_1[15:0]) +
	( 15'sd 15182) * $signed(input_fmap_2[15:0]) +
	( 16'sd 17332) * $signed(input_fmap_3[15:0]) +
	( 15'sd 8345) * $signed(input_fmap_4[15:0]) +
	( 16'sd 26884) * $signed(input_fmap_5[15:0]) +
	( 15'sd 8551) * $signed(input_fmap_6[15:0]) +
	( 15'sd 11255) * $signed(input_fmap_7[15:0]) +
	( 16'sd 21299) * $signed(input_fmap_8[15:0]) +
	( 15'sd 10953) * $signed(input_fmap_9[15:0]) +
	( 15'sd 11321) * $signed(input_fmap_10[15:0]) +
	( 16'sd 24851) * $signed(input_fmap_11[15:0]) +
	( 16'sd 30639) * $signed(input_fmap_12[15:0]) +
	( 15'sd 9423) * $signed(input_fmap_13[15:0]) +
	( 16'sd 16439) * $signed(input_fmap_14[15:0]) +
	( 16'sd 30372) * $signed(input_fmap_15[15:0]) +
	( 15'sd 13694) * $signed(input_fmap_16[15:0]) +
	( 15'sd 12140) * $signed(input_fmap_17[15:0]) +
	( 16'sd 19929) * $signed(input_fmap_18[15:0]) +
	( 16'sd 20842) * $signed(input_fmap_19[15:0]) +
	( 15'sd 15652) * $signed(input_fmap_20[15:0]) +
	( 16'sd 20816) * $signed(input_fmap_21[15:0]) +
	( 16'sd 28428) * $signed(input_fmap_22[15:0]) +
	( 16'sd 30131) * $signed(input_fmap_23[15:0]) +
	( 16'sd 22005) * $signed(input_fmap_24[15:0]) +
	( 16'sd 17854) * $signed(input_fmap_25[15:0]) +
	( 16'sd 26490) * $signed(input_fmap_26[15:0]) +
	( 13'sd 2249) * $signed(input_fmap_27[15:0]) +
	( 16'sd 25496) * $signed(input_fmap_28[15:0]) +
	( 16'sd 22790) * $signed(input_fmap_29[15:0]) +
	( 15'sd 12572) * $signed(input_fmap_30[15:0]) +
	( 16'sd 19567) * $signed(input_fmap_31[15:0]) +
	( 15'sd 10901) * $signed(input_fmap_32[15:0]) +
	( 16'sd 27500) * $signed(input_fmap_33[15:0]) +
	( 16'sd 26506) * $signed(input_fmap_34[15:0]) +
	( 16'sd 21228) * $signed(input_fmap_35[15:0]) +
	( 15'sd 12765) * $signed(input_fmap_36[15:0]) +
	( 15'sd 9704) * $signed(input_fmap_37[15:0]) +
	( 16'sd 31984) * $signed(input_fmap_38[15:0]) +
	( 14'sd 4534) * $signed(input_fmap_39[15:0]) +
	( 12'sd 2019) * $signed(input_fmap_40[15:0]) +
	( 16'sd 17828) * $signed(input_fmap_41[15:0]) +
	( 14'sd 5991) * $signed(input_fmap_42[15:0]) +
	( 12'sd 1139) * $signed(input_fmap_43[15:0]) +
	( 15'sd 12702) * $signed(input_fmap_44[15:0]) +
	( 16'sd 31671) * $signed(input_fmap_45[15:0]) +
	( 16'sd 31460) * $signed(input_fmap_46[15:0]) +
	( 16'sd 26761) * $signed(input_fmap_47[15:0]) +
	( 16'sd 20253) * $signed(input_fmap_48[15:0]) +
	( 16'sd 24979) * $signed(input_fmap_49[15:0]) +
	( 16'sd 26244) * $signed(input_fmap_50[15:0]) +
	( 16'sd 18268) * $signed(input_fmap_51[15:0]) +
	( 16'sd 29544) * $signed(input_fmap_52[15:0]) +
	( 16'sd 31379) * $signed(input_fmap_53[15:0]) +
	( 15'sd 12703) * $signed(input_fmap_54[15:0]) +
	( 11'sd 982) * $signed(input_fmap_55[15:0]) +
	( 16'sd 29147) * $signed(input_fmap_56[15:0]) +
	( 16'sd 30692) * $signed(input_fmap_57[15:0]) +
	( 16'sd 27367) * $signed(input_fmap_58[15:0]) +
	( 16'sd 25799) * $signed(input_fmap_59[15:0]) +
	( 12'sd 1405) * $signed(input_fmap_60[15:0]) +
	( 16'sd 27518) * $signed(input_fmap_61[15:0]) +
	( 16'sd 25321) * $signed(input_fmap_62[15:0]) +
	( 14'sd 4504) * $signed(input_fmap_63[15:0]) +
	( 16'sd 28792) * $signed(input_fmap_64[15:0]) +
	( 15'sd 9032) * $signed(input_fmap_65[15:0]) +
	( 12'sd 1819) * $signed(input_fmap_66[15:0]) +
	( 15'sd 12150) * $signed(input_fmap_67[15:0]) +
	( 16'sd 16878) * $signed(input_fmap_68[15:0]) +
	( 15'sd 11777) * $signed(input_fmap_69[15:0]) +
	( 16'sd 20192) * $signed(input_fmap_70[15:0]) +
	( 15'sd 9243) * $signed(input_fmap_71[15:0]) +
	( 16'sd 23399) * $signed(input_fmap_72[15:0]) +
	( 15'sd 14280) * $signed(input_fmap_73[15:0]) +
	( 14'sd 6018) * $signed(input_fmap_74[15:0]) +
	( 16'sd 23671) * $signed(input_fmap_75[15:0]) +
	( 14'sd 7670) * $signed(input_fmap_76[15:0]) +
	( 16'sd 27127) * $signed(input_fmap_77[15:0]) +
	( 16'sd 23274) * $signed(input_fmap_78[15:0]) +
	( 16'sd 24861) * $signed(input_fmap_79[15:0]) +
	( 10'sd 336) * $signed(input_fmap_80[15:0]) +
	( 16'sd 25165) * $signed(input_fmap_81[15:0]) +
	( 16'sd 16657) * $signed(input_fmap_82[15:0]) +
	( 16'sd 17129) * $signed(input_fmap_83[15:0]) +
	( 11'sd 520) * $signed(input_fmap_84[15:0]) +
	( 16'sd 26782) * $signed(input_fmap_85[15:0]) +
	( 12'sd 1839) * $signed(input_fmap_86[15:0]) +
	( 15'sd 15574) * $signed(input_fmap_87[15:0]) +
	( 15'sd 13359) * $signed(input_fmap_88[15:0]) +
	( 16'sd 17395) * $signed(input_fmap_89[15:0]) +
	( 15'sd 15571) * $signed(input_fmap_90[15:0]) +
	( 16'sd 26337) * $signed(input_fmap_91[15:0]) +
	( 16'sd 29231) * $signed(input_fmap_92[15:0]) +
	( 14'sd 4306) * $signed(input_fmap_93[15:0]) +
	( 16'sd 31301) * $signed(input_fmap_94[15:0]) +
	( 14'sd 5962) * $signed(input_fmap_95[15:0]) +
	( 15'sd 8203) * $signed(input_fmap_96[15:0]) +
	( 15'sd 12752) * $signed(input_fmap_97[15:0]) +
	( 14'sd 4114) * $signed(input_fmap_98[15:0]) +
	( 16'sd 29193) * $signed(input_fmap_99[15:0]) +
	( 16'sd 22372) * $signed(input_fmap_100[15:0]) +
	( 15'sd 16277) * $signed(input_fmap_101[15:0]) +
	( 14'sd 6034) * $signed(input_fmap_102[15:0]) +
	( 16'sd 16591) * $signed(input_fmap_103[15:0]) +
	( 15'sd 12647) * $signed(input_fmap_104[15:0]) +
	( 14'sd 5879) * $signed(input_fmap_105[15:0]) +
	( 16'sd 25431) * $signed(input_fmap_106[15:0]) +
	( 15'sd 12839) * $signed(input_fmap_107[15:0]) +
	( 15'sd 14188) * $signed(input_fmap_108[15:0]) +
	( 14'sd 4983) * $signed(input_fmap_109[15:0]) +
	( 15'sd 15230) * $signed(input_fmap_110[15:0]) +
	( 16'sd 23256) * $signed(input_fmap_111[15:0]) +
	( 16'sd 27576) * $signed(input_fmap_112[15:0]) +
	( 14'sd 5438) * $signed(input_fmap_113[15:0]) +
	( 10'sd 263) * $signed(input_fmap_114[15:0]) +
	( 16'sd 22207) * $signed(input_fmap_115[15:0]) +
	( 14'sd 5710) * $signed(input_fmap_116[15:0]) +
	( 16'sd 22756) * $signed(input_fmap_117[15:0]) +
	( 15'sd 11338) * $signed(input_fmap_118[15:0]) +
	( 15'sd 11848) * $signed(input_fmap_119[15:0]) +
	( 16'sd 27163) * $signed(input_fmap_120[15:0]) +
	( 15'sd 16241) * $signed(input_fmap_121[15:0]) +
	( 16'sd 27643) * $signed(input_fmap_122[15:0]) +
	( 16'sd 26425) * $signed(input_fmap_123[15:0]) +
	( 16'sd 32233) * $signed(input_fmap_124[15:0]) +
	( 12'sd 1386) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6001) * $signed(input_fmap_126[15:0]) +
	( 15'sd 11632) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 13'sd 2149) * $signed(input_fmap_0[15:0]) +
	( 15'sd 10169) * $signed(input_fmap_1[15:0]) +
	( 14'sd 6137) * $signed(input_fmap_2[15:0]) +
	( 16'sd 17559) * $signed(input_fmap_3[15:0]) +
	( 16'sd 31539) * $signed(input_fmap_4[15:0]) +
	( 15'sd 9605) * $signed(input_fmap_5[15:0]) +
	( 11'sd 820) * $signed(input_fmap_6[15:0]) +
	( 16'sd 21852) * $signed(input_fmap_7[15:0]) +
	( 14'sd 4749) * $signed(input_fmap_8[15:0]) +
	( 16'sd 18809) * $signed(input_fmap_9[15:0]) +
	( 16'sd 32168) * $signed(input_fmap_10[15:0]) +
	( 16'sd 32516) * $signed(input_fmap_11[15:0]) +
	( 10'sd 394) * $signed(input_fmap_12[15:0]) +
	( 15'sd 11121) * $signed(input_fmap_13[15:0]) +
	( 15'sd 15609) * $signed(input_fmap_14[15:0]) +
	( 14'sd 7395) * $signed(input_fmap_15[15:0]) +
	( 15'sd 8939) * $signed(input_fmap_16[15:0]) +
	( 14'sd 4488) * $signed(input_fmap_17[15:0]) +
	( 16'sd 17332) * $signed(input_fmap_18[15:0]) +
	( 15'sd 12507) * $signed(input_fmap_19[15:0]) +
	( 16'sd 17378) * $signed(input_fmap_20[15:0]) +
	( 16'sd 26855) * $signed(input_fmap_21[15:0]) +
	( 14'sd 8105) * $signed(input_fmap_22[15:0]) +
	( 16'sd 31624) * $signed(input_fmap_23[15:0]) +
	( 14'sd 7937) * $signed(input_fmap_24[15:0]) +
	( 16'sd 23616) * $signed(input_fmap_25[15:0]) +
	( 15'sd 15198) * $signed(input_fmap_26[15:0]) +
	( 14'sd 7497) * $signed(input_fmap_27[15:0]) +
	( 16'sd 24018) * $signed(input_fmap_28[15:0]) +
	( 15'sd 15354) * $signed(input_fmap_29[15:0]) +
	( 16'sd 27494) * $signed(input_fmap_30[15:0]) +
	( 16'sd 23630) * $signed(input_fmap_31[15:0]) +
	( 16'sd 25368) * $signed(input_fmap_32[15:0]) +
	( 16'sd 20660) * $signed(input_fmap_33[15:0]) +
	( 16'sd 19740) * $signed(input_fmap_34[15:0]) +
	( 16'sd 26268) * $signed(input_fmap_35[15:0]) +
	( 16'sd 18931) * $signed(input_fmap_36[15:0]) +
	( 15'sd 11363) * $signed(input_fmap_37[15:0]) +
	( 15'sd 14941) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24720) * $signed(input_fmap_39[15:0]) +
	( 15'sd 13223) * $signed(input_fmap_40[15:0]) +
	( 12'sd 1899) * $signed(input_fmap_41[15:0]) +
	( 15'sd 11975) * $signed(input_fmap_42[15:0]) +
	( 15'sd 11452) * $signed(input_fmap_43[15:0]) +
	( 16'sd 22731) * $signed(input_fmap_44[15:0]) +
	( 16'sd 31070) * $signed(input_fmap_45[15:0]) +
	( 16'sd 17161) * $signed(input_fmap_46[15:0]) +
	( 15'sd 9416) * $signed(input_fmap_47[15:0]) +
	( 16'sd 32652) * $signed(input_fmap_48[15:0]) +
	( 15'sd 12848) * $signed(input_fmap_49[15:0]) +
	( 16'sd 20023) * $signed(input_fmap_50[15:0]) +
	( 15'sd 14333) * $signed(input_fmap_51[15:0]) +
	( 15'sd 11038) * $signed(input_fmap_52[15:0]) +
	( 14'sd 6118) * $signed(input_fmap_53[15:0]) +
	( 11'sd 797) * $signed(input_fmap_54[15:0]) +
	( 15'sd 13609) * $signed(input_fmap_55[15:0]) +
	( 14'sd 4693) * $signed(input_fmap_56[15:0]) +
	( 16'sd 24801) * $signed(input_fmap_57[15:0]) +
	( 15'sd 12201) * $signed(input_fmap_58[15:0]) +
	( 14'sd 7022) * $signed(input_fmap_59[15:0]) +
	( 15'sd 13288) * $signed(input_fmap_60[15:0]) +
	( 14'sd 5317) * $signed(input_fmap_61[15:0]) +
	( 16'sd 22901) * $signed(input_fmap_62[15:0]) +
	( 16'sd 19838) * $signed(input_fmap_63[15:0]) +
	( 14'sd 5361) * $signed(input_fmap_64[15:0]) +
	( 16'sd 21744) * $signed(input_fmap_65[15:0]) +
	( 15'sd 15939) * $signed(input_fmap_66[15:0]) +
	( 16'sd 30807) * $signed(input_fmap_67[15:0]) +
	( 16'sd 21895) * $signed(input_fmap_68[15:0]) +
	( 16'sd 28933) * $signed(input_fmap_69[15:0]) +
	( 16'sd 25987) * $signed(input_fmap_70[15:0]) +
	( 14'sd 4510) * $signed(input_fmap_71[15:0]) +
	( 14'sd 7347) * $signed(input_fmap_72[15:0]) +
	( 16'sd 20613) * $signed(input_fmap_73[15:0]) +
	( 15'sd 9410) * $signed(input_fmap_74[15:0]) +
	( 15'sd 15798) * $signed(input_fmap_75[15:0]) +
	( 16'sd 30923) * $signed(input_fmap_76[15:0]) +
	( 13'sd 2576) * $signed(input_fmap_77[15:0]) +
	( 15'sd 13667) * $signed(input_fmap_78[15:0]) +
	( 14'sd 4475) * $signed(input_fmap_79[15:0]) +
	( 11'sd 621) * $signed(input_fmap_80[15:0]) +
	( 16'sd 29135) * $signed(input_fmap_81[15:0]) +
	( 15'sd 14334) * $signed(input_fmap_82[15:0]) +
	( 16'sd 29228) * $signed(input_fmap_83[15:0]) +
	( 15'sd 13757) * $signed(input_fmap_84[15:0]) +
	( 16'sd 19673) * $signed(input_fmap_85[15:0]) +
	( 14'sd 6110) * $signed(input_fmap_86[15:0]) +
	( 15'sd 15362) * $signed(input_fmap_87[15:0]) +
	( 16'sd 20727) * $signed(input_fmap_88[15:0]) +
	( 16'sd 17750) * $signed(input_fmap_89[15:0]) +
	( 12'sd 1483) * $signed(input_fmap_90[15:0]) +
	( 16'sd 20613) * $signed(input_fmap_91[15:0]) +
	( 16'sd 29702) * $signed(input_fmap_92[15:0]) +
	( 15'sd 13103) * $signed(input_fmap_93[15:0]) +
	( 16'sd 30079) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25642) * $signed(input_fmap_95[15:0]) +
	( 13'sd 2724) * $signed(input_fmap_96[15:0]) +
	( 12'sd 1915) * $signed(input_fmap_97[15:0]) +
	( 14'sd 4425) * $signed(input_fmap_98[15:0]) +
	( 15'sd 12122) * $signed(input_fmap_99[15:0]) +
	( 16'sd 26245) * $signed(input_fmap_100[15:0]) +
	( 15'sd 12317) * $signed(input_fmap_101[15:0]) +
	( 13'sd 3341) * $signed(input_fmap_102[15:0]) +
	( 16'sd 20955) * $signed(input_fmap_103[15:0]) +
	( 16'sd 24185) * $signed(input_fmap_104[15:0]) +
	( 14'sd 4168) * $signed(input_fmap_105[15:0]) +
	( 16'sd 18559) * $signed(input_fmap_106[15:0]) +
	( 15'sd 11731) * $signed(input_fmap_107[15:0]) +
	( 12'sd 1600) * $signed(input_fmap_108[15:0]) +
	( 14'sd 6966) * $signed(input_fmap_109[15:0]) +
	( 16'sd 23392) * $signed(input_fmap_110[15:0]) +
	( 14'sd 6953) * $signed(input_fmap_111[15:0]) +
	( 16'sd 27803) * $signed(input_fmap_112[15:0]) +
	( 16'sd 20916) * $signed(input_fmap_113[15:0]) +
	( 16'sd 18046) * $signed(input_fmap_114[15:0]) +
	( 16'sd 24639) * $signed(input_fmap_115[15:0]) +
	( 15'sd 14010) * $signed(input_fmap_116[15:0]) +
	( 15'sd 14599) * $signed(input_fmap_117[15:0]) +
	( 15'sd 11027) * $signed(input_fmap_118[15:0]) +
	( 16'sd 27384) * $signed(input_fmap_119[15:0]) +
	( 15'sd 11180) * $signed(input_fmap_120[15:0]) +
	( 12'sd 1943) * $signed(input_fmap_121[15:0]) +
	( 15'sd 8889) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21499) * $signed(input_fmap_123[15:0]) +
	( 16'sd 30096) * $signed(input_fmap_124[15:0]) +
	( 13'sd 3437) * $signed(input_fmap_125[15:0]) +
	( 15'sd 8779) * $signed(input_fmap_126[15:0]) +
	( 16'sd 22296) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 15'sd 14550) * $signed(input_fmap_0[15:0]) +
	( 15'sd 8737) * $signed(input_fmap_1[15:0]) +
	( 15'sd 9829) * $signed(input_fmap_2[15:0]) +
	( 15'sd 15793) * $signed(input_fmap_3[15:0]) +
	( 15'sd 8281) * $signed(input_fmap_4[15:0]) +
	( 15'sd 12255) * $signed(input_fmap_5[15:0]) +
	( 16'sd 27146) * $signed(input_fmap_6[15:0]) +
	( 16'sd 23583) * $signed(input_fmap_7[15:0]) +
	( 15'sd 11957) * $signed(input_fmap_8[15:0]) +
	( 12'sd 1636) * $signed(input_fmap_9[15:0]) +
	( 15'sd 11339) * $signed(input_fmap_10[15:0]) +
	( 11'sd 1018) * $signed(input_fmap_11[15:0]) +
	( 14'sd 6587) * $signed(input_fmap_12[15:0]) +
	( 14'sd 5270) * $signed(input_fmap_13[15:0]) +
	( 15'sd 11411) * $signed(input_fmap_14[15:0]) +
	( 16'sd 20879) * $signed(input_fmap_15[15:0]) +
	( 15'sd 10473) * $signed(input_fmap_16[15:0]) +
	( 14'sd 7194) * $signed(input_fmap_17[15:0]) +
	( 16'sd 26200) * $signed(input_fmap_18[15:0]) +
	( 16'sd 24066) * $signed(input_fmap_19[15:0]) +
	( 16'sd 30056) * $signed(input_fmap_20[15:0]) +
	( 16'sd 19442) * $signed(input_fmap_21[15:0]) +
	( 16'sd 30469) * $signed(input_fmap_22[15:0]) +
	( 15'sd 10475) * $signed(input_fmap_23[15:0]) +
	( 15'sd 13170) * $signed(input_fmap_24[15:0]) +
	( 15'sd 9457) * $signed(input_fmap_25[15:0]) +
	( 16'sd 26673) * $signed(input_fmap_26[15:0]) +
	( 16'sd 29018) * $signed(input_fmap_27[15:0]) +
	( 15'sd 14796) * $signed(input_fmap_28[15:0]) +
	( 16'sd 16959) * $signed(input_fmap_29[15:0]) +
	( 14'sd 5938) * $signed(input_fmap_30[15:0]) +
	( 16'sd 29372) * $signed(input_fmap_31[15:0]) +
	( 16'sd 32345) * $signed(input_fmap_32[15:0]) +
	( 13'sd 4015) * $signed(input_fmap_33[15:0]) +
	( 15'sd 15755) * $signed(input_fmap_34[15:0]) +
	( 16'sd 26742) * $signed(input_fmap_35[15:0]) +
	( 16'sd 24086) * $signed(input_fmap_36[15:0]) +
	( 16'sd 27238) * $signed(input_fmap_37[15:0]) +
	( 14'sd 4753) * $signed(input_fmap_38[15:0]) +
	( 16'sd 30082) * $signed(input_fmap_39[15:0]) +
	( 16'sd 24879) * $signed(input_fmap_40[15:0]) +
	( 16'sd 25017) * $signed(input_fmap_41[15:0]) +
	( 16'sd 27595) * $signed(input_fmap_42[15:0]) +
	( 15'sd 10598) * $signed(input_fmap_43[15:0]) +
	( 16'sd 21151) * $signed(input_fmap_44[15:0]) +
	( 12'sd 1444) * $signed(input_fmap_45[15:0]) +
	( 15'sd 13781) * $signed(input_fmap_46[15:0]) +
	( 16'sd 26340) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13266) * $signed(input_fmap_48[15:0]) +
	( 15'sd 10890) * $signed(input_fmap_49[15:0]) +
	( 14'sd 6617) * $signed(input_fmap_50[15:0]) +
	( 15'sd 10779) * $signed(input_fmap_51[15:0]) +
	( 16'sd 16648) * $signed(input_fmap_52[15:0]) +
	( 16'sd 25725) * $signed(input_fmap_53[15:0]) +
	( 15'sd 11258) * $signed(input_fmap_54[15:0]) +
	( 15'sd 9839) * $signed(input_fmap_55[15:0]) +
	( 16'sd 29241) * $signed(input_fmap_56[15:0]) +
	( 15'sd 11336) * $signed(input_fmap_57[15:0]) +
	( 14'sd 7493) * $signed(input_fmap_58[15:0]) +
	( 16'sd 17248) * $signed(input_fmap_59[15:0]) +
	( 13'sd 2983) * $signed(input_fmap_60[15:0]) +
	( 14'sd 7288) * $signed(input_fmap_61[15:0]) +
	( 16'sd 32646) * $signed(input_fmap_62[15:0]) +
	( 14'sd 6525) * $signed(input_fmap_63[15:0]) +
	( 15'sd 8383) * $signed(input_fmap_64[15:0]) +
	( 16'sd 28866) * $signed(input_fmap_65[15:0]) +
	( 15'sd 15499) * $signed(input_fmap_66[15:0]) +
	( 12'sd 1896) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26915) * $signed(input_fmap_68[15:0]) +
	( 14'sd 6782) * $signed(input_fmap_69[15:0]) +
	( 15'sd 11097) * $signed(input_fmap_70[15:0]) +
	( 15'sd 11055) * $signed(input_fmap_71[15:0]) +
	( 16'sd 25575) * $signed(input_fmap_72[15:0]) +
	( 16'sd 32030) * $signed(input_fmap_73[15:0]) +
	( 14'sd 7645) * $signed(input_fmap_74[15:0]) +
	( 16'sd 30464) * $signed(input_fmap_75[15:0]) +
	( 12'sd 2005) * $signed(input_fmap_76[15:0]) +
	( 16'sd 16827) * $signed(input_fmap_77[15:0]) +
	( 15'sd 16360) * $signed(input_fmap_78[15:0]) +
	( 14'sd 7929) * $signed(input_fmap_79[15:0]) +
	( 15'sd 10592) * $signed(input_fmap_80[15:0]) +
	( 16'sd 17140) * $signed(input_fmap_81[15:0]) +
	( 16'sd 25768) * $signed(input_fmap_82[15:0]) +
	( 15'sd 13677) * $signed(input_fmap_83[15:0]) +
	( 13'sd 2629) * $signed(input_fmap_84[15:0]) +
	( 13'sd 2068) * $signed(input_fmap_85[15:0]) +
	( 16'sd 23304) * $signed(input_fmap_86[15:0]) +
	( 14'sd 5034) * $signed(input_fmap_87[15:0]) +
	( 15'sd 10785) * $signed(input_fmap_88[15:0]) +
	( 15'sd 10824) * $signed(input_fmap_89[15:0]) +
	( 15'sd 10194) * $signed(input_fmap_90[15:0]) +
	( 15'sd 14168) * $signed(input_fmap_91[15:0]) +
	( 16'sd 30583) * $signed(input_fmap_92[15:0]) +
	( 16'sd 23595) * $signed(input_fmap_93[15:0]) +
	( 16'sd 26182) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25269) * $signed(input_fmap_95[15:0]) +
	( 16'sd 16751) * $signed(input_fmap_96[15:0]) +
	( 15'sd 10135) * $signed(input_fmap_97[15:0]) +
	( 16'sd 23941) * $signed(input_fmap_98[15:0]) +
	( 16'sd 17141) * $signed(input_fmap_99[15:0]) +
	( 13'sd 2096) * $signed(input_fmap_100[15:0]) +
	( 16'sd 27567) * $signed(input_fmap_101[15:0]) +
	( 16'sd 31105) * $signed(input_fmap_102[15:0]) +
	( 14'sd 5681) * $signed(input_fmap_103[15:0]) +
	( 16'sd 30897) * $signed(input_fmap_104[15:0]) +
	( 16'sd 27332) * $signed(input_fmap_105[15:0]) +
	( 15'sd 12529) * $signed(input_fmap_106[15:0]) +
	( 15'sd 10737) * $signed(input_fmap_107[15:0]) +
	( 16'sd 29616) * $signed(input_fmap_108[15:0]) +
	( 16'sd 30408) * $signed(input_fmap_109[15:0]) +
	( 16'sd 26043) * $signed(input_fmap_110[15:0]) +
	( 16'sd 21427) * $signed(input_fmap_111[15:0]) +
	( 16'sd 19590) * $signed(input_fmap_112[15:0]) +
	( 15'sd 9000) * $signed(input_fmap_113[15:0]) +
	( 16'sd 30488) * $signed(input_fmap_114[15:0]) +
	( 16'sd 21593) * $signed(input_fmap_115[15:0]) +
	( 16'sd 26569) * $signed(input_fmap_116[15:0]) +
	( 16'sd 18802) * $signed(input_fmap_117[15:0]) +
	( 15'sd 13384) * $signed(input_fmap_118[15:0]) +
	( 16'sd 27525) * $signed(input_fmap_119[15:0]) +
	( 15'sd 13919) * $signed(input_fmap_120[15:0]) +
	( 16'sd 26096) * $signed(input_fmap_121[15:0]) +
	( 16'sd 17819) * $signed(input_fmap_122[15:0]) +
	( 16'sd 23982) * $signed(input_fmap_123[15:0]) +
	( 16'sd 21633) * $signed(input_fmap_124[15:0]) +
	( 16'sd 19681) * $signed(input_fmap_125[15:0]) +
	( 14'sd 6255) * $signed(input_fmap_126[15:0]) +
	( 16'sd 26210) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 16'sd 28572) * $signed(input_fmap_0[15:0]) +
	( 15'sd 14616) * $signed(input_fmap_1[15:0]) +
	( 16'sd 27779) * $signed(input_fmap_2[15:0]) +
	( 12'sd 1971) * $signed(input_fmap_3[15:0]) +
	( 16'sd 29119) * $signed(input_fmap_4[15:0]) +
	( 16'sd 24829) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2899) * $signed(input_fmap_6[15:0]) +
	( 14'sd 5848) * $signed(input_fmap_7[15:0]) +
	( 16'sd 24902) * $signed(input_fmap_8[15:0]) +
	( 13'sd 3519) * $signed(input_fmap_9[15:0]) +
	( 16'sd 26960) * $signed(input_fmap_10[15:0]) +
	( 15'sd 8328) * $signed(input_fmap_11[15:0]) +
	( 16'sd 22182) * $signed(input_fmap_12[15:0]) +
	( 15'sd 9649) * $signed(input_fmap_13[15:0]) +
	( 15'sd 13590) * $signed(input_fmap_14[15:0]) +
	( 16'sd 30056) * $signed(input_fmap_15[15:0]) +
	( 16'sd 21556) * $signed(input_fmap_16[15:0]) +
	( 16'sd 30495) * $signed(input_fmap_17[15:0]) +
	( 13'sd 3677) * $signed(input_fmap_18[15:0]) +
	( 15'sd 8331) * $signed(input_fmap_19[15:0]) +
	( 14'sd 6199) * $signed(input_fmap_20[15:0]) +
	( 15'sd 13927) * $signed(input_fmap_21[15:0]) +
	( 16'sd 31578) * $signed(input_fmap_22[15:0]) +
	( 15'sd 10764) * $signed(input_fmap_23[15:0]) +
	( 16'sd 16455) * $signed(input_fmap_24[15:0]) +
	( 16'sd 30815) * $signed(input_fmap_25[15:0]) +
	( 15'sd 11032) * $signed(input_fmap_26[15:0]) +
	( 14'sd 5698) * $signed(input_fmap_27[15:0]) +
	( 14'sd 8104) * $signed(input_fmap_28[15:0]) +
	( 15'sd 8754) * $signed(input_fmap_29[15:0]) +
	( 16'sd 31334) * $signed(input_fmap_30[15:0]) +
	( 16'sd 16400) * $signed(input_fmap_31[15:0]) +
	( 16'sd 23189) * $signed(input_fmap_32[15:0]) +
	( 12'sd 1028) * $signed(input_fmap_33[15:0]) +
	( 16'sd 26728) * $signed(input_fmap_34[15:0]) +
	( 13'sd 3955) * $signed(input_fmap_35[15:0]) +
	( 16'sd 31926) * $signed(input_fmap_36[15:0]) +
	( 15'sd 12918) * $signed(input_fmap_37[15:0]) +
	( 15'sd 9670) * $signed(input_fmap_38[15:0]) +
	( 8'sd 104) * $signed(input_fmap_39[15:0]) +
	( 15'sd 11733) * $signed(input_fmap_40[15:0]) +
	( 15'sd 13909) * $signed(input_fmap_41[15:0]) +
	( 16'sd 28421) * $signed(input_fmap_42[15:0]) +
	( 16'sd 25196) * $signed(input_fmap_43[15:0]) +
	( 15'sd 14386) * $signed(input_fmap_44[15:0]) +
	( 16'sd 31990) * $signed(input_fmap_45[15:0]) +
	( 14'sd 5230) * $signed(input_fmap_46[15:0]) +
	( 13'sd 2507) * $signed(input_fmap_47[15:0]) +
	( 14'sd 4356) * $signed(input_fmap_48[15:0]) +
	( 16'sd 17451) * $signed(input_fmap_49[15:0]) +
	( 15'sd 11082) * $signed(input_fmap_50[15:0]) +
	( 16'sd 30281) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19307) * $signed(input_fmap_52[15:0]) +
	( 16'sd 29479) * $signed(input_fmap_53[15:0]) +
	( 16'sd 17680) * $signed(input_fmap_54[15:0]) +
	( 16'sd 19859) * $signed(input_fmap_55[15:0]) +
	( 16'sd 16879) * $signed(input_fmap_56[15:0]) +
	( 14'sd 8152) * $signed(input_fmap_57[15:0]) +
	( 14'sd 4600) * $signed(input_fmap_58[15:0]) +
	( 16'sd 29467) * $signed(input_fmap_59[15:0]) +
	( 16'sd 18302) * $signed(input_fmap_60[15:0]) +
	( 16'sd 30632) * $signed(input_fmap_61[15:0]) +
	( 15'sd 8248) * $signed(input_fmap_62[15:0]) +
	( 16'sd 27708) * $signed(input_fmap_63[15:0]) +
	( 14'sd 5498) * $signed(input_fmap_64[15:0]) +
	( 16'sd 24070) * $signed(input_fmap_65[15:0]) +
	( 16'sd 30437) * $signed(input_fmap_66[15:0]) +
	( 13'sd 3173) * $signed(input_fmap_67[15:0]) +
	( 13'sd 2229) * $signed(input_fmap_68[15:0]) +
	( 15'sd 15781) * $signed(input_fmap_69[15:0]) +
	( 16'sd 27847) * $signed(input_fmap_70[15:0]) +
	( 16'sd 26453) * $signed(input_fmap_71[15:0]) +
	( 16'sd 19347) * $signed(input_fmap_72[15:0]) +
	( 14'sd 4921) * $signed(input_fmap_73[15:0]) +
	( 16'sd 26711) * $signed(input_fmap_74[15:0]) +
	( 16'sd 20802) * $signed(input_fmap_75[15:0]) +
	( 16'sd 29518) * $signed(input_fmap_76[15:0]) +
	( 16'sd 27288) * $signed(input_fmap_77[15:0]) +
	( 14'sd 4833) * $signed(input_fmap_78[15:0]) +
	( 15'sd 12477) * $signed(input_fmap_79[15:0]) +
	( 14'sd 6765) * $signed(input_fmap_80[15:0]) +
	( 16'sd 22114) * $signed(input_fmap_81[15:0]) +
	( 14'sd 6380) * $signed(input_fmap_82[15:0]) +
	( 16'sd 26375) * $signed(input_fmap_83[15:0]) +
	( 13'sd 4091) * $signed(input_fmap_84[15:0]) +
	( 15'sd 11960) * $signed(input_fmap_85[15:0]) +
	( 15'sd 15575) * $signed(input_fmap_86[15:0]) +
	( 12'sd 1264) * $signed(input_fmap_87[15:0]) +
	( 15'sd 10400) * $signed(input_fmap_88[15:0]) +
	( 13'sd 3332) * $signed(input_fmap_89[15:0]) +
	( 15'sd 15335) * $signed(input_fmap_90[15:0]) +
	( 16'sd 23220) * $signed(input_fmap_91[15:0]) +
	( 16'sd 31277) * $signed(input_fmap_92[15:0]) +
	( 16'sd 21847) * $signed(input_fmap_93[15:0]) +
	( 15'sd 15960) * $signed(input_fmap_94[15:0]) +
	( 16'sd 29261) * $signed(input_fmap_95[15:0]) +
	( 16'sd 30902) * $signed(input_fmap_96[15:0]) +
	( 16'sd 18133) * $signed(input_fmap_97[15:0]) +
	( 13'sd 2787) * $signed(input_fmap_98[15:0]) +
	( 13'sd 3853) * $signed(input_fmap_99[15:0]) +
	( 16'sd 26161) * $signed(input_fmap_100[15:0]) +
	( 16'sd 25151) * $signed(input_fmap_101[15:0]) +
	( 16'sd 19410) * $signed(input_fmap_102[15:0]) +
	( 15'sd 15216) * $signed(input_fmap_103[15:0]) +
	( 15'sd 13154) * $signed(input_fmap_104[15:0]) +
	( 11'sd 1000) * $signed(input_fmap_105[15:0]) +
	( 16'sd 20906) * $signed(input_fmap_106[15:0]) +
	( 15'sd 15413) * $signed(input_fmap_107[15:0]) +
	( 16'sd 16696) * $signed(input_fmap_108[15:0]) +
	( 13'sd 3477) * $signed(input_fmap_109[15:0]) +
	( 14'sd 8157) * $signed(input_fmap_110[15:0]) +
	( 15'sd 14483) * $signed(input_fmap_111[15:0]) +
	( 14'sd 8001) * $signed(input_fmap_112[15:0]) +
	( 16'sd 31730) * $signed(input_fmap_113[15:0]) +
	( 15'sd 13833) * $signed(input_fmap_114[15:0]) +
	( 16'sd 28939) * $signed(input_fmap_115[15:0]) +
	( 16'sd 24060) * $signed(input_fmap_116[15:0]) +
	( 16'sd 21802) * $signed(input_fmap_117[15:0]) +
	( 16'sd 18567) * $signed(input_fmap_118[15:0]) +
	( 14'sd 6856) * $signed(input_fmap_119[15:0]) +
	( 16'sd 23200) * $signed(input_fmap_120[15:0]) +
	( 12'sd 1959) * $signed(input_fmap_121[15:0]) +
	( 16'sd 32701) * $signed(input_fmap_122[15:0]) +
	( 11'sd 583) * $signed(input_fmap_123[15:0]) +
	( 12'sd 1688) * $signed(input_fmap_124[15:0]) +
	( 12'sd 1754) * $signed(input_fmap_125[15:0]) +
	( 14'sd 4299) * $signed(input_fmap_126[15:0]) +
	( 10'sd 452) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 16'sd 21305) * $signed(input_fmap_0[15:0]) +
	( 13'sd 3658) * $signed(input_fmap_1[15:0]) +
	( 16'sd 16810) * $signed(input_fmap_2[15:0]) +
	( 14'sd 7367) * $signed(input_fmap_3[15:0]) +
	( 15'sd 9223) * $signed(input_fmap_4[15:0]) +
	( 15'sd 11713) * $signed(input_fmap_5[15:0]) +
	( 15'sd 10153) * $signed(input_fmap_6[15:0]) +
	( 16'sd 23557) * $signed(input_fmap_7[15:0]) +
	( 16'sd 22786) * $signed(input_fmap_8[15:0]) +
	( 15'sd 8207) * $signed(input_fmap_9[15:0]) +
	( 16'sd 19581) * $signed(input_fmap_10[15:0]) +
	( 15'sd 15103) * $signed(input_fmap_11[15:0]) +
	( 16'sd 26209) * $signed(input_fmap_12[15:0]) +
	( 16'sd 30380) * $signed(input_fmap_13[15:0]) +
	( 15'sd 13203) * $signed(input_fmap_14[15:0]) +
	( 16'sd 20804) * $signed(input_fmap_15[15:0]) +
	( 16'sd 24457) * $signed(input_fmap_16[15:0]) +
	( 15'sd 14744) * $signed(input_fmap_17[15:0]) +
	( 16'sd 18531) * $signed(input_fmap_18[15:0]) +
	( 16'sd 23207) * $signed(input_fmap_19[15:0]) +
	( 13'sd 2661) * $signed(input_fmap_20[15:0]) +
	( 15'sd 13495) * $signed(input_fmap_21[15:0]) +
	( 16'sd 31175) * $signed(input_fmap_22[15:0]) +
	( 16'sd 27383) * $signed(input_fmap_23[15:0]) +
	( 15'sd 15397) * $signed(input_fmap_24[15:0]) +
	( 16'sd 16561) * $signed(input_fmap_25[15:0]) +
	( 15'sd 15779) * $signed(input_fmap_26[15:0]) +
	( 9'sd 191) * $signed(input_fmap_27[15:0]) +
	( 11'sd 954) * $signed(input_fmap_28[15:0]) +
	( 16'sd 19138) * $signed(input_fmap_29[15:0]) +
	( 16'sd 21784) * $signed(input_fmap_30[15:0]) +
	( 16'sd 30432) * $signed(input_fmap_31[15:0]) +
	( 14'sd 4567) * $signed(input_fmap_32[15:0]) +
	( 16'sd 26497) * $signed(input_fmap_33[15:0]) +
	( 16'sd 16961) * $signed(input_fmap_34[15:0]) +
	( 15'sd 12797) * $signed(input_fmap_35[15:0]) +
	( 15'sd 9272) * $signed(input_fmap_36[15:0]) +
	( 16'sd 19494) * $signed(input_fmap_37[15:0]) +
	( 16'sd 19977) * $signed(input_fmap_38[15:0]) +
	( 16'sd 31950) * $signed(input_fmap_39[15:0]) +
	( 15'sd 12452) * $signed(input_fmap_40[15:0]) +
	( 16'sd 22986) * $signed(input_fmap_41[15:0]) +
	( 16'sd 26431) * $signed(input_fmap_42[15:0]) +
	( 16'sd 17351) * $signed(input_fmap_43[15:0]) +
	( 16'sd 22299) * $signed(input_fmap_44[15:0]) +
	( 14'sd 5770) * $signed(input_fmap_45[15:0]) +
	( 16'sd 17749) * $signed(input_fmap_46[15:0]) +
	( 16'sd 22352) * $signed(input_fmap_47[15:0]) +
	( 16'sd 28935) * $signed(input_fmap_48[15:0]) +
	( 15'sd 10377) * $signed(input_fmap_49[15:0]) +
	( 15'sd 9814) * $signed(input_fmap_50[15:0]) +
	( 13'sd 3081) * $signed(input_fmap_51[15:0]) +
	( 16'sd 29975) * $signed(input_fmap_52[15:0]) +
	( 16'sd 29401) * $signed(input_fmap_53[15:0]) +
	( 15'sd 13455) * $signed(input_fmap_54[15:0]) +
	( 16'sd 21474) * $signed(input_fmap_55[15:0]) +
	( 13'sd 3645) * $signed(input_fmap_56[15:0]) +
	( 16'sd 30699) * $signed(input_fmap_57[15:0]) +
	( 15'sd 15263) * $signed(input_fmap_58[15:0]) +
	( 16'sd 27382) * $signed(input_fmap_59[15:0]) +
	( 15'sd 8721) * $signed(input_fmap_60[15:0]) +
	( 16'sd 26796) * $signed(input_fmap_61[15:0]) +
	( 16'sd 31445) * $signed(input_fmap_62[15:0]) +
	( 16'sd 24405) * $signed(input_fmap_63[15:0]) +
	( 16'sd 24156) * $signed(input_fmap_64[15:0]) +
	( 15'sd 16143) * $signed(input_fmap_65[15:0]) +
	( 16'sd 28844) * $signed(input_fmap_66[15:0]) +
	( 16'sd 21690) * $signed(input_fmap_67[15:0]) +
	( 16'sd 26242) * $signed(input_fmap_68[15:0]) +
	( 16'sd 29557) * $signed(input_fmap_69[15:0]) +
	( 15'sd 13129) * $signed(input_fmap_70[15:0]) +
	( 14'sd 4259) * $signed(input_fmap_71[15:0]) +
	( 4'sd 5) * $signed(input_fmap_72[15:0]) +
	( 16'sd 26689) * $signed(input_fmap_73[15:0]) +
	( 14'sd 4911) * $signed(input_fmap_74[15:0]) +
	( 15'sd 14190) * $signed(input_fmap_75[15:0]) +
	( 16'sd 30138) * $signed(input_fmap_76[15:0]) +
	( 15'sd 14095) * $signed(input_fmap_77[15:0]) +
	( 16'sd 26307) * $signed(input_fmap_78[15:0]) +
	( 16'sd 20423) * $signed(input_fmap_79[15:0]) +
	( 14'sd 4491) * $signed(input_fmap_80[15:0]) +
	( 14'sd 6881) * $signed(input_fmap_81[15:0]) +
	( 16'sd 26208) * $signed(input_fmap_82[15:0]) +
	( 14'sd 5241) * $signed(input_fmap_83[15:0]) +
	( 15'sd 14565) * $signed(input_fmap_84[15:0]) +
	( 16'sd 17329) * $signed(input_fmap_85[15:0]) +
	( 15'sd 13430) * $signed(input_fmap_86[15:0]) +
	( 15'sd 13505) * $signed(input_fmap_87[15:0]) +
	( 16'sd 25631) * $signed(input_fmap_88[15:0]) +
	( 16'sd 30978) * $signed(input_fmap_89[15:0]) +
	( 14'sd 7180) * $signed(input_fmap_90[15:0]) +
	( 13'sd 2070) * $signed(input_fmap_91[15:0]) +
	( 15'sd 9669) * $signed(input_fmap_92[15:0]) +
	( 15'sd 10614) * $signed(input_fmap_93[15:0]) +
	( 16'sd 25486) * $signed(input_fmap_94[15:0]) +
	( 13'sd 2956) * $signed(input_fmap_95[15:0]) +
	( 16'sd 29573) * $signed(input_fmap_96[15:0]) +
	( 16'sd 31530) * $signed(input_fmap_97[15:0]) +
	( 16'sd 17416) * $signed(input_fmap_98[15:0]) +
	( 15'sd 8314) * $signed(input_fmap_99[15:0]) +
	( 16'sd 31004) * $signed(input_fmap_100[15:0]) +
	( 16'sd 20650) * $signed(input_fmap_101[15:0]) +
	( 16'sd 25218) * $signed(input_fmap_102[15:0]) +
	( 15'sd 14285) * $signed(input_fmap_103[15:0]) +
	( 14'sd 7756) * $signed(input_fmap_104[15:0]) +
	( 16'sd 32766) * $signed(input_fmap_105[15:0]) +
	( 16'sd 18337) * $signed(input_fmap_106[15:0]) +
	( 15'sd 8780) * $signed(input_fmap_107[15:0]) +
	( 16'sd 27355) * $signed(input_fmap_108[15:0]) +
	( 16'sd 18520) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22382) * $signed(input_fmap_110[15:0]) +
	( 16'sd 29747) * $signed(input_fmap_111[15:0]) +
	( 15'sd 14365) * $signed(input_fmap_112[15:0]) +
	( 14'sd 6582) * $signed(input_fmap_113[15:0]) +
	( 15'sd 13419) * $signed(input_fmap_114[15:0]) +
	( 15'sd 13732) * $signed(input_fmap_115[15:0]) +
	( 15'sd 12622) * $signed(input_fmap_116[15:0]) +
	( 16'sd 17672) * $signed(input_fmap_117[15:0]) +
	( 16'sd 22345) * $signed(input_fmap_118[15:0]) +
	( 13'sd 3959) * $signed(input_fmap_119[15:0]) +
	( 16'sd 28302) * $signed(input_fmap_120[15:0]) +
	( 15'sd 15232) * $signed(input_fmap_121[15:0]) +
	( 15'sd 12820) * $signed(input_fmap_122[15:0]) +
	( 16'sd 27211) * $signed(input_fmap_123[15:0]) +
	( 16'sd 28950) * $signed(input_fmap_124[15:0]) +
	( 14'sd 7665) * $signed(input_fmap_125[15:0]) +
	( 16'sd 23910) * $signed(input_fmap_126[15:0]) +
	( 16'sd 27914) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 16'sd 23150) * $signed(input_fmap_0[15:0]) +
	( 16'sd 17837) * $signed(input_fmap_1[15:0]) +
	( 16'sd 27207) * $signed(input_fmap_2[15:0]) +
	( 16'sd 28055) * $signed(input_fmap_3[15:0]) +
	( 16'sd 26793) * $signed(input_fmap_4[15:0]) +
	( 14'sd 5971) * $signed(input_fmap_5[15:0]) +
	( 15'sd 13390) * $signed(input_fmap_6[15:0]) +
	( 15'sd 12436) * $signed(input_fmap_7[15:0]) +
	( 16'sd 23107) * $signed(input_fmap_8[15:0]) +
	( 9'sd 233) * $signed(input_fmap_9[15:0]) +
	( 16'sd 24315) * $signed(input_fmap_10[15:0]) +
	( 11'sd 726) * $signed(input_fmap_11[15:0]) +
	( 16'sd 30773) * $signed(input_fmap_12[15:0]) +
	( 14'sd 6851) * $signed(input_fmap_13[15:0]) +
	( 16'sd 21538) * $signed(input_fmap_14[15:0]) +
	( 15'sd 13342) * $signed(input_fmap_15[15:0]) +
	( 16'sd 18287) * $signed(input_fmap_16[15:0]) +
	( 16'sd 29320) * $signed(input_fmap_17[15:0]) +
	( 13'sd 2206) * $signed(input_fmap_18[15:0]) +
	( 16'sd 18141) * $signed(input_fmap_19[15:0]) +
	( 15'sd 11910) * $signed(input_fmap_20[15:0]) +
	( 16'sd 26198) * $signed(input_fmap_21[15:0]) +
	( 16'sd 22751) * $signed(input_fmap_22[15:0]) +
	( 14'sd 6994) * $signed(input_fmap_23[15:0]) +
	( 16'sd 19510) * $signed(input_fmap_24[15:0]) +
	( 15'sd 15247) * $signed(input_fmap_25[15:0]) +
	( 15'sd 10330) * $signed(input_fmap_26[15:0]) +
	( 13'sd 3534) * $signed(input_fmap_27[15:0]) +
	( 16'sd 25555) * $signed(input_fmap_28[15:0]) +
	( 16'sd 30814) * $signed(input_fmap_29[15:0]) +
	( 16'sd 17749) * $signed(input_fmap_30[15:0]) +
	( 16'sd 26179) * $signed(input_fmap_31[15:0]) +
	( 16'sd 18037) * $signed(input_fmap_32[15:0]) +
	( 15'sd 10097) * $signed(input_fmap_33[15:0]) +
	( 13'sd 3424) * $signed(input_fmap_34[15:0]) +
	( 15'sd 11348) * $signed(input_fmap_35[15:0]) +
	( 16'sd 19650) * $signed(input_fmap_36[15:0]) +
	( 15'sd 12172) * $signed(input_fmap_37[15:0]) +
	( 12'sd 1045) * $signed(input_fmap_38[15:0]) +
	( 16'sd 24772) * $signed(input_fmap_39[15:0]) +
	( 9'sd 251) * $signed(input_fmap_40[15:0]) +
	( 15'sd 9499) * $signed(input_fmap_41[15:0]) +
	( 16'sd 23446) * $signed(input_fmap_42[15:0]) +
	( 14'sd 7600) * $signed(input_fmap_43[15:0]) +
	( 16'sd 20688) * $signed(input_fmap_44[15:0]) +
	( 16'sd 26741) * $signed(input_fmap_45[15:0]) +
	( 14'sd 8130) * $signed(input_fmap_46[15:0]) +
	( 16'sd 17056) * $signed(input_fmap_47[15:0]) +
	( 15'sd 10274) * $signed(input_fmap_48[15:0]) +
	( 15'sd 14363) * $signed(input_fmap_49[15:0]) +
	( 16'sd 22182) * $signed(input_fmap_50[15:0]) +
	( 8'sd 94) * $signed(input_fmap_51[15:0]) +
	( 16'sd 19350) * $signed(input_fmap_52[15:0]) +
	( 12'sd 1892) * $signed(input_fmap_53[15:0]) +
	( 16'sd 20238) * $signed(input_fmap_54[15:0]) +
	( 16'sd 18245) * $signed(input_fmap_55[15:0]) +
	( 16'sd 19057) * $signed(input_fmap_56[15:0]) +
	( 15'sd 11608) * $signed(input_fmap_57[15:0]) +
	( 16'sd 29554) * $signed(input_fmap_58[15:0]) +
	( 12'sd 1565) * $signed(input_fmap_59[15:0]) +
	( 16'sd 28544) * $signed(input_fmap_60[15:0]) +
	( 15'sd 14917) * $signed(input_fmap_61[15:0]) +
	( 16'sd 28728) * $signed(input_fmap_62[15:0]) +
	( 15'sd 14376) * $signed(input_fmap_63[15:0]) +
	( 11'sd 780) * $signed(input_fmap_64[15:0]) +
	( 16'sd 27264) * $signed(input_fmap_65[15:0]) +
	( 16'sd 18031) * $signed(input_fmap_66[15:0]) +
	( 15'sd 12435) * $signed(input_fmap_67[15:0]) +
	( 16'sd 16696) * $signed(input_fmap_68[15:0]) +
	( 16'sd 31095) * $signed(input_fmap_69[15:0]) +
	( 16'sd 23702) * $signed(input_fmap_70[15:0]) +
	( 16'sd 31566) * $signed(input_fmap_71[15:0]) +
	( 15'sd 14006) * $signed(input_fmap_72[15:0]) +
	( 14'sd 7622) * $signed(input_fmap_73[15:0]) +
	( 16'sd 30230) * $signed(input_fmap_74[15:0]) +
	( 16'sd 19595) * $signed(input_fmap_75[15:0]) +
	( 15'sd 8530) * $signed(input_fmap_76[15:0]) +
	( 14'sd 7939) * $signed(input_fmap_77[15:0]) +
	( 16'sd 16580) * $signed(input_fmap_78[15:0]) +
	( 15'sd 15861) * $signed(input_fmap_79[15:0]) +
	( 16'sd 19128) * $signed(input_fmap_80[15:0]) +
	( 16'sd 23242) * $signed(input_fmap_81[15:0]) +
	( 15'sd 9137) * $signed(input_fmap_82[15:0]) +
	( 16'sd 25389) * $signed(input_fmap_83[15:0]) +
	( 15'sd 9420) * $signed(input_fmap_84[15:0]) +
	( 16'sd 25986) * $signed(input_fmap_85[15:0]) +
	( 16'sd 16655) * $signed(input_fmap_86[15:0]) +
	( 16'sd 29783) * $signed(input_fmap_87[15:0]) +
	( 16'sd 30298) * $signed(input_fmap_88[15:0]) +
	( 11'sd 920) * $signed(input_fmap_89[15:0]) +
	( 16'sd 17457) * $signed(input_fmap_90[15:0]) +
	( 16'sd 24828) * $signed(input_fmap_91[15:0]) +
	( 16'sd 30417) * $signed(input_fmap_92[15:0]) +
	( 12'sd 1414) * $signed(input_fmap_93[15:0]) +
	( 16'sd 30094) * $signed(input_fmap_94[15:0]) +
	( 14'sd 4170) * $signed(input_fmap_95[15:0]) +
	( 14'sd 7414) * $signed(input_fmap_96[15:0]) +
	( 16'sd 27683) * $signed(input_fmap_97[15:0]) +
	( 15'sd 14260) * $signed(input_fmap_98[15:0]) +
	( 16'sd 24582) * $signed(input_fmap_99[15:0]) +
	( 15'sd 10866) * $signed(input_fmap_100[15:0]) +
	( 14'sd 5567) * $signed(input_fmap_101[15:0]) +
	( 16'sd 32236) * $signed(input_fmap_102[15:0]) +
	( 15'sd 15480) * $signed(input_fmap_103[15:0]) +
	( 16'sd 25689) * $signed(input_fmap_104[15:0]) +
	( 16'sd 30867) * $signed(input_fmap_105[15:0]) +
	( 12'sd 2001) * $signed(input_fmap_106[15:0]) +
	( 16'sd 22872) * $signed(input_fmap_107[15:0]) +
	( 15'sd 15997) * $signed(input_fmap_108[15:0]) +
	( 16'sd 25124) * $signed(input_fmap_109[15:0]) +
	( 16'sd 22710) * $signed(input_fmap_110[15:0]) +
	( 16'sd 20014) * $signed(input_fmap_111[15:0]) +
	( 16'sd 25790) * $signed(input_fmap_112[15:0]) +
	( 16'sd 29272) * $signed(input_fmap_113[15:0]) +
	( 16'sd 26782) * $signed(input_fmap_114[15:0]) +
	( 9'sd 148) * $signed(input_fmap_115[15:0]) +
	( 15'sd 15892) * $signed(input_fmap_116[15:0]) +
	( 16'sd 31446) * $signed(input_fmap_117[15:0]) +
	( 16'sd 18512) * $signed(input_fmap_118[15:0]) +
	( 16'sd 16624) * $signed(input_fmap_119[15:0]) +
	( 16'sd 18068) * $signed(input_fmap_120[15:0]) +
	( 16'sd 27838) * $signed(input_fmap_121[15:0]) +
	( 16'sd 16891) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21653) * $signed(input_fmap_123[15:0]) +
	( 16'sd 23407) * $signed(input_fmap_124[15:0]) +
	( 15'sd 15962) * $signed(input_fmap_125[15:0]) +
	( 15'sd 12886) * $signed(input_fmap_126[15:0]) +
	( 15'sd 13670) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 16'sd 23498) * $signed(input_fmap_0[15:0]) +
	( 15'sd 13591) * $signed(input_fmap_1[15:0]) +
	( 16'sd 22622) * $signed(input_fmap_2[15:0]) +
	( 16'sd 25820) * $signed(input_fmap_3[15:0]) +
	( 16'sd 24181) * $signed(input_fmap_4[15:0]) +
	( 15'sd 11288) * $signed(input_fmap_5[15:0]) +
	( 13'sd 2529) * $signed(input_fmap_6[15:0]) +
	( 12'sd 1151) * $signed(input_fmap_7[15:0]) +
	( 16'sd 16867) * $signed(input_fmap_8[15:0]) +
	( 16'sd 19337) * $signed(input_fmap_9[15:0]) +
	( 16'sd 16688) * $signed(input_fmap_10[15:0]) +
	( 16'sd 25456) * $signed(input_fmap_11[15:0]) +
	( 15'sd 12482) * $signed(input_fmap_12[15:0]) +
	( 13'sd 3875) * $signed(input_fmap_13[15:0]) +
	( 14'sd 5591) * $signed(input_fmap_14[15:0]) +
	( 15'sd 12922) * $signed(input_fmap_15[15:0]) +
	( 16'sd 26221) * $signed(input_fmap_16[15:0]) +
	( 11'sd 669) * $signed(input_fmap_17[15:0]) +
	( 16'sd 19582) * $signed(input_fmap_18[15:0]) +
	( 7'sd 46) * $signed(input_fmap_19[15:0]) +
	( 15'sd 12631) * $signed(input_fmap_20[15:0]) +
	( 16'sd 25067) * $signed(input_fmap_21[15:0]) +
	( 15'sd 14550) * $signed(input_fmap_22[15:0]) +
	( 16'sd 22868) * $signed(input_fmap_23[15:0]) +
	( 16'sd 23669) * $signed(input_fmap_24[15:0]) +
	( 16'sd 28630) * $signed(input_fmap_25[15:0]) +
	( 16'sd 32475) * $signed(input_fmap_26[15:0]) +
	( 15'sd 15401) * $signed(input_fmap_27[15:0]) +
	( 16'sd 29107) * $signed(input_fmap_28[15:0]) +
	( 16'sd 22806) * $signed(input_fmap_29[15:0]) +
	( 14'sd 6421) * $signed(input_fmap_30[15:0]) +
	( 16'sd 24439) * $signed(input_fmap_31[15:0]) +
	( 15'sd 11681) * $signed(input_fmap_32[15:0]) +
	( 16'sd 23643) * $signed(input_fmap_33[15:0]) +
	( 12'sd 1545) * $signed(input_fmap_34[15:0]) +
	( 13'sd 2315) * $signed(input_fmap_35[15:0]) +
	( 13'sd 2256) * $signed(input_fmap_36[15:0]) +
	( 16'sd 20376) * $signed(input_fmap_37[15:0]) +
	( 16'sd 25526) * $signed(input_fmap_38[15:0]) +
	( 15'sd 9372) * $signed(input_fmap_39[15:0]) +
	( 16'sd 19483) * $signed(input_fmap_40[15:0]) +
	( 16'sd 17998) * $signed(input_fmap_41[15:0]) +
	( 15'sd 11031) * $signed(input_fmap_42[15:0]) +
	( 16'sd 17167) * $signed(input_fmap_43[15:0]) +
	( 16'sd 26684) * $signed(input_fmap_44[15:0]) +
	( 16'sd 18758) * $signed(input_fmap_45[15:0]) +
	( 15'sd 13619) * $signed(input_fmap_46[15:0]) +
	( 16'sd 26074) * $signed(input_fmap_47[15:0]) +
	( 16'sd 22389) * $signed(input_fmap_48[15:0]) +
	( 16'sd 23374) * $signed(input_fmap_49[15:0]) +
	( 15'sd 11284) * $signed(input_fmap_50[15:0]) +
	( 14'sd 6225) * $signed(input_fmap_51[15:0]) +
	( 16'sd 28818) * $signed(input_fmap_52[15:0]) +
	( 16'sd 21654) * $signed(input_fmap_53[15:0]) +
	( 16'sd 28404) * $signed(input_fmap_54[15:0]) +
	( 16'sd 18392) * $signed(input_fmap_55[15:0]) +
	( 16'sd 21052) * $signed(input_fmap_56[15:0]) +
	( 14'sd 4107) * $signed(input_fmap_57[15:0]) +
	( 15'sd 9616) * $signed(input_fmap_58[15:0]) +
	( 16'sd 29540) * $signed(input_fmap_59[15:0]) +
	( 16'sd 17825) * $signed(input_fmap_60[15:0]) +
	( 16'sd 22598) * $signed(input_fmap_61[15:0]) +
	( 16'sd 16717) * $signed(input_fmap_62[15:0]) +
	( 15'sd 13822) * $signed(input_fmap_63[15:0]) +
	( 16'sd 26367) * $signed(input_fmap_64[15:0]) +
	( 14'sd 5522) * $signed(input_fmap_65[15:0]) +
	( 16'sd 31255) * $signed(input_fmap_66[15:0]) +
	( 16'sd 22557) * $signed(input_fmap_67[15:0]) +
	( 16'sd 30938) * $signed(input_fmap_68[15:0]) +
	( 16'sd 28775) * $signed(input_fmap_69[15:0]) +
	( 15'sd 11974) * $signed(input_fmap_70[15:0]) +
	( 15'sd 9782) * $signed(input_fmap_71[15:0]) +
	( 16'sd 22612) * $signed(input_fmap_72[15:0]) +
	( 13'sd 2394) * $signed(input_fmap_73[15:0]) +
	( 13'sd 2533) * $signed(input_fmap_74[15:0]) +
	( 13'sd 3961) * $signed(input_fmap_75[15:0]) +
	( 16'sd 26122) * $signed(input_fmap_76[15:0]) +
	( 16'sd 30853) * $signed(input_fmap_77[15:0]) +
	( 14'sd 6780) * $signed(input_fmap_78[15:0]) +
	( 15'sd 14717) * $signed(input_fmap_79[15:0]) +
	( 15'sd 8720) * $signed(input_fmap_80[15:0]) +
	( 13'sd 2587) * $signed(input_fmap_81[15:0]) +
	( 14'sd 4651) * $signed(input_fmap_82[15:0]) +
	( 14'sd 7692) * $signed(input_fmap_83[15:0]) +
	( 16'sd 23329) * $signed(input_fmap_84[15:0]) +
	( 16'sd 25387) * $signed(input_fmap_85[15:0]) +
	( 15'sd 13541) * $signed(input_fmap_86[15:0]) +
	( 16'sd 27739) * $signed(input_fmap_87[15:0]) +
	( 16'sd 31434) * $signed(input_fmap_88[15:0]) +
	( 16'sd 16431) * $signed(input_fmap_89[15:0]) +
	( 14'sd 6431) * $signed(input_fmap_90[15:0]) +
	( 15'sd 11434) * $signed(input_fmap_91[15:0]) +
	( 16'sd 32373) * $signed(input_fmap_92[15:0]) +
	( 15'sd 11487) * $signed(input_fmap_93[15:0]) +
	( 16'sd 19833) * $signed(input_fmap_94[15:0]) +
	( 16'sd 25125) * $signed(input_fmap_95[15:0]) +
	( 16'sd 22217) * $signed(input_fmap_96[15:0]) +
	( 16'sd 25424) * $signed(input_fmap_97[15:0]) +
	( 16'sd 17852) * $signed(input_fmap_98[15:0]) +
	( 14'sd 5750) * $signed(input_fmap_99[15:0]) +
	( 13'sd 3235) * $signed(input_fmap_100[15:0]) +
	( 14'sd 4342) * $signed(input_fmap_101[15:0]) +
	( 16'sd 18584) * $signed(input_fmap_102[15:0]) +
	( 16'sd 31923) * $signed(input_fmap_103[15:0]) +
	( 14'sd 5291) * $signed(input_fmap_104[15:0]) +
	( 14'sd 5648) * $signed(input_fmap_105[15:0]) +
	( 16'sd 29923) * $signed(input_fmap_106[15:0]) +
	( 16'sd 17453) * $signed(input_fmap_107[15:0]) +
	( 16'sd 22449) * $signed(input_fmap_108[15:0]) +
	( 16'sd 30117) * $signed(input_fmap_109[15:0]) +
	( 15'sd 13336) * $signed(input_fmap_110[15:0]) +
	( 15'sd 11857) * $signed(input_fmap_111[15:0]) +
	( 16'sd 26261) * $signed(input_fmap_112[15:0]) +
	( 15'sd 12183) * $signed(input_fmap_113[15:0]) +
	( 14'sd 6828) * $signed(input_fmap_114[15:0]) +
	( 16'sd 24006) * $signed(input_fmap_115[15:0]) +
	( 14'sd 7030) * $signed(input_fmap_116[15:0]) +
	( 15'sd 13070) * $signed(input_fmap_117[15:0]) +
	( 16'sd 31787) * $signed(input_fmap_118[15:0]) +
	( 15'sd 14718) * $signed(input_fmap_119[15:0]) +
	( 16'sd 29209) * $signed(input_fmap_120[15:0]) +
	( 16'sd 25597) * $signed(input_fmap_121[15:0]) +
	( 16'sd 23965) * $signed(input_fmap_122[15:0]) +
	( 16'sd 21066) * $signed(input_fmap_123[15:0]) +
	( 16'sd 21373) * $signed(input_fmap_124[15:0]) +
	( 16'sd 24847) * $signed(input_fmap_125[15:0]) +
	( 14'sd 4920) * $signed(input_fmap_126[15:0]) +
	( 16'sd 24653) * $signed(input_fmap_127[15:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 16'sd 19950) * $signed(input_fmap_0[15:0]) +
	( 14'sd 4549) * $signed(input_fmap_1[15:0]) +
	( 14'sd 5562) * $signed(input_fmap_2[15:0]) +
	( 14'sd 5153) * $signed(input_fmap_3[15:0]) +
	( 16'sd 22672) * $signed(input_fmap_4[15:0]) +
	( 15'sd 14387) * $signed(input_fmap_5[15:0]) +
	( 15'sd 10626) * $signed(input_fmap_6[15:0]) +
	( 16'sd 31177) * $signed(input_fmap_7[15:0]) +
	( 16'sd 30962) * $signed(input_fmap_8[15:0]) +
	( 15'sd 10625) * $signed(input_fmap_9[15:0]) +
	( 16'sd 32379) * $signed(input_fmap_10[15:0]) +
	( 15'sd 15735) * $signed(input_fmap_11[15:0]) +
	( 15'sd 10129) * $signed(input_fmap_12[15:0]) +
	( 16'sd 29296) * $signed(input_fmap_13[15:0]) +
	( 16'sd 27484) * $signed(input_fmap_14[15:0]) +
	( 16'sd 32221) * $signed(input_fmap_15[15:0]) +
	( 16'sd 19424) * $signed(input_fmap_16[15:0]) +
	( 16'sd 19885) * $signed(input_fmap_17[15:0]) +
	( 16'sd 24605) * $signed(input_fmap_18[15:0]) +
	( 16'sd 17971) * $signed(input_fmap_19[15:0]) +
	( 16'sd 19636) * $signed(input_fmap_20[15:0]) +
	( 15'sd 8521) * $signed(input_fmap_21[15:0]) +
	( 15'sd 8735) * $signed(input_fmap_22[15:0]) +
	( 16'sd 25208) * $signed(input_fmap_23[15:0]) +
	( 12'sd 1756) * $signed(input_fmap_24[15:0]) +
	( 16'sd 19412) * $signed(input_fmap_25[15:0]) +
	( 15'sd 11433) * $signed(input_fmap_26[15:0]) +
	( 16'sd 25998) * $signed(input_fmap_27[15:0]) +
	( 14'sd 6239) * $signed(input_fmap_28[15:0]) +
	( 16'sd 17736) * $signed(input_fmap_29[15:0]) +
	( 16'sd 25689) * $signed(input_fmap_30[15:0]) +
	( 16'sd 17700) * $signed(input_fmap_31[15:0]) +
	( 15'sd 14888) * $signed(input_fmap_32[15:0]) +
	( 16'sd 18507) * $signed(input_fmap_33[15:0]) +
	( 15'sd 9006) * $signed(input_fmap_34[15:0]) +
	( 16'sd 24209) * $signed(input_fmap_35[15:0]) +
	( 16'sd 26225) * $signed(input_fmap_36[15:0]) +
	( 16'sd 27027) * $signed(input_fmap_37[15:0]) +
	( 16'sd 28594) * $signed(input_fmap_38[15:0]) +
	( 15'sd 15719) * $signed(input_fmap_39[15:0]) +
	( 16'sd 19161) * $signed(input_fmap_40[15:0]) +
	( 15'sd 11088) * $signed(input_fmap_41[15:0]) +
	( 16'sd 20419) * $signed(input_fmap_42[15:0]) +
	( 16'sd 32738) * $signed(input_fmap_43[15:0]) +
	( 16'sd 30831) * $signed(input_fmap_44[15:0]) +
	( 16'sd 26675) * $signed(input_fmap_45[15:0]) +
	( 16'sd 28379) * $signed(input_fmap_46[15:0]) +
	( 11'sd 688) * $signed(input_fmap_47[15:0]) +
	( 15'sd 13912) * $signed(input_fmap_48[15:0]) +
	( 9'sd 143) * $signed(input_fmap_49[15:0]) +
	( 16'sd 20573) * $signed(input_fmap_50[15:0]) +
	( 15'sd 14324) * $signed(input_fmap_51[15:0]) +
	( 16'sd 21220) * $signed(input_fmap_52[15:0]) +
	( 16'sd 20667) * $signed(input_fmap_53[15:0]) +
	( 15'sd 12380) * $signed(input_fmap_54[15:0]) +
	( 15'sd 13284) * $signed(input_fmap_55[15:0]) +
	( 16'sd 32489) * $signed(input_fmap_56[15:0]) +
	( 16'sd 27158) * $signed(input_fmap_57[15:0]) +
	( 16'sd 29696) * $signed(input_fmap_58[15:0]) +
	( 16'sd 28420) * $signed(input_fmap_59[15:0]) +
	( 16'sd 20342) * $signed(input_fmap_60[15:0]) +
	( 15'sd 12691) * $signed(input_fmap_61[15:0]) +
	( 16'sd 18698) * $signed(input_fmap_62[15:0]) +
	( 15'sd 14794) * $signed(input_fmap_63[15:0]) +
	( 16'sd 21739) * $signed(input_fmap_64[15:0]) +
	( 16'sd 19758) * $signed(input_fmap_65[15:0]) +
	( 16'sd 25598) * $signed(input_fmap_66[15:0]) +
	( 16'sd 32379) * $signed(input_fmap_67[15:0]) +
	( 16'sd 30340) * $signed(input_fmap_68[15:0]) +
	( 15'sd 15357) * $signed(input_fmap_69[15:0]) +
	( 16'sd 30444) * $signed(input_fmap_70[15:0]) +
	( 15'sd 13066) * $signed(input_fmap_71[15:0]) +
	( 14'sd 5770) * $signed(input_fmap_72[15:0]) +
	( 15'sd 9802) * $signed(input_fmap_73[15:0]) +
	( 16'sd 19858) * $signed(input_fmap_74[15:0]) +
	( 16'sd 27668) * $signed(input_fmap_75[15:0]) +
	( 15'sd 10790) * $signed(input_fmap_76[15:0]) +
	( 15'sd 11423) * $signed(input_fmap_77[15:0]) +
	( 15'sd 16262) * $signed(input_fmap_78[15:0]) +
	( 13'sd 2672) * $signed(input_fmap_79[15:0]) +
	( 16'sd 16577) * $signed(input_fmap_80[15:0]) +
	( 13'sd 2489) * $signed(input_fmap_81[15:0]) +
	( 16'sd 26343) * $signed(input_fmap_82[15:0]) +
	( 15'sd 8514) * $signed(input_fmap_83[15:0]) +
	( 14'sd 5896) * $signed(input_fmap_84[15:0]) +
	( 10'sd 279) * $signed(input_fmap_85[15:0]) +
	( 13'sd 2079) * $signed(input_fmap_86[15:0]) +
	( 16'sd 30606) * $signed(input_fmap_87[15:0]) +
	( 15'sd 12652) * $signed(input_fmap_88[15:0]) +
	( 14'sd 5558) * $signed(input_fmap_89[15:0]) +
	( 15'sd 13996) * $signed(input_fmap_90[15:0]) +
	( 13'sd 2982) * $signed(input_fmap_91[15:0]) +
	( 14'sd 7466) * $signed(input_fmap_92[15:0]) +
	( 16'sd 26284) * $signed(input_fmap_93[15:0]) +
	( 13'sd 2489) * $signed(input_fmap_94[15:0]) +
	( 16'sd 18603) * $signed(input_fmap_95[15:0]) +
	( 16'sd 22151) * $signed(input_fmap_96[15:0]) +
	( 16'sd 17713) * $signed(input_fmap_97[15:0]) +
	( 16'sd 28112) * $signed(input_fmap_98[15:0]) +
	( 15'sd 14287) * $signed(input_fmap_99[15:0]) +
	( 16'sd 17347) * $signed(input_fmap_100[15:0]) +
	( 16'sd 27243) * $signed(input_fmap_101[15:0]) +
	( 15'sd 11294) * $signed(input_fmap_102[15:0]) +
	( 15'sd 8826) * $signed(input_fmap_103[15:0]) +
	( 15'sd 14315) * $signed(input_fmap_104[15:0]) +
	( 15'sd 9679) * $signed(input_fmap_105[15:0]) +
	( 16'sd 26921) * $signed(input_fmap_106[15:0]) +
	( 8'sd 76) * $signed(input_fmap_107[15:0]) +
	( 12'sd 1786) * $signed(input_fmap_108[15:0]) +
	( 15'sd 12070) * $signed(input_fmap_109[15:0]) +
	( 16'sd 23075) * $signed(input_fmap_110[15:0]) +
	( 15'sd 11895) * $signed(input_fmap_111[15:0]) +
	( 15'sd 12091) * $signed(input_fmap_112[15:0]) +
	( 16'sd 26632) * $signed(input_fmap_113[15:0]) +
	( 16'sd 31031) * $signed(input_fmap_114[15:0]) +
	( 15'sd 14876) * $signed(input_fmap_115[15:0]) +
	( 16'sd 23733) * $signed(input_fmap_116[15:0]) +
	( 16'sd 27729) * $signed(input_fmap_117[15:0]) +
	( 16'sd 26131) * $signed(input_fmap_118[15:0]) +
	( 16'sd 18914) * $signed(input_fmap_119[15:0]) +
	( 13'sd 2878) * $signed(input_fmap_120[15:0]) +
	( 15'sd 13688) * $signed(input_fmap_121[15:0]) +
	( 14'sd 4630) * $signed(input_fmap_122[15:0]) +
	( 16'sd 24737) * $signed(input_fmap_123[15:0]) +
	( 16'sd 25828) * $signed(input_fmap_124[15:0]) +
	( 15'sd 10173) * $signed(input_fmap_125[15:0]) +
	( 15'sd 11083) * $signed(input_fmap_126[15:0]) +
	( 16'sd 29374) * $signed(input_fmap_127[15:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 16'd27712;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 16'd18066;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 15'd13774;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 15'd12566;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 12'd1318;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 16'd19624;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 12'd1068;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 10'd355;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 15'd9122;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 16'd22721;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 16'd24781;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 10'd438;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 13'd2687;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 14'd5094;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 15'd11100;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 16'd17215;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 12'd1560;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 16'd27114;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 15'd10068;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 16'd30263;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 16'd25331;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 4'd7;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 16'd29162;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 15'd14436;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 15'd8706;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 16'd20294;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 11'd808;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 12'd1760;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 16'd20222;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 16'd20768;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 11'd675;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 16'd30298;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 16'd25482;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 16'd19389;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 16'd28916;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 16'd20881;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 16'd20547;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 14'd7135;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 16'd20548;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 15'd12623;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 15'd10827;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 16'd17558;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 16'd32691;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 15'd8840;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 14'd4209;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 16'd16912;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 15'd9625;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 16'd23036;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 16'd27663;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 15'd16061;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 16'd20302;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 15'd11849;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 15'd12239;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 16'd21962;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 13'd3866;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 13'd2765;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 14'd5148;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 15'd13195;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 16'd27621;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 14'd4395;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 16'd21446;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 16'd16452;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 12'd1151;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 15'd11739;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64 + 16'd20421;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 15'd9830;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 14'd5431;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67 + 14'd4986;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 16'd26111;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 14'd6037;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 14'd7367;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 16'd23491;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 16'd28885;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 16'd18178;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74 + 15'd11112;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 11'd649;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 15'd16255;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 15'd15895;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 16'd29834;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79 + 15'd11230;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80 + 16'd26354;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81 + 14'd8050;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 16'd26807;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 16'd25214;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 15'd15864;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 12'd1211;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 16'd25522;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 16'd17351;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 16'd29073;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 16'd27686;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 16'd30432;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91 + 15'd15851;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 15'd15124;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 15'd14066;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 16'd30727;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 16'd26852;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 13'd2761;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97 + 15'd11867;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 13'd3930;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 15'd13494;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 16'd18486;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 16'd19502;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102 + 13'd2445;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 14'd7942;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 16'd29572;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 15'd8940;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 16'd19100;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 15'd8796;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108 + 15'd14844;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 16'd26205;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 16'd26240;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 16'd19180;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 16'd29249;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113 + 5'd12;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 13'd2544;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 16'd19033;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116 + 12'd1820;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117 + 16'd20530;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 16'd25782;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 16'd18665;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 16'd24082;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 16'd22849;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 16'd23464;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 16'd30365;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124 + 15'd11203;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 14'd4653;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 16'd31996;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 16'd18431;

logic [15:0] relu_0;
assign relu_0[15:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[29:15]}} :'d6) : '0;
logic [15:0] relu_1;
assign relu_1[15:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[29:15]}} :'d6) : '0;
logic [15:0] relu_2;
assign relu_2[15:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[29:15]}} :'d6) : '0;
logic [15:0] relu_3;
assign relu_3[15:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[29:15]}} :'d6) : '0;
logic [15:0] relu_4;
assign relu_4[15:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[29:15]}} :'d6) : '0;
logic [15:0] relu_5;
assign relu_5[15:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[29:15]}} :'d6) : '0;
logic [15:0] relu_6;
assign relu_6[15:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[29:15]}} :'d6) : '0;
logic [15:0] relu_7;
assign relu_7[15:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[29:15]}} :'d6) : '0;
logic [15:0] relu_8;
assign relu_8[15:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[29:15]}} :'d6) : '0;
logic [15:0] relu_9;
assign relu_9[15:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[29:15]}} :'d6) : '0;
logic [15:0] relu_10;
assign relu_10[15:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[29:15]}} :'d6) : '0;
logic [15:0] relu_11;
assign relu_11[15:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[29:15]}} :'d6) : '0;
logic [15:0] relu_12;
assign relu_12[15:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[29:15]}} :'d6) : '0;
logic [15:0] relu_13;
assign relu_13[15:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[29:15]}} :'d6) : '0;
logic [15:0] relu_14;
assign relu_14[15:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[29:15]}} :'d6) : '0;
logic [15:0] relu_15;
assign relu_15[15:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[29:15]}} :'d6) : '0;
logic [15:0] relu_16;
assign relu_16[15:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[29:15]}} :'d6) : '0;
logic [15:0] relu_17;
assign relu_17[15:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[29:15]}} :'d6) : '0;
logic [15:0] relu_18;
assign relu_18[15:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[29:15]}} :'d6) : '0;
logic [15:0] relu_19;
assign relu_19[15:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[29:15]}} :'d6) : '0;
logic [15:0] relu_20;
assign relu_20[15:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[29:15]}} :'d6) : '0;
logic [15:0] relu_21;
assign relu_21[15:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[29:15]}} :'d6) : '0;
logic [15:0] relu_22;
assign relu_22[15:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[29:15]}} :'d6) : '0;
logic [15:0] relu_23;
assign relu_23[15:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[29:15]}} :'d6) : '0;
logic [15:0] relu_24;
assign relu_24[15:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[29:15]}} :'d6) : '0;
logic [15:0] relu_25;
assign relu_25[15:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[29:15]}} :'d6) : '0;
logic [15:0] relu_26;
assign relu_26[15:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[29:15]}} :'d6) : '0;
logic [15:0] relu_27;
assign relu_27[15:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[29:15]}} :'d6) : '0;
logic [15:0] relu_28;
assign relu_28[15:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[29:15]}} :'d6) : '0;
logic [15:0] relu_29;
assign relu_29[15:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[29:15]}} :'d6) : '0;
logic [15:0] relu_30;
assign relu_30[15:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[29:15]}} :'d6) : '0;
logic [15:0] relu_31;
assign relu_31[15:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[29:15]}} :'d6) : '0;
logic [15:0] relu_32;
assign relu_32[15:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[29:15]}} :'d6) : '0;
logic [15:0] relu_33;
assign relu_33[15:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[29:15]}} :'d6) : '0;
logic [15:0] relu_34;
assign relu_34[15:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[29:15]}} :'d6) : '0;
logic [15:0] relu_35;
assign relu_35[15:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[29:15]}} :'d6) : '0;
logic [15:0] relu_36;
assign relu_36[15:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[29:15]}} :'d6) : '0;
logic [15:0] relu_37;
assign relu_37[15:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[29:15]}} :'d6) : '0;
logic [15:0] relu_38;
assign relu_38[15:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[29:15]}} :'d6) : '0;
logic [15:0] relu_39;
assign relu_39[15:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[29:15]}} :'d6) : '0;
logic [15:0] relu_40;
assign relu_40[15:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[29:15]}} :'d6) : '0;
logic [15:0] relu_41;
assign relu_41[15:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[29:15]}} :'d6) : '0;
logic [15:0] relu_42;
assign relu_42[15:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[29:15]}} :'d6) : '0;
logic [15:0] relu_43;
assign relu_43[15:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[29:15]}} :'d6) : '0;
logic [15:0] relu_44;
assign relu_44[15:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[29:15]}} :'d6) : '0;
logic [15:0] relu_45;
assign relu_45[15:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[29:15]}} :'d6) : '0;
logic [15:0] relu_46;
assign relu_46[15:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[29:15]}} :'d6) : '0;
logic [15:0] relu_47;
assign relu_47[15:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[29:15]}} :'d6) : '0;
logic [15:0] relu_48;
assign relu_48[15:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[29:15]}} :'d6) : '0;
logic [15:0] relu_49;
assign relu_49[15:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[29:15]}} :'d6) : '0;
logic [15:0] relu_50;
assign relu_50[15:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[29:15]}} :'d6) : '0;
logic [15:0] relu_51;
assign relu_51[15:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[29:15]}} :'d6) : '0;
logic [15:0] relu_52;
assign relu_52[15:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[29:15]}} :'d6) : '0;
logic [15:0] relu_53;
assign relu_53[15:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[29:15]}} :'d6) : '0;
logic [15:0] relu_54;
assign relu_54[15:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[29:15]}} :'d6) : '0;
logic [15:0] relu_55;
assign relu_55[15:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[29:15]}} :'d6) : '0;
logic [15:0] relu_56;
assign relu_56[15:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[29:15]}} :'d6) : '0;
logic [15:0] relu_57;
assign relu_57[15:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[29:15]}} :'d6) : '0;
logic [15:0] relu_58;
assign relu_58[15:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[29:15]}} :'d6) : '0;
logic [15:0] relu_59;
assign relu_59[15:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[29:15]}} :'d6) : '0;
logic [15:0] relu_60;
assign relu_60[15:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[29:15]}} :'d6) : '0;
logic [15:0] relu_61;
assign relu_61[15:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[29:15]}} :'d6) : '0;
logic [15:0] relu_62;
assign relu_62[15:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[29:15]}} :'d6) : '0;
logic [15:0] relu_63;
assign relu_63[15:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[29:15]}} :'d6) : '0;
logic [15:0] relu_64;
assign relu_64[15:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[29:15]}} :'d6) : '0;
logic [15:0] relu_65;
assign relu_65[15:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[29:15]}} :'d6) : '0;
logic [15:0] relu_66;
assign relu_66[15:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[29:15]}} :'d6) : '0;
logic [15:0] relu_67;
assign relu_67[15:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[29:15]}} :'d6) : '0;
logic [15:0] relu_68;
assign relu_68[15:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[29:15]}} :'d6) : '0;
logic [15:0] relu_69;
assign relu_69[15:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[29:15]}} :'d6) : '0;
logic [15:0] relu_70;
assign relu_70[15:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[29:15]}} :'d6) : '0;
logic [15:0] relu_71;
assign relu_71[15:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[29:15]}} :'d6) : '0;
logic [15:0] relu_72;
assign relu_72[15:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[29:15]}} :'d6) : '0;
logic [15:0] relu_73;
assign relu_73[15:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[29:15]}} :'d6) : '0;
logic [15:0] relu_74;
assign relu_74[15:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[29:15]}} :'d6) : '0;
logic [15:0] relu_75;
assign relu_75[15:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[29:15]}} :'d6) : '0;
logic [15:0] relu_76;
assign relu_76[15:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[29:15]}} :'d6) : '0;
logic [15:0] relu_77;
assign relu_77[15:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[29:15]}} :'d6) : '0;
logic [15:0] relu_78;
assign relu_78[15:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[29:15]}} :'d6) : '0;
logic [15:0] relu_79;
assign relu_79[15:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[29:15]}} :'d6) : '0;
logic [15:0] relu_80;
assign relu_80[15:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[29:15]}} :'d6) : '0;
logic [15:0] relu_81;
assign relu_81[15:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[29:15]}} :'d6) : '0;
logic [15:0] relu_82;
assign relu_82[15:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[29:15]}} :'d6) : '0;
logic [15:0] relu_83;
assign relu_83[15:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[29:15]}} :'d6) : '0;
logic [15:0] relu_84;
assign relu_84[15:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[29:15]}} :'d6) : '0;
logic [15:0] relu_85;
assign relu_85[15:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[29:15]}} :'d6) : '0;
logic [15:0] relu_86;
assign relu_86[15:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[29:15]}} :'d6) : '0;
logic [15:0] relu_87;
assign relu_87[15:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[29:15]}} :'d6) : '0;
logic [15:0] relu_88;
assign relu_88[15:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[29:15]}} :'d6) : '0;
logic [15:0] relu_89;
assign relu_89[15:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[29:15]}} :'d6) : '0;
logic [15:0] relu_90;
assign relu_90[15:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[29:15]}} :'d6) : '0;
logic [15:0] relu_91;
assign relu_91[15:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[29:15]}} :'d6) : '0;
logic [15:0] relu_92;
assign relu_92[15:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[29:15]}} :'d6) : '0;
logic [15:0] relu_93;
assign relu_93[15:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[29:15]}} :'d6) : '0;
logic [15:0] relu_94;
assign relu_94[15:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[29:15]}} :'d6) : '0;
logic [15:0] relu_95;
assign relu_95[15:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[29:15]}} :'d6) : '0;
logic [15:0] relu_96;
assign relu_96[15:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[29:15]}} :'d6) : '0;
logic [15:0] relu_97;
assign relu_97[15:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[29:15]}} :'d6) : '0;
logic [15:0] relu_98;
assign relu_98[15:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[29:15]}} :'d6) : '0;
logic [15:0] relu_99;
assign relu_99[15:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[29:15]}} :'d6) : '0;
logic [15:0] relu_100;
assign relu_100[15:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[29:15]}} :'d6) : '0;
logic [15:0] relu_101;
assign relu_101[15:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[29:15]}} :'d6) : '0;
logic [15:0] relu_102;
assign relu_102[15:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[29:15]}} :'d6) : '0;
logic [15:0] relu_103;
assign relu_103[15:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[29:15]}} :'d6) : '0;
logic [15:0] relu_104;
assign relu_104[15:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[29:15]}} :'d6) : '0;
logic [15:0] relu_105;
assign relu_105[15:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[29:15]}} :'d6) : '0;
logic [15:0] relu_106;
assign relu_106[15:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[29:15]}} :'d6) : '0;
logic [15:0] relu_107;
assign relu_107[15:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[29:15]}} :'d6) : '0;
logic [15:0] relu_108;
assign relu_108[15:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[29:15]}} :'d6) : '0;
logic [15:0] relu_109;
assign relu_109[15:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[29:15]}} :'d6) : '0;
logic [15:0] relu_110;
assign relu_110[15:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[29:15]}} :'d6) : '0;
logic [15:0] relu_111;
assign relu_111[15:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[29:15]}} :'d6) : '0;
logic [15:0] relu_112;
assign relu_112[15:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[29:15]}} :'d6) : '0;
logic [15:0] relu_113;
assign relu_113[15:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[29:15]}} :'d6) : '0;
logic [15:0] relu_114;
assign relu_114[15:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[29:15]}} :'d6) : '0;
logic [15:0] relu_115;
assign relu_115[15:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[29:15]}} :'d6) : '0;
logic [15:0] relu_116;
assign relu_116[15:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[29:15]}} :'d6) : '0;
logic [15:0] relu_117;
assign relu_117[15:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[29:15]}} :'d6) : '0;
logic [15:0] relu_118;
assign relu_118[15:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[29:15]}} :'d6) : '0;
logic [15:0] relu_119;
assign relu_119[15:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[29:15]}} :'d6) : '0;
logic [15:0] relu_120;
assign relu_120[15:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[29:15]}} :'d6) : '0;
logic [15:0] relu_121;
assign relu_121[15:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[29:15]}} :'d6) : '0;
logic [15:0] relu_122;
assign relu_122[15:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[29:15]}} :'d6) : '0;
logic [15:0] relu_123;
assign relu_123[15:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[29:15]}} :'d6) : '0;
logic [15:0] relu_124;
assign relu_124[15:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[29:15]}} :'d6) : '0;
logic [15:0] relu_125;
assign relu_125[15:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[29:15]}} :'d6) : '0;
logic [15:0] relu_126;
assign relu_126[15:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[29:15]}} :'d6) : '0;
logic [15:0] relu_127;
assign relu_127[15:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[29:15]}} :'d6) : '0;

assign output_act = {
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
