module conv2 (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [2400-1:0] input_act,
    output logic [256-1:0] output_act,
    output logic ready
);

logic [2400-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [399:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[399:0];
logic [399:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[799:400];
logic [399:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[1199:800];
logic [399:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[1599:1200];
logic [399:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[1999:1600];
logic [399:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[2399:2000];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	-2'sd 1 * $signed(input_fmap_0[31:16]) +
	-2'sd 1 * $signed(input_fmap_0[47:32]) +
	-2'sd 1 * $signed(input_fmap_0[63:48]) +
	-2'sd 1 * $signed(input_fmap_0[79:64]) +
	-3'sd 3 * $signed(input_fmap_0[95:80]) +
	-2'sd 1 * $signed(input_fmap_0[111:96]) +
	 4'sd 4 * $signed(input_fmap_0[127:112]) +
	 4'sd 5 * $signed(input_fmap_0[143:128]) +
	 3'sd 3 * $signed(input_fmap_0[159:144]) +
	-4'sd 4 * $signed(input_fmap_0[175:160]) +
	 2'sd 1 * $signed(input_fmap_0[191:176]) +
	 4'sd 6 * $signed(input_fmap_0[207:192]) +
	 4'sd 6 * $signed(input_fmap_0[223:208]) +
	 3'sd 3 * $signed(input_fmap_0[239:224]) +
	-3'sd 3 * $signed(input_fmap_0[255:240]) +
	-3'sd 2 * $signed(input_fmap_0[271:256]) +
	-3'sd 2 * $signed(input_fmap_0[287:272]) +
	-3'sd 2 * $signed(input_fmap_0[303:288]) +
	 2'sd 1 * $signed(input_fmap_0[319:304]) +
	-2'sd 1 * $signed(input_fmap_0[335:320]) +
	 2'sd 1 * $signed(input_fmap_0[351:336]) +
	 3'sd 2 * $signed(input_fmap_0[367:352]) +
	 3'sd 3 * $signed(input_fmap_0[383:368]) +
	 2'sd 1 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[47:32]) +
	-2'sd 1 * $signed(input_fmap_1[63:48]) +
	-2'sd 1 * $signed(input_fmap_1[79:64]) +
	 2'sd 1 * $signed(input_fmap_1[111:96]) +
	-2'sd 1 * $signed(input_fmap_1[159:144]) +
	 3'sd 2 * $signed(input_fmap_1[191:176]) +
	 2'sd 1 * $signed(input_fmap_1[207:192]) +
	-3'sd 2 * $signed(input_fmap_1[255:240]) +
	-2'sd 1 * $signed(input_fmap_1[271:256]) +
	-2'sd 1 * $signed(input_fmap_1[287:272]) +
	-3'sd 3 * $signed(input_fmap_1[335:320]) +
	-3'sd 2 * $signed(input_fmap_1[351:336]) +
	-3'sd 3 * $signed(input_fmap_1[367:352]) +
	-2'sd 1 * $signed(input_fmap_1[383:368]) +
	-2'sd 1 * $signed(input_fmap_2[15:0]) +
	-2'sd 1 * $signed(input_fmap_2[47:32]) +
	-2'sd 1 * $signed(input_fmap_2[63:48]) +
	 3'sd 2 * $signed(input_fmap_2[111:96]) +
	 2'sd 1 * $signed(input_fmap_2[127:112]) +
	 2'sd 1 * $signed(input_fmap_2[175:160]) +
	 3'sd 3 * $signed(input_fmap_2[191:176]) +
	 3'sd 2 * $signed(input_fmap_2[207:192]) +
	 3'sd 2 * $signed(input_fmap_2[223:208]) +
	 2'sd 1 * $signed(input_fmap_2[239:224]) +
	-3'sd 2 * $signed(input_fmap_2[255:240]) +
	-2'sd 1 * $signed(input_fmap_2[271:256]) +
	-2'sd 1 * $signed(input_fmap_2[287:272]) +
	-3'sd 2 * $signed(input_fmap_2[335:320]) +
	-3'sd 2 * $signed(input_fmap_2[351:336]) +
	-3'sd 3 * $signed(input_fmap_2[367:352]) +
	-2'sd 1 * $signed(input_fmap_2[383:368]) +
	-2'sd 1 * $signed(input_fmap_3[15:0]) +
	-2'sd 1 * $signed(input_fmap_3[47:32]) +
	-2'sd 1 * $signed(input_fmap_3[63:48]) +
	-2'sd 1 * $signed(input_fmap_3[79:64]) +
	 2'sd 1 * $signed(input_fmap_3[111:96]) +
	 2'sd 1 * $signed(input_fmap_3[127:112]) +
	 2'sd 1 * $signed(input_fmap_3[175:160]) +
	 3'sd 2 * $signed(input_fmap_3[191:176]) +
	 3'sd 2 * $signed(input_fmap_3[207:192]) +
	 2'sd 1 * $signed(input_fmap_3[223:208]) +
	 2'sd 1 * $signed(input_fmap_3[239:224]) +
	-3'sd 2 * $signed(input_fmap_3[255:240]) +
	-2'sd 1 * $signed(input_fmap_3[271:256]) +
	-2'sd 1 * $signed(input_fmap_3[287:272]) +
	-3'sd 2 * $signed(input_fmap_3[335:320]) +
	-3'sd 2 * $signed(input_fmap_3[351:336]) +
	-3'sd 3 * $signed(input_fmap_3[367:352]) +
	-3'sd 2 * $signed(input_fmap_3[383:368]) +
	-2'sd 1 * $signed(input_fmap_4[15:0]) +
	-3'sd 2 * $signed(input_fmap_4[31:16]) +
	-3'sd 2 * $signed(input_fmap_4[47:32]) +
	-2'sd 1 * $signed(input_fmap_4[63:48]) +
	-2'sd 1 * $signed(input_fmap_4[95:80]) +
	 3'sd 2 * $signed(input_fmap_4[111:96]) +
	 2'sd 1 * $signed(input_fmap_4[127:112]) +
	 2'sd 1 * $signed(input_fmap_4[159:144]) +
	 2'sd 1 * $signed(input_fmap_4[175:160]) +
	 4'sd 4 * $signed(input_fmap_4[191:176]) +
	 3'sd 3 * $signed(input_fmap_4[207:192]) +
	 3'sd 2 * $signed(input_fmap_4[223:208]) +
	 2'sd 1 * $signed(input_fmap_4[239:224]) +
	-2'sd 1 * $signed(input_fmap_4[255:240]) +
	 2'sd 1 * $signed(input_fmap_4[287:272]) +
	 3'sd 2 * $signed(input_fmap_4[303:288]) +
	 2'sd 1 * $signed(input_fmap_4[319:304]) +
	-2'sd 1 * $signed(input_fmap_4[335:320]) +
	-3'sd 2 * $signed(input_fmap_4[351:336]) +
	-3'sd 3 * $signed(input_fmap_4[367:352]) +
	-2'sd 1 * $signed(input_fmap_4[383:368]) +
	-2'sd 1 * $signed(input_fmap_5[15:0]) +
	-2'sd 1 * $signed(input_fmap_5[31:16]) +
	-3'sd 2 * $signed(input_fmap_5[47:32]) +
	-2'sd 1 * $signed(input_fmap_5[63:48]) +
	 2'sd 1 * $signed(input_fmap_5[111:96]) +
	 2'sd 1 * $signed(input_fmap_5[175:160]) +
	 4'sd 4 * $signed(input_fmap_5[191:176]) +
	 3'sd 2 * $signed(input_fmap_5[207:192]) +
	 3'sd 2 * $signed(input_fmap_5[223:208]) +
	 2'sd 1 * $signed(input_fmap_5[239:224]) +
	-2'sd 1 * $signed(input_fmap_5[255:240]) +
	 2'sd 1 * $signed(input_fmap_5[303:288]) +
	 2'sd 1 * $signed(input_fmap_5[319:304]) +
	-3'sd 2 * $signed(input_fmap_5[335:320]) +
	-3'sd 2 * $signed(input_fmap_5[351:336]) +
	-3'sd 3 * $signed(input_fmap_5[367:352]) +
	-2'sd 1 * $signed(input_fmap_5[383:368]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	 3'sd 2 * $signed(input_fmap_0[15:0]) +
	 4'sd 4 * $signed(input_fmap_0[31:16]) +
	 4'sd 4 * $signed(input_fmap_0[47:32]) +
	 3'sd 3 * $signed(input_fmap_0[63:48]) +
	 3'sd 2 * $signed(input_fmap_0[79:64]) +
	 3'sd 2 * $signed(input_fmap_0[95:80]) +
	 4'sd 4 * $signed(input_fmap_0[111:96]) +
	 3'sd 3 * $signed(input_fmap_0[127:112]) +
	-3'sd 2 * $signed(input_fmap_0[175:160]) +
	-3'sd 3 * $signed(input_fmap_0[191:176]) +
	-4'sd 6 * $signed(input_fmap_0[207:192]) +
	-4'sd 5 * $signed(input_fmap_0[223:208]) +
	-2'sd 1 * $signed(input_fmap_0[239:224]) +
	 2'sd 1 * $signed(input_fmap_0[255:240]) +
	 2'sd 1 * $signed(input_fmap_0[271:256]) +
	-3'sd 3 * $signed(input_fmap_0[287:272]) +
	-3'sd 3 * $signed(input_fmap_0[303:288]) +
	-4'sd 4 * $signed(input_fmap_0[319:304]) +
	 4'sd 4 * $signed(input_fmap_0[335:320]) +
	 4'sd 4 * $signed(input_fmap_0[351:336]) +
	 3'sd 2 * $signed(input_fmap_0[367:352]) +
	 3'sd 2 * $signed(input_fmap_0[383:368]) +
	 3'sd 3 * $signed(input_fmap_0[399:384]) +
	 2'sd 1 * $signed(input_fmap_1[15:0]) +
	 2'sd 1 * $signed(input_fmap_1[31:16]) +
	 2'sd 1 * $signed(input_fmap_1[47:32]) +
	-2'sd 1 * $signed(input_fmap_1[63:48]) +
	-2'sd 1 * $signed(input_fmap_1[79:64]) +
	 2'sd 1 * $signed(input_fmap_1[95:80]) +
	 3'sd 2 * $signed(input_fmap_1[111:96]) +
	 3'sd 2 * $signed(input_fmap_1[127:112]) +
	 2'sd 1 * $signed(input_fmap_1[143:128]) +
	 2'sd 1 * $signed(input_fmap_1[159:144]) +
	-2'sd 1 * $signed(input_fmap_1[175:160]) +
	-2'sd 1 * $signed(input_fmap_1[207:192]) +
	 3'sd 2 * $signed(input_fmap_1[239:224]) +
	-3'sd 2 * $signed(input_fmap_1[255:240]) +
	-3'sd 3 * $signed(input_fmap_1[271:256]) +
	-3'sd 3 * $signed(input_fmap_1[287:272]) +
	-3'sd 2 * $signed(input_fmap_1[303:288]) +
	 2'sd 1 * $signed(input_fmap_1[335:320]) +
	-3'sd 2 * $signed(input_fmap_1[351:336]) +
	-3'sd 2 * $signed(input_fmap_1[367:352]) +
	-2'sd 1 * $signed(input_fmap_1[383:368]) +
	-3'sd 2 * $signed(input_fmap_1[399:384]) +
	 2'sd 1 * $signed(input_fmap_2[31:16]) +
	 2'sd 1 * $signed(input_fmap_2[47:32]) +
	-2'sd 1 * $signed(input_fmap_2[79:64]) +
	 2'sd 1 * $signed(input_fmap_2[95:80]) +
	 3'sd 2 * $signed(input_fmap_2[111:96]) +
	 3'sd 2 * $signed(input_fmap_2[127:112]) +
	 2'sd 1 * $signed(input_fmap_2[143:128]) +
	 3'sd 2 * $signed(input_fmap_2[159:144]) +
	-2'sd 1 * $signed(input_fmap_2[175:160]) +
	 3'sd 2 * $signed(input_fmap_2[239:224]) +
	-3'sd 2 * $signed(input_fmap_2[255:240]) +
	-3'sd 3 * $signed(input_fmap_2[271:256]) +
	-3'sd 3 * $signed(input_fmap_2[287:272]) +
	-3'sd 3 * $signed(input_fmap_2[303:288]) +
	-2'sd 1 * $signed(input_fmap_2[319:304]) +
	-2'sd 1 * $signed(input_fmap_2[351:336]) +
	-2'sd 1 * $signed(input_fmap_2[367:352]) +
	-2'sd 1 * $signed(input_fmap_2[383:368]) +
	-2'sd 1 * $signed(input_fmap_2[399:384]) +
	 2'sd 1 * $signed(input_fmap_3[31:16]) +
	-2'sd 1 * $signed(input_fmap_3[79:64]) +
	 2'sd 1 * $signed(input_fmap_3[95:80]) +
	 3'sd 2 * $signed(input_fmap_3[111:96]) +
	 3'sd 2 * $signed(input_fmap_3[127:112]) +
	 2'sd 1 * $signed(input_fmap_3[143:128]) +
	 3'sd 2 * $signed(input_fmap_3[159:144]) +
	-2'sd 1 * $signed(input_fmap_3[175:160]) +
	-2'sd 1 * $signed(input_fmap_3[207:192]) +
	 3'sd 2 * $signed(input_fmap_3[239:224]) +
	-3'sd 2 * $signed(input_fmap_3[255:240]) +
	-3'sd 3 * $signed(input_fmap_3[271:256]) +
	-3'sd 3 * $signed(input_fmap_3[287:272]) +
	-3'sd 3 * $signed(input_fmap_3[303:288]) +
	-2'sd 1 * $signed(input_fmap_3[319:304]) +
	-2'sd 1 * $signed(input_fmap_3[351:336]) +
	-3'sd 2 * $signed(input_fmap_3[367:352]) +
	-2'sd 1 * $signed(input_fmap_3[383:368]) +
	-2'sd 1 * $signed(input_fmap_3[399:384]) +
	 2'sd 1 * $signed(input_fmap_4[31:16]) +
	-2'sd 1 * $signed(input_fmap_4[79:64]) +
	 3'sd 2 * $signed(input_fmap_4[95:80]) +
	 3'sd 3 * $signed(input_fmap_4[111:96]) +
	 3'sd 2 * $signed(input_fmap_4[127:112]) +
	 3'sd 2 * $signed(input_fmap_4[143:128]) +
	 3'sd 2 * $signed(input_fmap_4[159:144]) +
	 2'sd 1 * $signed(input_fmap_4[191:176]) +
	 2'sd 1 * $signed(input_fmap_4[207:192]) +
	 2'sd 1 * $signed(input_fmap_4[223:208]) +
	 4'sd 4 * $signed(input_fmap_4[239:224]) +
	-3'sd 3 * $signed(input_fmap_4[255:240]) +
	-4'sd 4 * $signed(input_fmap_4[271:256]) +
	-3'sd 3 * $signed(input_fmap_4[287:272]) +
	-3'sd 2 * $signed(input_fmap_4[303:288]) +
	-2'sd 1 * $signed(input_fmap_4[335:320]) +
	-2'sd 1 * $signed(input_fmap_4[351:336]) +
	-3'sd 2 * $signed(input_fmap_4[367:352]) +
	-2'sd 1 * $signed(input_fmap_4[383:368]) +
	-3'sd 3 * $signed(input_fmap_4[399:384]) +
	 2'sd 1 * $signed(input_fmap_5[31:16]) +
	-2'sd 1 * $signed(input_fmap_5[79:64]) +
	 3'sd 2 * $signed(input_fmap_5[95:80]) +
	 3'sd 2 * $signed(input_fmap_5[111:96]) +
	 3'sd 2 * $signed(input_fmap_5[127:112]) +
	 3'sd 2 * $signed(input_fmap_5[143:128]) +
	 3'sd 2 * $signed(input_fmap_5[159:144]) +
	-2'sd 1 * $signed(input_fmap_5[175:160]) +
	 2'sd 1 * $signed(input_fmap_5[223:208]) +
	 3'sd 3 * $signed(input_fmap_5[239:224]) +
	-3'sd 2 * $signed(input_fmap_5[255:240]) +
	-4'sd 4 * $signed(input_fmap_5[271:256]) +
	-3'sd 3 * $signed(input_fmap_5[287:272]) +
	-3'sd 2 * $signed(input_fmap_5[303:288]) +
	-2'sd 1 * $signed(input_fmap_5[319:304]) +
	-2'sd 1 * $signed(input_fmap_5[351:336]) +
	-3'sd 2 * $signed(input_fmap_5[367:352]) +
	-2'sd 1 * $signed(input_fmap_5[383:368]) +
	-3'sd 2 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	-3'sd 2 * $signed(input_fmap_0[15:0]) +
	-3'sd 2 * $signed(input_fmap_0[31:16]) +
	-4'sd 5 * $signed(input_fmap_0[47:32]) +
	-3'sd 3 * $signed(input_fmap_0[63:48]) +
	 3'sd 3 * $signed(input_fmap_0[79:64]) +
	-3'sd 2 * $signed(input_fmap_0[95:80]) +
	-4'sd 5 * $signed(input_fmap_0[111:96]) +
	-4'sd 5 * $signed(input_fmap_0[127:112]) +
	-2'sd 1 * $signed(input_fmap_0[143:128]) +
	 2'sd 1 * $signed(input_fmap_0[159:144]) +
	-4'sd 5 * $signed(input_fmap_0[175:160]) +
	-4'sd 5 * $signed(input_fmap_0[191:176]) +
	-2'sd 1 * $signed(input_fmap_0[207:192]) +
	-3'sd 2 * $signed(input_fmap_0[223:208]) +
	-4'sd 4 * $signed(input_fmap_0[239:224]) +
	-4'sd 5 * $signed(input_fmap_0[255:240]) +
	-3'sd 2 * $signed(input_fmap_0[271:256]) +
	 3'sd 2 * $signed(input_fmap_0[287:272]) +
	 3'sd 2 * $signed(input_fmap_0[303:288]) +
	 2'sd 1 * $signed(input_fmap_0[319:304]) +
	-2'sd 1 * $signed(input_fmap_0[335:320]) +
	 3'sd 2 * $signed(input_fmap_0[351:336]) +
	 3'sd 2 * $signed(input_fmap_0[367:352]) +
	 3'sd 2 * $signed(input_fmap_0[383:368]) +
	 3'sd 3 * $signed(input_fmap_0[399:384]) +
	 3'sd 2 * $signed(input_fmap_1[15:0]) +
	 3'sd 2 * $signed(input_fmap_1[31:16]) +
	-2'sd 1 * $signed(input_fmap_1[47:32]) +
	-3'sd 2 * $signed(input_fmap_1[63:48]) +
	-2'sd 1 * $signed(input_fmap_1[79:64]) +
	 4'sd 4 * $signed(input_fmap_1[95:80]) +
	 2'sd 1 * $signed(input_fmap_1[111:96]) +
	-3'sd 3 * $signed(input_fmap_1[127:112]) +
	-3'sd 2 * $signed(input_fmap_1[143:128]) +
	 4'sd 4 * $signed(input_fmap_1[175:160]) +
	 2'sd 1 * $signed(input_fmap_1[191:176]) +
	-3'sd 3 * $signed(input_fmap_1[207:192]) +
	-2'sd 1 * $signed(input_fmap_1[223:208]) +
	-3'sd 2 * $signed(input_fmap_1[239:224]) +
	 3'sd 2 * $signed(input_fmap_1[255:240]) +
	 2'sd 1 * $signed(input_fmap_1[271:256]) +
	-2'sd 1 * $signed(input_fmap_1[287:272]) +
	 3'sd 2 * $signed(input_fmap_1[335:320]) +
	 2'sd 1 * $signed(input_fmap_1[351:336]) +
	 2'sd 1 * $signed(input_fmap_1[367:352]) +
	 3'sd 2 * $signed(input_fmap_1[383:368]) +
	 2'sd 1 * $signed(input_fmap_1[399:384]) +
	 3'sd 2 * $signed(input_fmap_2[31:16]) +
	-2'sd 1 * $signed(input_fmap_2[63:48]) +
	-2'sd 1 * $signed(input_fmap_2[79:64]) +
	 2'sd 1 * $signed(input_fmap_2[95:80]) +
	 2'sd 1 * $signed(input_fmap_2[111:96]) +
	-3'sd 2 * $signed(input_fmap_2[127:112]) +
	-3'sd 2 * $signed(input_fmap_2[143:128]) +
	 3'sd 2 * $signed(input_fmap_2[175:160]) +
	 2'sd 1 * $signed(input_fmap_2[191:176]) +
	-3'sd 2 * $signed(input_fmap_2[207:192]) +
	-3'sd 3 * $signed(input_fmap_2[223:208]) +
	-3'sd 2 * $signed(input_fmap_2[239:224]) +
	 3'sd 2 * $signed(input_fmap_2[255:240]) +
	 2'sd 1 * $signed(input_fmap_2[271:256]) +
	 2'sd 1 * $signed(input_fmap_2[335:320]) +
	 2'sd 1 * $signed(input_fmap_2[351:336]) +
	 2'sd 1 * $signed(input_fmap_2[367:352]) +
	 3'sd 2 * $signed(input_fmap_2[383:368]) +
	 3'sd 2 * $signed(input_fmap_2[399:384]) +
	 3'sd 2 * $signed(input_fmap_3[31:16]) +
	-2'sd 1 * $signed(input_fmap_3[63:48]) +
	-2'sd 1 * $signed(input_fmap_3[79:64]) +
	 3'sd 2 * $signed(input_fmap_3[95:80]) +
	 3'sd 2 * $signed(input_fmap_3[111:96]) +
	-3'sd 2 * $signed(input_fmap_3[127:112]) +
	-3'sd 3 * $signed(input_fmap_3[143:128]) +
	 3'sd 3 * $signed(input_fmap_3[175:160]) +
	 2'sd 1 * $signed(input_fmap_3[191:176]) +
	-3'sd 2 * $signed(input_fmap_3[207:192]) +
	-3'sd 2 * $signed(input_fmap_3[223:208]) +
	-3'sd 2 * $signed(input_fmap_3[239:224]) +
	 3'sd 2 * $signed(input_fmap_3[255:240]) +
	 2'sd 1 * $signed(input_fmap_3[271:256]) +
	 3'sd 2 * $signed(input_fmap_3[335:320]) +
	 3'sd 2 * $signed(input_fmap_3[351:336]) +
	 2'sd 1 * $signed(input_fmap_3[367:352]) +
	 3'sd 2 * $signed(input_fmap_3[383:368]) +
	 2'sd 1 * $signed(input_fmap_3[399:384]) +
	-2'sd 1 * $signed(input_fmap_4[63:48]) +
	-2'sd 1 * $signed(input_fmap_4[79:64]) +
	-2'sd 1 * $signed(input_fmap_4[127:112]) +
	-3'sd 2 * $signed(input_fmap_4[143:128]) +
	 2'sd 1 * $signed(input_fmap_4[191:176]) +
	-3'sd 2 * $signed(input_fmap_4[207:192]) +
	-3'sd 3 * $signed(input_fmap_4[223:208]) +
	-3'sd 3 * $signed(input_fmap_4[239:224]) +
	 2'sd 1 * $signed(input_fmap_4[255:240]) +
	 2'sd 1 * $signed(input_fmap_4[271:256]) +
	-2'sd 1 * $signed(input_fmap_4[287:272]) +
	-2'sd 1 * $signed(input_fmap_4[303:288]) +
	-2'sd 1 * $signed(input_fmap_4[319:304]) +
	 2'sd 1 * $signed(input_fmap_4[335:320]) +
	 2'sd 1 * $signed(input_fmap_4[351:336]) +
	 2'sd 1 * $signed(input_fmap_4[367:352]) +
	 3'sd 2 * $signed(input_fmap_4[383:368]) +
	 3'sd 2 * $signed(input_fmap_4[399:384]) +
	 2'sd 1 * $signed(input_fmap_5[31:16]) +
	-2'sd 1 * $signed(input_fmap_5[63:48]) +
	-2'sd 1 * $signed(input_fmap_5[79:64]) +
	 2'sd 1 * $signed(input_fmap_5[95:80]) +
	 2'sd 1 * $signed(input_fmap_5[111:96]) +
	-3'sd 2 * $signed(input_fmap_5[127:112]) +
	-3'sd 2 * $signed(input_fmap_5[143:128]) +
	 3'sd 2 * $signed(input_fmap_5[175:160]) +
	 2'sd 1 * $signed(input_fmap_5[191:176]) +
	-3'sd 2 * $signed(input_fmap_5[207:192]) +
	-3'sd 3 * $signed(input_fmap_5[223:208]) +
	-3'sd 2 * $signed(input_fmap_5[239:224]) +
	 3'sd 2 * $signed(input_fmap_5[255:240]) +
	 2'sd 1 * $signed(input_fmap_5[271:256]) +
	-2'sd 1 * $signed(input_fmap_5[287:272]) +
	-2'sd 1 * $signed(input_fmap_5[303:288]) +
	 2'sd 1 * $signed(input_fmap_5[335:320]) +
	 2'sd 1 * $signed(input_fmap_5[351:336]) +
	 2'sd 1 * $signed(input_fmap_5[367:352]) +
	 3'sd 2 * $signed(input_fmap_5[383:368]) +
	 3'sd 2 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	-2'sd 1 * $signed(input_fmap_0[47:32]) +
	 3'sd 2 * $signed(input_fmap_0[95:80]) +
	 3'sd 3 * $signed(input_fmap_0[207:192]) +
	 4'sd 6 * $signed(input_fmap_0[223:208]) +
	 4'sd 6 * $signed(input_fmap_0[239:224]) +
	-4'sd 6 * $signed(input_fmap_0[255:240]) +
	-5'sd 8 * $signed(input_fmap_0[271:256]) +
	-4'sd 6 * $signed(input_fmap_0[287:272]) +
	-3'sd 2 * $signed(input_fmap_0[303:288]) +
	 2'sd 1 * $signed(input_fmap_0[319:304]) +
	-2'sd 1 * $signed(input_fmap_0[335:320]) +
	 2'sd 1 * $signed(input_fmap_0[367:352]) +
	 2'sd 1 * $signed(input_fmap_0[383:368]) +
	-3'sd 2 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[79:64]) +
	 2'sd 1 * $signed(input_fmap_1[95:80]) +
	-2'sd 1 * $signed(input_fmap_1[111:96]) +
	-2'sd 1 * $signed(input_fmap_1[143:128]) +
	-3'sd 2 * $signed(input_fmap_1[159:144]) +
	 2'sd 1 * $signed(input_fmap_1[191:176]) +
	 3'sd 2 * $signed(input_fmap_1[207:192]) +
	 2'sd 1 * $signed(input_fmap_1[223:208]) +
	 2'sd 1 * $signed(input_fmap_1[239:224]) +
	-3'sd 3 * $signed(input_fmap_1[255:240]) +
	-3'sd 2 * $signed(input_fmap_1[271:256]) +
	 2'sd 1 * $signed(input_fmap_1[319:304]) +
	-4'sd 5 * $signed(input_fmap_1[335:320]) +
	-3'sd 3 * $signed(input_fmap_1[351:336]) +
	-3'sd 2 * $signed(input_fmap_1[367:352]) +
	-3'sd 2 * $signed(input_fmap_1[383:368]) +
	-3'sd 2 * $signed(input_fmap_1[399:384]) +
	-2'sd 1 * $signed(input_fmap_2[15:0]) +
	-2'sd 1 * $signed(input_fmap_2[31:16]) +
	-2'sd 1 * $signed(input_fmap_2[47:32]) +
	 2'sd 1 * $signed(input_fmap_2[95:80]) +
	-2'sd 1 * $signed(input_fmap_2[143:128]) +
	-2'sd 1 * $signed(input_fmap_2[159:144]) +
	 2'sd 1 * $signed(input_fmap_2[175:160]) +
	 3'sd 2 * $signed(input_fmap_2[191:176]) +
	 3'sd 3 * $signed(input_fmap_2[207:192]) +
	 3'sd 3 * $signed(input_fmap_2[223:208]) +
	 2'sd 1 * $signed(input_fmap_2[239:224]) +
	-3'sd 3 * $signed(input_fmap_2[255:240]) +
	-3'sd 3 * $signed(input_fmap_2[271:256]) +
	 3'sd 2 * $signed(input_fmap_2[303:288]) +
	 3'sd 2 * $signed(input_fmap_2[319:304]) +
	-4'sd 4 * $signed(input_fmap_2[335:320]) +
	-4'sd 4 * $signed(input_fmap_2[351:336]) +
	-3'sd 3 * $signed(input_fmap_2[367:352]) +
	-3'sd 3 * $signed(input_fmap_2[383:368]) +
	-3'sd 2 * $signed(input_fmap_2[399:384]) +
	-2'sd 1 * $signed(input_fmap_3[15:0]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	-2'sd 1 * $signed(input_fmap_3[47:32]) +
	-2'sd 1 * $signed(input_fmap_3[79:64]) +
	 2'sd 1 * $signed(input_fmap_3[95:80]) +
	-2'sd 1 * $signed(input_fmap_3[143:128]) +
	-3'sd 2 * $signed(input_fmap_3[159:144]) +
	 2'sd 1 * $signed(input_fmap_3[175:160]) +
	 3'sd 2 * $signed(input_fmap_3[191:176]) +
	 3'sd 2 * $signed(input_fmap_3[207:192]) +
	 3'sd 2 * $signed(input_fmap_3[223:208]) +
	 2'sd 1 * $signed(input_fmap_3[239:224]) +
	-3'sd 3 * $signed(input_fmap_3[255:240]) +
	-3'sd 3 * $signed(input_fmap_3[271:256]) +
	 2'sd 1 * $signed(input_fmap_3[303:288]) +
	 2'sd 1 * $signed(input_fmap_3[319:304]) +
	-4'sd 4 * $signed(input_fmap_3[335:320]) +
	-4'sd 4 * $signed(input_fmap_3[351:336]) +
	-3'sd 3 * $signed(input_fmap_3[367:352]) +
	-3'sd 3 * $signed(input_fmap_3[383:368]) +
	-3'sd 2 * $signed(input_fmap_3[399:384]) +
	-2'sd 1 * $signed(input_fmap_4[15:0]) +
	-3'sd 2 * $signed(input_fmap_4[31:16]) +
	-2'sd 1 * $signed(input_fmap_4[47:32]) +
	-2'sd 1 * $signed(input_fmap_4[127:112]) +
	-2'sd 1 * $signed(input_fmap_4[143:128]) +
	 3'sd 2 * $signed(input_fmap_4[175:160]) +
	 4'sd 4 * $signed(input_fmap_4[191:176]) +
	 4'sd 4 * $signed(input_fmap_4[207:192]) +
	 3'sd 2 * $signed(input_fmap_4[223:208]) +
	 2'sd 1 * $signed(input_fmap_4[239:224]) +
	-3'sd 2 * $signed(input_fmap_4[255:240]) +
	-2'sd 1 * $signed(input_fmap_4[271:256]) +
	 3'sd 2 * $signed(input_fmap_4[287:272]) +
	 3'sd 3 * $signed(input_fmap_4[303:288]) +
	 3'sd 2 * $signed(input_fmap_4[319:304]) +
	-4'sd 4 * $signed(input_fmap_4[335:320]) +
	-4'sd 4 * $signed(input_fmap_4[351:336]) +
	-4'sd 4 * $signed(input_fmap_4[367:352]) +
	-3'sd 2 * $signed(input_fmap_4[383:368]) +
	-2'sd 1 * $signed(input_fmap_4[399:384]) +
	-2'sd 1 * $signed(input_fmap_5[15:0]) +
	-2'sd 1 * $signed(input_fmap_5[31:16]) +
	-2'sd 1 * $signed(input_fmap_5[47:32]) +
	 2'sd 1 * $signed(input_fmap_5[95:80]) +
	-2'sd 1 * $signed(input_fmap_5[127:112]) +
	-2'sd 1 * $signed(input_fmap_5[143:128]) +
	-2'sd 1 * $signed(input_fmap_5[159:144]) +
	 3'sd 2 * $signed(input_fmap_5[175:160]) +
	 3'sd 3 * $signed(input_fmap_5[191:176]) +
	 3'sd 3 * $signed(input_fmap_5[207:192]) +
	 3'sd 2 * $signed(input_fmap_5[223:208]) +
	 2'sd 1 * $signed(input_fmap_5[239:224]) +
	-3'sd 2 * $signed(input_fmap_5[255:240]) +
	-2'sd 1 * $signed(input_fmap_5[271:256]) +
	 2'sd 1 * $signed(input_fmap_5[287:272]) +
	 3'sd 2 * $signed(input_fmap_5[303:288]) +
	 3'sd 2 * $signed(input_fmap_5[319:304]) +
	-4'sd 4 * $signed(input_fmap_5[335:320]) +
	-4'sd 4 * $signed(input_fmap_5[351:336]) +
	-3'sd 3 * $signed(input_fmap_5[367:352]) +
	-3'sd 2 * $signed(input_fmap_5[383:368]) +
	-2'sd 1 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 32'sd 0;

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	-4'sd 4 * $signed(input_fmap_0[31:16]) +
	-4'sd 7 * $signed(input_fmap_0[47:32]) +
	-4'sd 6 * $signed(input_fmap_0[63:48]) +
	 3'sd 2 * $signed(input_fmap_0[79:64]) +
	 4'sd 4 * $signed(input_fmap_0[95:80]) +
	 3'sd 2 * $signed(input_fmap_0[111:96]) +
	-3'sd 3 * $signed(input_fmap_0[127:112]) +
	-4'sd 6 * $signed(input_fmap_0[143:128]) +
	-5'sd 9 * $signed(input_fmap_0[159:144]) +
	 3'sd 3 * $signed(input_fmap_0[175:160]) +
	 4'sd 4 * $signed(input_fmap_0[191:176]) +
	 4'sd 4 * $signed(input_fmap_0[207:192]) +
	 4'sd 4 * $signed(input_fmap_0[223:208]) +
	 3'sd 3 * $signed(input_fmap_0[239:224]) +
	 4'sd 4 * $signed(input_fmap_0[303:288]) +
	 4'sd 5 * $signed(input_fmap_0[319:304]) +
	-2'sd 1 * $signed(input_fmap_0[335:320]) +
	-4'sd 4 * $signed(input_fmap_0[351:336]) +
	-4'sd 4 * $signed(input_fmap_0[367:352]) +
	-3'sd 2 * $signed(input_fmap_0[383:368]) +
	-2'sd 1 * $signed(input_fmap_0[399:384]) +
	-3'sd 3 * $signed(input_fmap_1[15:0]) +
	-3'sd 2 * $signed(input_fmap_1[31:16]) +
	-3'sd 3 * $signed(input_fmap_1[47:32]) +
	-2'sd 1 * $signed(input_fmap_1[63:48]) +
	 4'sd 4 * $signed(input_fmap_1[79:64]) +
	-2'sd 1 * $signed(input_fmap_1[95:80]) +
	-3'sd 3 * $signed(input_fmap_1[111:96]) +
	-4'sd 4 * $signed(input_fmap_1[127:112]) +
	-4'sd 4 * $signed(input_fmap_1[143:128]) +
	 2'sd 1 * $signed(input_fmap_1[175:160]) +
	-2'sd 1 * $signed(input_fmap_1[191:176]) +
	-3'sd 2 * $signed(input_fmap_1[223:208]) +
	-3'sd 2 * $signed(input_fmap_1[239:224]) +
	 2'sd 1 * $signed(input_fmap_1[255:240]) +
	 2'sd 1 * $signed(input_fmap_1[271:256]) +
	 2'sd 1 * $signed(input_fmap_1[287:272]) +
	 2'sd 1 * $signed(input_fmap_1[351:336]) +
	 2'sd 1 * $signed(input_fmap_1[367:352]) +
	 2'sd 1 * $signed(input_fmap_1[383:368]) +
	-3'sd 3 * $signed(input_fmap_2[15:0]) +
	-3'sd 3 * $signed(input_fmap_2[31:16]) +
	-3'sd 3 * $signed(input_fmap_2[47:32]) +
	-2'sd 1 * $signed(input_fmap_2[63:48]) +
	 3'sd 3 * $signed(input_fmap_2[79:64]) +
	-2'sd 1 * $signed(input_fmap_2[111:96]) +
	-3'sd 3 * $signed(input_fmap_2[127:112]) +
	-4'sd 6 * $signed(input_fmap_2[143:128]) +
	-3'sd 3 * $signed(input_fmap_2[159:144]) +
	 3'sd 2 * $signed(input_fmap_2[175:160]) +
	 2'sd 1 * $signed(input_fmap_2[191:176]) +
	 2'sd 1 * $signed(input_fmap_2[207:192]) +
	-2'sd 1 * $signed(input_fmap_2[239:224]) +
	 2'sd 1 * $signed(input_fmap_2[255:240]) +
	 2'sd 1 * $signed(input_fmap_2[271:256]) +
	 3'sd 2 * $signed(input_fmap_2[287:272]) +
	 3'sd 2 * $signed(input_fmap_2[303:288]) +
	 3'sd 2 * $signed(input_fmap_2[319:304]) +
	-2'sd 1 * $signed(input_fmap_2[335:320]) +
	 2'sd 1 * $signed(input_fmap_2[367:352]) +
	 2'sd 1 * $signed(input_fmap_2[399:384]) +
	-3'sd 3 * $signed(input_fmap_3[15:0]) +
	-3'sd 3 * $signed(input_fmap_3[31:16]) +
	-3'sd 3 * $signed(input_fmap_3[47:32]) +
	-3'sd 2 * $signed(input_fmap_3[63:48]) +
	 3'sd 3 * $signed(input_fmap_3[79:64]) +
	-3'sd 2 * $signed(input_fmap_3[111:96]) +
	-3'sd 3 * $signed(input_fmap_3[127:112]) +
	-4'sd 6 * $signed(input_fmap_3[143:128]) +
	-3'sd 2 * $signed(input_fmap_3[159:144]) +
	 2'sd 1 * $signed(input_fmap_3[175:160]) +
	 2'sd 1 * $signed(input_fmap_3[191:176]) +
	-2'sd 1 * $signed(input_fmap_3[223:208]) +
	-3'sd 2 * $signed(input_fmap_3[239:224]) +
	 2'sd 1 * $signed(input_fmap_3[255:240]) +
	 2'sd 1 * $signed(input_fmap_3[271:256]) +
	 3'sd 2 * $signed(input_fmap_3[287:272]) +
	 2'sd 1 * $signed(input_fmap_3[303:288]) +
	 2'sd 1 * $signed(input_fmap_3[319:304]) +
	-2'sd 1 * $signed(input_fmap_3[335:320]) +
	 2'sd 1 * $signed(input_fmap_3[367:352]) +
	 2'sd 1 * $signed(input_fmap_3[399:384]) +
	-3'sd 3 * $signed(input_fmap_4[15:0]) +
	-3'sd 3 * $signed(input_fmap_4[31:16]) +
	-3'sd 2 * $signed(input_fmap_4[47:32]) +
	 3'sd 3 * $signed(input_fmap_4[79:64]) +
	-3'sd 2 * $signed(input_fmap_4[111:96]) +
	-4'sd 4 * $signed(input_fmap_4[127:112]) +
	-4'sd 6 * $signed(input_fmap_4[143:128]) +
	-2'sd 1 * $signed(input_fmap_4[159:144]) +
	 3'sd 3 * $signed(input_fmap_4[175:160]) +
	 3'sd 2 * $signed(input_fmap_4[191:176]) +
	 2'sd 1 * $signed(input_fmap_4[207:192]) +
	-3'sd 2 * $signed(input_fmap_4[223:208]) +
	-3'sd 3 * $signed(input_fmap_4[239:224]) +
	 2'sd 1 * $signed(input_fmap_4[255:240]) +
	 3'sd 3 * $signed(input_fmap_4[271:256]) +
	 3'sd 3 * $signed(input_fmap_4[287:272]) +
	 3'sd 3 * $signed(input_fmap_4[303:288]) +
	 3'sd 2 * $signed(input_fmap_4[319:304]) +
	-2'sd 1 * $signed(input_fmap_4[335:320]) +
	 2'sd 1 * $signed(input_fmap_4[367:352]) +
	 3'sd 2 * $signed(input_fmap_4[383:368]) +
	 2'sd 1 * $signed(input_fmap_4[399:384]) +
	-3'sd 3 * $signed(input_fmap_5[15:0]) +
	-3'sd 3 * $signed(input_fmap_5[31:16]) +
	-3'sd 3 * $signed(input_fmap_5[47:32]) +
	-2'sd 1 * $signed(input_fmap_5[63:48]) +
	 3'sd 3 * $signed(input_fmap_5[79:64]) +
	-3'sd 2 * $signed(input_fmap_5[111:96]) +
	-4'sd 4 * $signed(input_fmap_5[127:112]) +
	-4'sd 6 * $signed(input_fmap_5[143:128]) +
	-3'sd 2 * $signed(input_fmap_5[159:144]) +
	 3'sd 2 * $signed(input_fmap_5[175:160]) +
	 2'sd 1 * $signed(input_fmap_5[191:176]) +
	 2'sd 1 * $signed(input_fmap_5[207:192]) +
	-2'sd 1 * $signed(input_fmap_5[223:208]) +
	-3'sd 2 * $signed(input_fmap_5[239:224]) +
	 2'sd 1 * $signed(input_fmap_5[255:240]) +
	 3'sd 2 * $signed(input_fmap_5[271:256]) +
	 3'sd 2 * $signed(input_fmap_5[287:272]) +
	 3'sd 2 * $signed(input_fmap_5[303:288]) +
	 3'sd 2 * $signed(input_fmap_5[319:304]) +
	 2'sd 1 * $signed(input_fmap_5[367:352]) +
	 2'sd 1 * $signed(input_fmap_5[383:368]) +
	 2'sd 1 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	 3'sd 3 * $signed(input_fmap_0[15:0]) +
	 2'sd 1 * $signed(input_fmap_0[31:16]) +
	-2'sd 1 * $signed(input_fmap_0[47:32]) +
	-4'sd 4 * $signed(input_fmap_0[63:48]) +
	-4'sd 4 * $signed(input_fmap_0[79:64]) +
	 3'sd 3 * $signed(input_fmap_0[95:80]) +
	 3'sd 3 * $signed(input_fmap_0[111:96]) +
	-3'sd 2 * $signed(input_fmap_0[127:112]) +
	-4'sd 5 * $signed(input_fmap_0[143:128]) +
	-3'sd 3 * $signed(input_fmap_0[159:144]) +
	 3'sd 3 * $signed(input_fmap_0[175:160]) +
	 2'sd 1 * $signed(input_fmap_0[191:176]) +
	-3'sd 3 * $signed(input_fmap_0[207:192]) +
	-4'sd 4 * $signed(input_fmap_0[223:208]) +
	 2'sd 1 * $signed(input_fmap_0[239:224]) +
	 4'sd 4 * $signed(input_fmap_0[255:240]) +
	-3'sd 2 * $signed(input_fmap_0[271:256]) +
	-4'sd 5 * $signed(input_fmap_0[287:272]) +
	-3'sd 3 * $signed(input_fmap_0[303:288]) +
	-2'sd 1 * $signed(input_fmap_0[319:304]) +
	-2'sd 1 * $signed(input_fmap_0[335:320]) +
	-4'sd 4 * $signed(input_fmap_0[351:336]) +
	-3'sd 3 * $signed(input_fmap_0[367:352]) +
	-3'sd 2 * $signed(input_fmap_0[383:368]) +
	-3'sd 2 * $signed(input_fmap_1[31:16]) +
	 3'sd 2 * $signed(input_fmap_1[63:48]) +
	 2'sd 1 * $signed(input_fmap_1[127:112]) +
	 3'sd 3 * $signed(input_fmap_1[143:128]) +
	-2'sd 1 * $signed(input_fmap_1[159:144]) +
	 3'sd 2 * $signed(input_fmap_1[175:160]) +
	 3'sd 2 * $signed(input_fmap_1[191:176]) +
	 2'sd 1 * $signed(input_fmap_1[207:192]) +
	 2'sd 1 * $signed(input_fmap_1[223:208]) +
	-2'sd 1 * $signed(input_fmap_1[239:224]) +
	 3'sd 2 * $signed(input_fmap_1[255:240]) +
	-2'sd 1 * $signed(input_fmap_1[319:304]) +
	 2'sd 1 * $signed(input_fmap_1[335:320]) +
	-2'sd 1 * $signed(input_fmap_1[351:336]) +
	-2'sd 1 * $signed(input_fmap_1[399:384]) +
	-2'sd 1 * $signed(input_fmap_2[31:16]) +
	-2'sd 1 * $signed(input_fmap_2[47:32]) +
	 2'sd 1 * $signed(input_fmap_2[63:48]) +
	 2'sd 1 * $signed(input_fmap_2[79:64]) +
	-2'sd 1 * $signed(input_fmap_2[127:112]) +
	 2'sd 1 * $signed(input_fmap_2[143:128]) +
	 2'sd 1 * $signed(input_fmap_2[159:144]) +
	 2'sd 1 * $signed(input_fmap_2[191:176]) +
	 3'sd 2 * $signed(input_fmap_2[223:208]) +
	-2'sd 1 * $signed(input_fmap_2[287:272]) +
	 2'sd 1 * $signed(input_fmap_2[303:288]) +
	 2'sd 1 * $signed(input_fmap_2[335:320]) +
	-2'sd 1 * $signed(input_fmap_2[367:352]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	-2'sd 1 * $signed(input_fmap_3[47:32]) +
	 2'sd 1 * $signed(input_fmap_3[63:48]) +
	 2'sd 1 * $signed(input_fmap_3[79:64]) +
	-2'sd 1 * $signed(input_fmap_3[95:80]) +
	-2'sd 1 * $signed(input_fmap_3[127:112]) +
	 3'sd 2 * $signed(input_fmap_3[143:128]) +
	 2'sd 1 * $signed(input_fmap_3[159:144]) +
	 2'sd 1 * $signed(input_fmap_3[191:176]) +
	 3'sd 2 * $signed(input_fmap_3[223:208]) +
	 2'sd 1 * $signed(input_fmap_3[255:240]) +
	 2'sd 1 * $signed(input_fmap_3[271:256]) +
	-2'sd 1 * $signed(input_fmap_3[287:272]) +
	 2'sd 1 * $signed(input_fmap_3[303:288]) +
	 2'sd 1 * $signed(input_fmap_3[335:320]) +
	-2'sd 1 * $signed(input_fmap_3[367:352]) +
	-2'sd 1 * $signed(input_fmap_3[399:384]) +
	 2'sd 1 * $signed(input_fmap_4[15:0]) +
	 2'sd 1 * $signed(input_fmap_4[47:32]) +
	-2'sd 1 * $signed(input_fmap_4[79:64]) +
	 2'sd 1 * $signed(input_fmap_4[95:80]) +
	-3'sd 2 * $signed(input_fmap_4[127:112]) +
	 2'sd 1 * $signed(input_fmap_4[191:176]) +
	-2'sd 1 * $signed(input_fmap_4[207:192]) +
	 2'sd 1 * $signed(input_fmap_4[223:208]) +
	 2'sd 1 * $signed(input_fmap_4[239:224]) +
	-2'sd 1 * $signed(input_fmap_4[287:272]) +
	 2'sd 1 * $signed(input_fmap_4[303:288]) +
	 2'sd 1 * $signed(input_fmap_4[319:304]) +
	-2'sd 1 * $signed(input_fmap_4[367:352]) +
	-2'sd 1 * $signed(input_fmap_4[399:384]) +
	 2'sd 1 * $signed(input_fmap_5[63:48]) +
	 2'sd 1 * $signed(input_fmap_5[143:128]) +
	 2'sd 1 * $signed(input_fmap_5[159:144]) +
	 2'sd 1 * $signed(input_fmap_5[175:160]) +
	 2'sd 1 * $signed(input_fmap_5[191:176]) +
	 2'sd 1 * $signed(input_fmap_5[223:208]) +
	 2'sd 1 * $signed(input_fmap_5[335:320]) +
	-2'sd 1 * $signed(input_fmap_5[367:352]) +
	-2'sd 1 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	-3'sd 2 * $signed(input_fmap_0[15:0]) +
	-2'sd 1 * $signed(input_fmap_0[31:16]) +
	-2'sd 1 * $signed(input_fmap_0[63:48]) +
	-2'sd 1 * $signed(input_fmap_0[79:64]) +
	 4'sd 4 * $signed(input_fmap_0[95:80]) +
	 4'sd 6 * $signed(input_fmap_0[111:96]) +
	 4'sd 7 * $signed(input_fmap_0[127:112]) +
	 4'sd 4 * $signed(input_fmap_0[143:128]) +
	 4'sd 4 * $signed(input_fmap_0[175:160]) +
	 4'sd 4 * $signed(input_fmap_0[191:176]) +
	 2'sd 1 * $signed(input_fmap_0[207:192]) +
	-3'sd 2 * $signed(input_fmap_0[223:208]) +
	-2'sd 1 * $signed(input_fmap_0[239:224]) +
	-3'sd 3 * $signed(input_fmap_0[255:240]) +
	-4'sd 4 * $signed(input_fmap_0[271:256]) +
	-3'sd 3 * $signed(input_fmap_0[287:272]) +
	-2'sd 1 * $signed(input_fmap_0[303:288]) +
	-2'sd 1 * $signed(input_fmap_0[319:304]) +
	 4'sd 5 * $signed(input_fmap_0[335:320]) +
	 4'sd 5 * $signed(input_fmap_0[351:336]) +
	 3'sd 3 * $signed(input_fmap_0[367:352]) +
	 2'sd 1 * $signed(input_fmap_0[383:368]) +
	-3'sd 2 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[31:16]) +
	-2'sd 1 * $signed(input_fmap_1[47:32]) +
	 2'sd 1 * $signed(input_fmap_1[79:64]) +
	 2'sd 1 * $signed(input_fmap_1[95:80]) +
	 2'sd 1 * $signed(input_fmap_1[111:96]) +
	 2'sd 1 * $signed(input_fmap_1[127:112]) +
	 2'sd 1 * $signed(input_fmap_1[159:144]) +
	 2'sd 1 * $signed(input_fmap_1[175:160]) +
	 2'sd 1 * $signed(input_fmap_1[191:176]) +
	 2'sd 1 * $signed(input_fmap_1[207:192]) +
	 2'sd 1 * $signed(input_fmap_1[239:224]) +
	-3'sd 2 * $signed(input_fmap_1[255:240]) +
	-3'sd 2 * $signed(input_fmap_1[271:256]) +
	-3'sd 2 * $signed(input_fmap_1[287:272]) +
	-3'sd 2 * $signed(input_fmap_1[303:288]) +
	 2'sd 1 * $signed(input_fmap_1[319:304]) +
	-3'sd 2 * $signed(input_fmap_1[335:320]) +
	-3'sd 3 * $signed(input_fmap_1[351:336]) +
	-2'sd 1 * $signed(input_fmap_1[367:352]) +
	-3'sd 2 * $signed(input_fmap_1[383:368]) +
	-2'sd 1 * $signed(input_fmap_1[399:384]) +
	-2'sd 1 * $signed(input_fmap_2[15:0]) +
	-2'sd 1 * $signed(input_fmap_2[47:32]) +
	-2'sd 1 * $signed(input_fmap_2[63:48]) +
	 2'sd 1 * $signed(input_fmap_2[95:80]) +
	 3'sd 2 * $signed(input_fmap_2[111:96]) +
	 3'sd 2 * $signed(input_fmap_2[127:112]) +
	 3'sd 2 * $signed(input_fmap_2[143:128]) +
	 2'sd 1 * $signed(input_fmap_2[159:144]) +
	 3'sd 2 * $signed(input_fmap_2[175:160]) +
	 3'sd 2 * $signed(input_fmap_2[191:176]) +
	 2'sd 1 * $signed(input_fmap_2[207:192]) +
	 2'sd 1 * $signed(input_fmap_2[223:208]) +
	 2'sd 1 * $signed(input_fmap_2[239:224]) +
	-3'sd 2 * $signed(input_fmap_2[255:240]) +
	-3'sd 2 * $signed(input_fmap_2[271:256]) +
	-3'sd 2 * $signed(input_fmap_2[287:272]) +
	-2'sd 1 * $signed(input_fmap_2[303:288]) +
	 2'sd 1 * $signed(input_fmap_2[319:304]) +
	-2'sd 1 * $signed(input_fmap_2[335:320]) +
	-3'sd 2 * $signed(input_fmap_2[351:336]) +
	-2'sd 1 * $signed(input_fmap_2[367:352]) +
	-2'sd 1 * $signed(input_fmap_2[383:368]) +
	-2'sd 1 * $signed(input_fmap_2[399:384]) +
	-2'sd 1 * $signed(input_fmap_3[15:0]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	-3'sd 2 * $signed(input_fmap_3[47:32]) +
	-2'sd 1 * $signed(input_fmap_3[63:48]) +
	 2'sd 1 * $signed(input_fmap_3[95:80]) +
	 2'sd 1 * $signed(input_fmap_3[111:96]) +
	 2'sd 1 * $signed(input_fmap_3[127:112]) +
	 2'sd 1 * $signed(input_fmap_3[143:128]) +
	 2'sd 1 * $signed(input_fmap_3[159:144]) +
	 2'sd 1 * $signed(input_fmap_3[175:160]) +
	 2'sd 1 * $signed(input_fmap_3[191:176]) +
	 2'sd 1 * $signed(input_fmap_3[207:192]) +
	 2'sd 1 * $signed(input_fmap_3[239:224]) +
	-3'sd 2 * $signed(input_fmap_3[255:240]) +
	-3'sd 2 * $signed(input_fmap_3[271:256]) +
	-3'sd 2 * $signed(input_fmap_3[287:272]) +
	-3'sd 2 * $signed(input_fmap_3[303:288]) +
	 2'sd 1 * $signed(input_fmap_3[319:304]) +
	-2'sd 1 * $signed(input_fmap_3[335:320]) +
	-3'sd 2 * $signed(input_fmap_3[351:336]) +
	-3'sd 2 * $signed(input_fmap_3[367:352]) +
	-2'sd 1 * $signed(input_fmap_3[383:368]) +
	-2'sd 1 * $signed(input_fmap_4[15:0]) +
	-2'sd 1 * $signed(input_fmap_4[31:16]) +
	-3'sd 2 * $signed(input_fmap_4[47:32]) +
	-3'sd 2 * $signed(input_fmap_4[63:48]) +
	-2'sd 1 * $signed(input_fmap_4[79:64]) +
	 2'sd 1 * $signed(input_fmap_4[111:96]) +
	 2'sd 1 * $signed(input_fmap_4[127:112]) +
	 2'sd 1 * $signed(input_fmap_4[143:128]) +
	 2'sd 1 * $signed(input_fmap_4[159:144]) +
	 3'sd 3 * $signed(input_fmap_4[175:160]) +
	 3'sd 3 * $signed(input_fmap_4[191:176]) +
	 3'sd 2 * $signed(input_fmap_4[207:192]) +
	 2'sd 1 * $signed(input_fmap_4[223:208]) +
	 3'sd 2 * $signed(input_fmap_4[239:224]) +
	-2'sd 1 * $signed(input_fmap_4[255:240]) +
	-2'sd 1 * $signed(input_fmap_4[271:256]) +
	-2'sd 1 * $signed(input_fmap_4[287:272]) +
	 2'sd 1 * $signed(input_fmap_4[319:304]) +
	-2'sd 1 * $signed(input_fmap_4[335:320]) +
	-3'sd 2 * $signed(input_fmap_4[351:336]) +
	-3'sd 2 * $signed(input_fmap_4[367:352]) +
	-3'sd 2 * $signed(input_fmap_4[383:368]) +
	-2'sd 1 * $signed(input_fmap_4[399:384]) +
	-2'sd 1 * $signed(input_fmap_5[15:0]) +
	-2'sd 1 * $signed(input_fmap_5[31:16]) +
	-3'sd 2 * $signed(input_fmap_5[47:32]) +
	-2'sd 1 * $signed(input_fmap_5[63:48]) +
	 2'sd 1 * $signed(input_fmap_5[111:96]) +
	 2'sd 1 * $signed(input_fmap_5[127:112]) +
	 2'sd 1 * $signed(input_fmap_5[143:128]) +
	 2'sd 1 * $signed(input_fmap_5[159:144]) +
	 3'sd 2 * $signed(input_fmap_5[175:160]) +
	 3'sd 2 * $signed(input_fmap_5[191:176]) +
	 2'sd 1 * $signed(input_fmap_5[207:192]) +
	 2'sd 1 * $signed(input_fmap_5[223:208]) +
	 2'sd 1 * $signed(input_fmap_5[239:224]) +
	-2'sd 1 * $signed(input_fmap_5[255:240]) +
	-2'sd 1 * $signed(input_fmap_5[271:256]) +
	-2'sd 1 * $signed(input_fmap_5[287:272]) +
	-2'sd 1 * $signed(input_fmap_5[303:288]) +
	 2'sd 1 * $signed(input_fmap_5[319:304]) +
	-2'sd 1 * $signed(input_fmap_5[335:320]) +
	-3'sd 2 * $signed(input_fmap_5[351:336]) +
	-2'sd 1 * $signed(input_fmap_5[367:352]) +
	-2'sd 1 * $signed(input_fmap_5[383:368]) +
	-2'sd 1 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	-2'sd 1 * $signed(input_fmap_0[31:16]) +
	-2'sd 1 * $signed(input_fmap_0[47:32]) +
	-3'sd 3 * $signed(input_fmap_0[63:48]) +
	-4'sd 5 * $signed(input_fmap_0[79:64]) +
	 3'sd 3 * $signed(input_fmap_0[95:80]) +
	-4'sd 7 * $signed(input_fmap_0[127:112]) +
	-4'sd 6 * $signed(input_fmap_0[143:128]) +
	 4'sd 4 * $signed(input_fmap_0[175:160]) +
	-3'sd 2 * $signed(input_fmap_0[191:176]) +
	-5'sd 10 * $signed(input_fmap_0[207:192]) +
	-3'sd 3 * $signed(input_fmap_0[223:208]) +
	 4'sd 4 * $signed(input_fmap_0[239:224]) +
	 3'sd 3 * $signed(input_fmap_0[255:240]) +
	-3'sd 2 * $signed(input_fmap_0[271:256]) +
	-4'sd 5 * $signed(input_fmap_0[287:272]) +
	 3'sd 2 * $signed(input_fmap_0[319:304]) +
	 3'sd 2 * $signed(input_fmap_0[335:320]) +
	-2'sd 1 * $signed(input_fmap_0[351:336]) +
	-3'sd 3 * $signed(input_fmap_0[367:352]) +
	 3'sd 2 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[31:16]) +
	 3'sd 2 * $signed(input_fmap_1[47:32]) +
	 3'sd 3 * $signed(input_fmap_1[63:48]) +
	-3'sd 2 * $signed(input_fmap_1[79:64]) +
	-2'sd 1 * $signed(input_fmap_1[95:80]) +
	 3'sd 3 * $signed(input_fmap_1[127:112]) +
	 3'sd 2 * $signed(input_fmap_1[143:128]) +
	-3'sd 3 * $signed(input_fmap_1[159:144]) +
	-2'sd 1 * $signed(input_fmap_1[175:160]) +
	 2'sd 1 * $signed(input_fmap_1[191:176]) +
	 3'sd 2 * $signed(input_fmap_1[207:192]) +
	 2'sd 1 * $signed(input_fmap_1[223:208]) +
	-3'sd 2 * $signed(input_fmap_1[239:224]) +
	 2'sd 1 * $signed(input_fmap_1[271:256]) +
	 3'sd 2 * $signed(input_fmap_1[287:272]) +
	-3'sd 2 * $signed(input_fmap_1[319:304]) +
	 2'sd 1 * $signed(input_fmap_1[351:336]) +
	 2'sd 1 * $signed(input_fmap_1[367:352]) +
	-2'sd 1 * $signed(input_fmap_1[383:368]) +
	-3'sd 2 * $signed(input_fmap_1[399:384]) +
	 3'sd 2 * $signed(input_fmap_2[63:48]) +
	-2'sd 1 * $signed(input_fmap_2[79:64]) +
	-2'sd 1 * $signed(input_fmap_2[95:80]) +
	 2'sd 1 * $signed(input_fmap_2[127:112]) +
	 3'sd 2 * $signed(input_fmap_2[143:128]) +
	-2'sd 1 * $signed(input_fmap_2[159:144]) +
	 2'sd 1 * $signed(input_fmap_2[207:192]) +
	 3'sd 2 * $signed(input_fmap_2[223:208]) +
	-2'sd 1 * $signed(input_fmap_2[239:224]) +
	 2'sd 1 * $signed(input_fmap_2[287:272]) +
	 2'sd 1 * $signed(input_fmap_2[303:288]) +
	-2'sd 1 * $signed(input_fmap_2[319:304]) +
	 2'sd 1 * $signed(input_fmap_2[335:320]) +
	 2'sd 1 * $signed(input_fmap_2[367:352]) +
	-2'sd 1 * $signed(input_fmap_2[399:384]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	 3'sd 2 * $signed(input_fmap_3[63:48]) +
	-2'sd 1 * $signed(input_fmap_3[95:80]) +
	-2'sd 1 * $signed(input_fmap_3[111:96]) +
	 3'sd 2 * $signed(input_fmap_3[127:112]) +
	 3'sd 3 * $signed(input_fmap_3[143:128]) +
	-3'sd 2 * $signed(input_fmap_3[159:144]) +
	 3'sd 2 * $signed(input_fmap_3[207:192]) +
	 3'sd 2 * $signed(input_fmap_3[223:208]) +
	-2'sd 1 * $signed(input_fmap_3[239:224]) +
	 2'sd 1 * $signed(input_fmap_3[287:272]) +
	 2'sd 1 * $signed(input_fmap_3[303:288]) +
	-2'sd 1 * $signed(input_fmap_3[319:304]) +
	 2'sd 1 * $signed(input_fmap_3[335:320]) +
	 2'sd 1 * $signed(input_fmap_3[367:352]) +
	-2'sd 1 * $signed(input_fmap_3[399:384]) +
	 2'sd 1 * $signed(input_fmap_4[31:16]) +
	-2'sd 1 * $signed(input_fmap_4[63:48]) +
	-2'sd 1 * $signed(input_fmap_4[79:64]) +
	-2'sd 1 * $signed(input_fmap_4[95:80]) +
	 2'sd 1 * $signed(input_fmap_4[127:112]) +
	 2'sd 1 * $signed(input_fmap_4[143:128]) +
	-2'sd 1 * $signed(input_fmap_4[159:144]) +
	-2'sd 1 * $signed(input_fmap_4[175:160]) +
	 2'sd 1 * $signed(input_fmap_4[207:192]) +
	 3'sd 2 * $signed(input_fmap_4[223:208]) +
	 2'sd 1 * $signed(input_fmap_4[303:288]) +
	 2'sd 1 * $signed(input_fmap_4[335:320]) +
	-2'sd 1 * $signed(input_fmap_4[399:384]) +
	 2'sd 1 * $signed(input_fmap_5[63:48]) +
	-2'sd 1 * $signed(input_fmap_5[79:64]) +
	-2'sd 1 * $signed(input_fmap_5[95:80]) +
	 3'sd 2 * $signed(input_fmap_5[127:112]) +
	 3'sd 2 * $signed(input_fmap_5[143:128]) +
	-3'sd 2 * $signed(input_fmap_5[159:144]) +
	-2'sd 1 * $signed(input_fmap_5[175:160]) +
	 2'sd 1 * $signed(input_fmap_5[207:192]) +
	 3'sd 2 * $signed(input_fmap_5[223:208]) +
	-2'sd 1 * $signed(input_fmap_5[239:224]) +
	 2'sd 1 * $signed(input_fmap_5[287:272]) +
	 2'sd 1 * $signed(input_fmap_5[303:288]) +
	-2'sd 1 * $signed(input_fmap_5[319:304]) +
	 2'sd 1 * $signed(input_fmap_5[335:320]) +
	 2'sd 1 * $signed(input_fmap_5[351:336]) +
	 2'sd 1 * $signed(input_fmap_5[367:352]) +
	-2'sd 1 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	 4'sd 4 * $signed(input_fmap_0[15:0]) +
	 3'sd 2 * $signed(input_fmap_0[31:16]) +
	-3'sd 3 * $signed(input_fmap_0[47:32]) +
	-4'sd 7 * $signed(input_fmap_0[63:48]) +
	-3'sd 3 * $signed(input_fmap_0[79:64]) +
	 3'sd 3 * $signed(input_fmap_0[95:80]) +
	 3'sd 2 * $signed(input_fmap_0[111:96]) +
	-2'sd 1 * $signed(input_fmap_0[127:112]) +
	-4'sd 4 * $signed(input_fmap_0[143:128]) +
	-4'sd 5 * $signed(input_fmap_0[159:144]) +
	 3'sd 2 * $signed(input_fmap_0[175:160]) +
	 3'sd 3 * $signed(input_fmap_0[191:176]) +
	 3'sd 3 * $signed(input_fmap_0[207:192]) +
	 3'sd 2 * $signed(input_fmap_0[223:208]) +
	 3'sd 2 * $signed(input_fmap_0[255:240]) +
	-3'sd 2 * $signed(input_fmap_0[271:256]) +
	-3'sd 2 * $signed(input_fmap_0[287:272]) +
	 2'sd 1 * $signed(input_fmap_0[319:304]) +
	 3'sd 2 * $signed(input_fmap_0[335:320]) +
	-2'sd 1 * $signed(input_fmap_0[351:336]) +
	-3'sd 3 * $signed(input_fmap_0[367:352]) +
	-3'sd 2 * $signed(input_fmap_0[383:368]) +
	-3'sd 2 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[31:16]) +
	-3'sd 2 * $signed(input_fmap_1[47:32]) +
	 2'sd 1 * $signed(input_fmap_1[63:48]) +
	 3'sd 2 * $signed(input_fmap_1[79:64]) +
	 2'sd 1 * $signed(input_fmap_1[95:80]) +
	-3'sd 2 * $signed(input_fmap_1[111:96]) +
	-3'sd 3 * $signed(input_fmap_1[127:112]) +
	 2'sd 1 * $signed(input_fmap_1[143:128]) +
	 3'sd 2 * $signed(input_fmap_1[159:144]) +
	 2'sd 1 * $signed(input_fmap_1[175:160]) +
	 2'sd 1 * $signed(input_fmap_1[191:176]) +
	-2'sd 1 * $signed(input_fmap_1[207:192]) +
	-2'sd 1 * $signed(input_fmap_1[223:208]) +
	 2'sd 1 * $signed(input_fmap_1[239:224]) +
	-2'sd 1 * $signed(input_fmap_1[287:272]) +
	-2'sd 1 * $signed(input_fmap_1[303:288]) +
	 2'sd 1 * $signed(input_fmap_1[319:304]) +
	-3'sd 2 * $signed(input_fmap_1[335:320]) +
	-2'sd 1 * $signed(input_fmap_1[351:336]) +
	 2'sd 1 * $signed(input_fmap_1[367:352]) +
	-2'sd 1 * $signed(input_fmap_1[383:368]) +
	-2'sd 1 * $signed(input_fmap_2[31:16]) +
	-3'sd 3 * $signed(input_fmap_2[47:32]) +
	 3'sd 2 * $signed(input_fmap_2[79:64]) +
	-3'sd 3 * $signed(input_fmap_2[127:112]) +
	-2'sd 1 * $signed(input_fmap_2[143:128]) +
	 2'sd 1 * $signed(input_fmap_2[159:144]) +
	 2'sd 1 * $signed(input_fmap_2[175:160]) +
	 3'sd 2 * $signed(input_fmap_2[191:176]) +
	 2'sd 1 * $signed(input_fmap_2[207:192]) +
	-2'sd 1 * $signed(input_fmap_2[223:208]) +
	 2'sd 1 * $signed(input_fmap_2[239:224]) +
	 2'sd 1 * $signed(input_fmap_2[319:304]) +
	-3'sd 2 * $signed(input_fmap_2[335:320]) +
	-3'sd 2 * $signed(input_fmap_2[351:336]) +
	-2'sd 1 * $signed(input_fmap_2[367:352]) +
	-2'sd 1 * $signed(input_fmap_3[15:0]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	-3'sd 3 * $signed(input_fmap_3[47:32]) +
	 2'sd 1 * $signed(input_fmap_3[63:48]) +
	 3'sd 2 * $signed(input_fmap_3[79:64]) +
	-3'sd 3 * $signed(input_fmap_3[127:112]) +
	-2'sd 1 * $signed(input_fmap_3[143:128]) +
	 2'sd 1 * $signed(input_fmap_3[159:144]) +
	 2'sd 1 * $signed(input_fmap_3[175:160]) +
	 3'sd 2 * $signed(input_fmap_3[191:176]) +
	-2'sd 1 * $signed(input_fmap_3[223:208]) +
	 2'sd 1 * $signed(input_fmap_3[239:224]) +
	-2'sd 1 * $signed(input_fmap_3[287:272]) +
	 2'sd 1 * $signed(input_fmap_3[319:304]) +
	-3'sd 2 * $signed(input_fmap_3[335:320]) +
	-3'sd 2 * $signed(input_fmap_3[351:336]) +
	-2'sd 1 * $signed(input_fmap_3[367:352]) +
	-3'sd 2 * $signed(input_fmap_4[31:16]) +
	-3'sd 3 * $signed(input_fmap_4[47:32]) +
	 2'sd 1 * $signed(input_fmap_4[79:64]) +
	 3'sd 2 * $signed(input_fmap_4[95:80]) +
	-4'sd 4 * $signed(input_fmap_4[127:112]) +
	-2'sd 1 * $signed(input_fmap_4[143:128]) +
	 3'sd 2 * $signed(input_fmap_4[159:144]) +
	 3'sd 2 * $signed(input_fmap_4[175:160]) +
	 3'sd 3 * $signed(input_fmap_4[191:176]) +
	-3'sd 2 * $signed(input_fmap_4[223:208]) +
	 2'sd 1 * $signed(input_fmap_4[239:224]) +
	 3'sd 2 * $signed(input_fmap_4[271:256]) +
	 2'sd 1 * $signed(input_fmap_4[287:272]) +
	 3'sd 2 * $signed(input_fmap_4[319:304]) +
	-3'sd 2 * $signed(input_fmap_4[335:320]) +
	-3'sd 2 * $signed(input_fmap_4[351:336]) +
	-2'sd 1 * $signed(input_fmap_4[367:352]) +
	-2'sd 1 * $signed(input_fmap_4[383:368]) +
	-2'sd 1 * $signed(input_fmap_4[399:384]) +
	-2'sd 1 * $signed(input_fmap_5[31:16]) +
	-3'sd 3 * $signed(input_fmap_5[47:32]) +
	 3'sd 2 * $signed(input_fmap_5[79:64]) +
	 2'sd 1 * $signed(input_fmap_5[95:80]) +
	-3'sd 3 * $signed(input_fmap_5[127:112]) +
	-2'sd 1 * $signed(input_fmap_5[143:128]) +
	 3'sd 2 * $signed(input_fmap_5[159:144]) +
	 2'sd 1 * $signed(input_fmap_5[175:160]) +
	 3'sd 2 * $signed(input_fmap_5[191:176]) +
	-2'sd 1 * $signed(input_fmap_5[223:208]) +
	 2'sd 1 * $signed(input_fmap_5[239:224]) +
	 2'sd 1 * $signed(input_fmap_5[271:256]) +
	 2'sd 1 * $signed(input_fmap_5[319:304]) +
	-3'sd 2 * $signed(input_fmap_5[335:320]) +
	-3'sd 2 * $signed(input_fmap_5[351:336]) +
	-2'sd 1 * $signed(input_fmap_5[367:352]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	 3'sd 2 * $signed(input_fmap_0[15:0]) +
	 3'sd 3 * $signed(input_fmap_0[31:16]) +
	 4'sd 5 * $signed(input_fmap_0[47:32]) +
	 4'sd 4 * $signed(input_fmap_0[63:48]) +
	 4'sd 4 * $signed(input_fmap_0[95:80]) +
	 4'sd 5 * $signed(input_fmap_0[111:96]) +
	 3'sd 2 * $signed(input_fmap_0[127:112]) +
	-2'sd 1 * $signed(input_fmap_0[143:128]) +
	-4'sd 4 * $signed(input_fmap_0[159:144]) +
	-2'sd 1 * $signed(input_fmap_0[175:160]) +
	-4'sd 4 * $signed(input_fmap_0[191:176]) +
	-3'sd 2 * $signed(input_fmap_0[207:192]) +
	-2'sd 1 * $signed(input_fmap_0[223:208]) +
	-4'sd 4 * $signed(input_fmap_0[239:224]) +
	 2'sd 1 * $signed(input_fmap_0[255:240]) +
	 4'sd 4 * $signed(input_fmap_0[271:256]) +
	 3'sd 2 * $signed(input_fmap_0[287:272]) +
	-3'sd 2 * $signed(input_fmap_0[303:288]) +
	-4'sd 6 * $signed(input_fmap_0[319:304]) +
	 4'sd 5 * $signed(input_fmap_0[335:320]) +
	 4'sd 5 * $signed(input_fmap_0[351:336]) +
	 2'sd 1 * $signed(input_fmap_0[367:352]) +
	-4'sd 6 * $signed(input_fmap_0[383:368]) +
	-4'sd 4 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[47:32]) +
	-2'sd 1 * $signed(input_fmap_1[63:48]) +
	-2'sd 1 * $signed(input_fmap_1[79:64]) +
	 2'sd 1 * $signed(input_fmap_1[95:80]) +
	 2'sd 1 * $signed(input_fmap_1[111:96]) +
	-2'sd 1 * $signed(input_fmap_1[127:112]) +
	-2'sd 1 * $signed(input_fmap_1[143:128]) +
	-2'sd 1 * $signed(input_fmap_1[175:160]) +
	-2'sd 1 * $signed(input_fmap_1[191:176]) +
	-2'sd 1 * $signed(input_fmap_1[207:192]) +
	 2'sd 1 * $signed(input_fmap_1[223:208]) +
	 2'sd 1 * $signed(input_fmap_1[239:224]) +
	-3'sd 2 * $signed(input_fmap_1[255:240]) +
	-3'sd 2 * $signed(input_fmap_1[271:256]) +
	 2'sd 1 * $signed(input_fmap_1[303:288]) +
	 2'sd 1 * $signed(input_fmap_1[351:336]) +
	 2'sd 1 * $signed(input_fmap_1[367:352]) +
	 2'sd 1 * $signed(input_fmap_1[383:368]) +
	-2'sd 1 * $signed(input_fmap_2[15:0]) +
	 2'sd 1 * $signed(input_fmap_2[31:16]) +
	-2'sd 1 * $signed(input_fmap_2[79:64]) +
	 3'sd 2 * $signed(input_fmap_2[95:80]) +
	 3'sd 2 * $signed(input_fmap_2[111:96]) +
	 2'sd 1 * $signed(input_fmap_2[127:112]) +
	-2'sd 1 * $signed(input_fmap_2[159:144]) +
	-3'sd 2 * $signed(input_fmap_2[175:160]) +
	-2'sd 1 * $signed(input_fmap_2[207:192]) +
	 2'sd 1 * $signed(input_fmap_2[239:224]) +
	-3'sd 2 * $signed(input_fmap_2[255:240]) +
	-3'sd 2 * $signed(input_fmap_2[271:256]) +
	-2'sd 1 * $signed(input_fmap_2[287:272]) +
	 2'sd 1 * $signed(input_fmap_2[303:288]) +
	 3'sd 2 * $signed(input_fmap_2[319:304]) +
	 2'sd 1 * $signed(input_fmap_2[367:352]) +
	 2'sd 1 * $signed(input_fmap_2[399:384]) +
	-2'sd 1 * $signed(input_fmap_3[15:0]) +
	-2'sd 1 * $signed(input_fmap_3[79:64]) +
	 2'sd 1 * $signed(input_fmap_3[95:80]) +
	 2'sd 1 * $signed(input_fmap_3[111:96]) +
	-2'sd 1 * $signed(input_fmap_3[159:144]) +
	-2'sd 1 * $signed(input_fmap_3[175:160]) +
	-2'sd 1 * $signed(input_fmap_3[207:192]) +
	 2'sd 1 * $signed(input_fmap_3[239:224]) +
	-3'sd 2 * $signed(input_fmap_3[255:240]) +
	-3'sd 2 * $signed(input_fmap_3[271:256]) +
	-2'sd 1 * $signed(input_fmap_3[287:272]) +
	 2'sd 1 * $signed(input_fmap_3[303:288]) +
	 3'sd 2 * $signed(input_fmap_3[319:304]) +
	 2'sd 1 * $signed(input_fmap_3[399:384]) +
	-2'sd 1 * $signed(input_fmap_4[15:0]) +
	-2'sd 1 * $signed(input_fmap_4[63:48]) +
	 3'sd 3 * $signed(input_fmap_4[95:80]) +
	 3'sd 2 * $signed(input_fmap_4[111:96]) +
	 3'sd 2 * $signed(input_fmap_4[127:112]) +
	 2'sd 1 * $signed(input_fmap_4[143:128]) +
	 2'sd 1 * $signed(input_fmap_4[191:176]) +
	 2'sd 1 * $signed(input_fmap_4[223:208]) +
	-2'sd 1 * $signed(input_fmap_4[255:240]) +
	-2'sd 1 * $signed(input_fmap_4[271:256]) +
	-2'sd 1 * $signed(input_fmap_4[335:320]) +
	-2'sd 1 * $signed(input_fmap_4[351:336]) +
	 2'sd 1 * $signed(input_fmap_4[399:384]) +
	-2'sd 1 * $signed(input_fmap_5[15:0]) +
	-2'sd 1 * $signed(input_fmap_5[79:64]) +
	 3'sd 2 * $signed(input_fmap_5[95:80]) +
	 3'sd 2 * $signed(input_fmap_5[111:96]) +
	 2'sd 1 * $signed(input_fmap_5[127:112]) +
	-2'sd 1 * $signed(input_fmap_5[175:160]) +
	-3'sd 2 * $signed(input_fmap_5[255:240]) +
	-3'sd 2 * $signed(input_fmap_5[271:256]) +
	 2'sd 1 * $signed(input_fmap_5[319:304]) +
	-2'sd 1 * $signed(input_fmap_5[335:320]) +
	 2'sd 1 * $signed(input_fmap_5[383:368]) +
	 2'sd 1 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	 3'sd 2 * $signed(input_fmap_0[15:0]) +
	 3'sd 2 * $signed(input_fmap_0[31:16]) +
	-2'sd 1 * $signed(input_fmap_0[47:32]) +
	-3'sd 2 * $signed(input_fmap_0[63:48]) +
	-3'sd 2 * $signed(input_fmap_0[79:64]) +
	 4'sd 6 * $signed(input_fmap_0[95:80]) +
	 3'sd 2 * $signed(input_fmap_0[111:96]) +
	-3'sd 3 * $signed(input_fmap_0[127:112]) +
	-3'sd 3 * $signed(input_fmap_0[143:128]) +
	-4'sd 4 * $signed(input_fmap_0[159:144]) +
	 4'sd 4 * $signed(input_fmap_0[175:160]) +
	-2'sd 1 * $signed(input_fmap_0[191:176]) +
	-3'sd 2 * $signed(input_fmap_0[207:192]) +
	-3'sd 3 * $signed(input_fmap_0[223:208]) +
	-4'sd 6 * $signed(input_fmap_0[239:224]) +
	-2'sd 1 * $signed(input_fmap_0[255:240]) +
	-2'sd 1 * $signed(input_fmap_0[271:256]) +
	-3'sd 3 * $signed(input_fmap_0[303:288]) +
	-5'sd 9 * $signed(input_fmap_0[319:304]) +
	-2'sd 1 * $signed(input_fmap_0[335:320]) +
	 3'sd 2 * $signed(input_fmap_0[351:336]) +
	 3'sd 2 * $signed(input_fmap_0[367:352]) +
	-4'sd 4 * $signed(input_fmap_0[383:368]) +
	-4'sd 7 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[15:0]) +
	-2'sd 1 * $signed(input_fmap_1[31:16]) +
	 2'sd 1 * $signed(input_fmap_1[79:64]) +
	-2'sd 1 * $signed(input_fmap_1[111:96]) +
	-3'sd 2 * $signed(input_fmap_1[127:112]) +
	 3'sd 2 * $signed(input_fmap_1[143:128]) +
	 3'sd 3 * $signed(input_fmap_1[159:144]) +
	 3'sd 2 * $signed(input_fmap_1[175:160]) +
	-3'sd 2 * $signed(input_fmap_1[191:176]) +
	-3'sd 3 * $signed(input_fmap_1[207:192]) +
	 3'sd 3 * $signed(input_fmap_1[223:208]) +
	 3'sd 3 * $signed(input_fmap_1[239:224]) +
	 2'sd 1 * $signed(input_fmap_1[255:240]) +
	-3'sd 3 * $signed(input_fmap_1[271:256]) +
	 3'sd 3 * $signed(input_fmap_1[303:288]) +
	 3'sd 2 * $signed(input_fmap_1[319:304]) +
	-2'sd 1 * $signed(input_fmap_1[335:320]) +
	 2'sd 1 * $signed(input_fmap_1[351:336]) +
	 3'sd 3 * $signed(input_fmap_1[367:352]) +
	 3'sd 3 * $signed(input_fmap_1[383:368]) +
	 2'sd 1 * $signed(input_fmap_1[399:384]) +
	-2'sd 1 * $signed(input_fmap_2[47:32]) +
	 2'sd 1 * $signed(input_fmap_2[79:64]) +
	-2'sd 1 * $signed(input_fmap_2[111:96]) +
	-3'sd 3 * $signed(input_fmap_2[127:112]) +
	 3'sd 2 * $signed(input_fmap_2[159:144]) +
	 3'sd 2 * $signed(input_fmap_2[175:160]) +
	-2'sd 1 * $signed(input_fmap_2[191:176]) +
	-3'sd 3 * $signed(input_fmap_2[207:192]) +
	 2'sd 1 * $signed(input_fmap_2[223:208]) +
	 3'sd 2 * $signed(input_fmap_2[239:224]) +
	 2'sd 1 * $signed(input_fmap_2[255:240]) +
	-3'sd 2 * $signed(input_fmap_2[271:256]) +
	-2'sd 1 * $signed(input_fmap_2[287:272]) +
	 3'sd 2 * $signed(input_fmap_2[303:288]) +
	 3'sd 2 * $signed(input_fmap_2[319:304]) +
	-2'sd 1 * $signed(input_fmap_2[335:320]) +
	 3'sd 2 * $signed(input_fmap_2[367:352]) +
	 3'sd 3 * $signed(input_fmap_2[383:368]) +
	 3'sd 2 * $signed(input_fmap_2[399:384]) +
	-2'sd 1 * $signed(input_fmap_3[15:0]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	-2'sd 1 * $signed(input_fmap_3[47:32]) +
	 2'sd 1 * $signed(input_fmap_3[79:64]) +
	 2'sd 1 * $signed(input_fmap_3[95:80]) +
	-3'sd 2 * $signed(input_fmap_3[127:112]) +
	 3'sd 2 * $signed(input_fmap_3[159:144]) +
	 3'sd 2 * $signed(input_fmap_3[175:160]) +
	-2'sd 1 * $signed(input_fmap_3[191:176]) +
	-4'sd 4 * $signed(input_fmap_3[207:192]) +
	 2'sd 1 * $signed(input_fmap_3[223:208]) +
	 3'sd 3 * $signed(input_fmap_3[239:224]) +
	 3'sd 2 * $signed(input_fmap_3[255:240]) +
	-3'sd 2 * $signed(input_fmap_3[271:256]) +
	-2'sd 1 * $signed(input_fmap_3[287:272]) +
	 3'sd 2 * $signed(input_fmap_3[303:288]) +
	 3'sd 2 * $signed(input_fmap_3[319:304]) +
	-2'sd 1 * $signed(input_fmap_3[335:320]) +
	-2'sd 1 * $signed(input_fmap_3[351:336]) +
	 2'sd 1 * $signed(input_fmap_3[367:352]) +
	 3'sd 3 * $signed(input_fmap_3[383:368]) +
	 3'sd 2 * $signed(input_fmap_3[399:384]) +
	-2'sd 1 * $signed(input_fmap_4[31:16]) +
	-2'sd 1 * $signed(input_fmap_4[47:32]) +
	 2'sd 1 * $signed(input_fmap_4[79:64]) +
	-2'sd 1 * $signed(input_fmap_4[111:96]) +
	-3'sd 2 * $signed(input_fmap_4[127:112]) +
	 2'sd 1 * $signed(input_fmap_4[143:128]) +
	 2'sd 1 * $signed(input_fmap_4[159:144]) +
	 2'sd 1 * $signed(input_fmap_4[175:160]) +
	-3'sd 3 * $signed(input_fmap_4[191:176]) +
	-3'sd 3 * $signed(input_fmap_4[207:192]) +
	 2'sd 1 * $signed(input_fmap_4[239:224]) +
	-3'sd 2 * $signed(input_fmap_4[271:256]) +
	-2'sd 1 * $signed(input_fmap_4[287:272]) +
	 2'sd 1 * $signed(input_fmap_4[319:304]) +
	-2'sd 1 * $signed(input_fmap_4[335:320]) +
	-2'sd 1 * $signed(input_fmap_4[351:336]) +
	 2'sd 1 * $signed(input_fmap_4[367:352]) +
	 2'sd 1 * $signed(input_fmap_4[383:368]) +
	 2'sd 1 * $signed(input_fmap_4[399:384]) +
	-2'sd 1 * $signed(input_fmap_5[31:16]) +
	-2'sd 1 * $signed(input_fmap_5[47:32]) +
	 2'sd 1 * $signed(input_fmap_5[79:64]) +
	-2'sd 1 * $signed(input_fmap_5[111:96]) +
	-3'sd 2 * $signed(input_fmap_5[127:112]) +
	 3'sd 2 * $signed(input_fmap_5[159:144]) +
	 2'sd 1 * $signed(input_fmap_5[175:160]) +
	-3'sd 2 * $signed(input_fmap_5[191:176]) +
	-3'sd 3 * $signed(input_fmap_5[207:192]) +
	 3'sd 2 * $signed(input_fmap_5[239:224]) +
	 2'sd 1 * $signed(input_fmap_5[255:240]) +
	-3'sd 2 * $signed(input_fmap_5[271:256]) +
	-2'sd 1 * $signed(input_fmap_5[287:272]) +
	 2'sd 1 * $signed(input_fmap_5[303:288]) +
	 3'sd 2 * $signed(input_fmap_5[319:304]) +
	-2'sd 1 * $signed(input_fmap_5[335:320]) +
	-2'sd 1 * $signed(input_fmap_5[351:336]) +
	 2'sd 1 * $signed(input_fmap_5[367:352]) +
	 3'sd 2 * $signed(input_fmap_5[383:368]) +
	 2'sd 1 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	 3'sd 2 * $signed(input_fmap_0[15:0]) +
	 2'sd 1 * $signed(input_fmap_0[31:16]) +
	-2'sd 1 * $signed(input_fmap_0[47:32]) +
	-2'sd 1 * $signed(input_fmap_0[63:48]) +
	-2'sd 1 * $signed(input_fmap_0[79:64]) +
	 4'sd 4 * $signed(input_fmap_0[95:80]) +
	-3'sd 2 * $signed(input_fmap_0[111:96]) +
	-3'sd 3 * $signed(input_fmap_0[127:112]) +
	-2'sd 1 * $signed(input_fmap_0[143:128]) +
	-2'sd 1 * $signed(input_fmap_0[159:144]) +
	 3'sd 2 * $signed(input_fmap_0[175:160]) +
	-2'sd 1 * $signed(input_fmap_0[191:176]) +
	 2'sd 1 * $signed(input_fmap_0[207:192]) +
	-3'sd 2 * $signed(input_fmap_0[223:208]) +
	-4'sd 5 * $signed(input_fmap_0[239:224]) +
	 2'sd 1 * $signed(input_fmap_0[271:256]) +
	-4'sd 4 * $signed(input_fmap_0[303:288]) +
	-5'sd 9 * $signed(input_fmap_0[319:304]) +
	 2'sd 1 * $signed(input_fmap_0[335:320]) +
	 3'sd 2 * $signed(input_fmap_0[351:336]) +
	 2'sd 1 * $signed(input_fmap_0[367:352]) +
	-4'sd 6 * $signed(input_fmap_0[383:368]) +
	-4'sd 5 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[31:16]) +
	 2'sd 1 * $signed(input_fmap_1[47:32]) +
	 2'sd 1 * $signed(input_fmap_1[63:48]) +
	-3'sd 2 * $signed(input_fmap_1[111:96]) +
	 3'sd 2 * $signed(input_fmap_1[143:128]) +
	 2'sd 1 * $signed(input_fmap_1[159:144]) +
	-2'sd 1 * $signed(input_fmap_1[175:160]) +
	-3'sd 3 * $signed(input_fmap_1[191:176]) +
	 2'sd 1 * $signed(input_fmap_1[207:192]) +
	 3'sd 3 * $signed(input_fmap_1[223:208]) +
	 2'sd 1 * $signed(input_fmap_1[239:224]) +
	-3'sd 2 * $signed(input_fmap_1[255:240]) +
	 3'sd 3 * $signed(input_fmap_1[287:272]) +
	 3'sd 2 * $signed(input_fmap_1[303:288]) +
	-2'sd 1 * $signed(input_fmap_1[335:320]) +
	 2'sd 1 * $signed(input_fmap_1[351:336]) +
	 3'sd 3 * $signed(input_fmap_1[367:352]) +
	 3'sd 2 * $signed(input_fmap_1[383:368]) +
	-2'sd 1 * $signed(input_fmap_2[31:16]) +
	 2'sd 1 * $signed(input_fmap_2[63:48]) +
	 2'sd 1 * $signed(input_fmap_2[79:64]) +
	-3'sd 2 * $signed(input_fmap_2[111:96]) +
	-2'sd 1 * $signed(input_fmap_2[127:112]) +
	 2'sd 1 * $signed(input_fmap_2[143:128]) +
	 2'sd 1 * $signed(input_fmap_2[159:144]) +
	 2'sd 1 * $signed(input_fmap_2[175:160]) +
	-3'sd 3 * $signed(input_fmap_2[191:176]) +
	 3'sd 2 * $signed(input_fmap_2[223:208]) +
	 2'sd 1 * $signed(input_fmap_2[239:224]) +
	-3'sd 2 * $signed(input_fmap_2[271:256]) +
	 2'sd 1 * $signed(input_fmap_2[287:272]) +
	 3'sd 2 * $signed(input_fmap_2[303:288]) +
	 2'sd 1 * $signed(input_fmap_2[319:304]) +
	-2'sd 1 * $signed(input_fmap_2[335:320]) +
	 2'sd 1 * $signed(input_fmap_2[351:336]) +
	 3'sd 2 * $signed(input_fmap_2[367:352]) +
	 3'sd 2 * $signed(input_fmap_2[383:368]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	 2'sd 1 * $signed(input_fmap_3[63:48]) +
	 2'sd 1 * $signed(input_fmap_3[95:80]) +
	-3'sd 2 * $signed(input_fmap_3[111:96]) +
	-2'sd 1 * $signed(input_fmap_3[127:112]) +
	 3'sd 2 * $signed(input_fmap_3[143:128]) +
	 2'sd 1 * $signed(input_fmap_3[159:144]) +
	 2'sd 1 * $signed(input_fmap_3[175:160]) +
	-3'sd 3 * $signed(input_fmap_3[191:176]) +
	-2'sd 1 * $signed(input_fmap_3[207:192]) +
	 3'sd 2 * $signed(input_fmap_3[223:208]) +
	 2'sd 1 * $signed(input_fmap_3[239:224]) +
	-3'sd 2 * $signed(input_fmap_3[271:256]) +
	 3'sd 2 * $signed(input_fmap_3[287:272]) +
	 3'sd 2 * $signed(input_fmap_3[303:288]) +
	 2'sd 1 * $signed(input_fmap_3[319:304]) +
	-2'sd 1 * $signed(input_fmap_3[335:320]) +
	 3'sd 3 * $signed(input_fmap_3[367:352]) +
	 3'sd 2 * $signed(input_fmap_3[383:368]) +
	-2'sd 1 * $signed(input_fmap_4[31:16]) +
	 2'sd 1 * $signed(input_fmap_4[47:32]) +
	 2'sd 1 * $signed(input_fmap_4[63:48]) +
	-2'sd 1 * $signed(input_fmap_4[95:80]) +
	-3'sd 2 * $signed(input_fmap_4[111:96]) +
	 2'sd 1 * $signed(input_fmap_4[143:128]) +
	 2'sd 1 * $signed(input_fmap_4[159:144]) +
	-3'sd 2 * $signed(input_fmap_4[191:176]) +
	 2'sd 1 * $signed(input_fmap_4[223:208]) +
	-2'sd 1 * $signed(input_fmap_4[271:256]) +
	 2'sd 1 * $signed(input_fmap_4[303:288]) +
	 2'sd 1 * $signed(input_fmap_4[319:304]) +
	 2'sd 1 * $signed(input_fmap_4[367:352]) +
	 2'sd 1 * $signed(input_fmap_4[383:368]) +
	-2'sd 1 * $signed(input_fmap_5[31:16]) +
	 2'sd 1 * $signed(input_fmap_5[63:48]) +
	-3'sd 2 * $signed(input_fmap_5[111:96]) +
	-2'sd 1 * $signed(input_fmap_5[127:112]) +
	 2'sd 1 * $signed(input_fmap_5[143:128]) +
	 2'sd 1 * $signed(input_fmap_5[159:144]) +
	 2'sd 1 * $signed(input_fmap_5[175:160]) +
	-3'sd 3 * $signed(input_fmap_5[191:176]) +
	 2'sd 1 * $signed(input_fmap_5[223:208]) +
	 2'sd 1 * $signed(input_fmap_5[239:224]) +
	-3'sd 2 * $signed(input_fmap_5[271:256]) +
	 2'sd 1 * $signed(input_fmap_5[287:272]) +
	 3'sd 2 * $signed(input_fmap_5[303:288]) +
	 2'sd 1 * $signed(input_fmap_5[319:304]) +
	-2'sd 1 * $signed(input_fmap_5[335:320]) +
	 3'sd 2 * $signed(input_fmap_5[367:352]) +
	 3'sd 2 * $signed(input_fmap_5[383:368]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	 3'sd 3 * $signed(input_fmap_0[15:0]) +
	-2'sd 1 * $signed(input_fmap_0[47:32]) +
	-3'sd 2 * $signed(input_fmap_0[79:64]) +
	 2'sd 1 * $signed(input_fmap_0[95:80]) +
	 2'sd 1 * $signed(input_fmap_0[143:128]) +
	 3'sd 2 * $signed(input_fmap_0[159:144]) +
	 2'sd 1 * $signed(input_fmap_0[175:160]) +
	 4'sd 4 * $signed(input_fmap_0[191:176]) +
	 4'sd 4 * $signed(input_fmap_0[207:192]) +
	 3'sd 3 * $signed(input_fmap_0[223:208]) +
	 2'sd 1 * $signed(input_fmap_0[239:224]) +
	 4'sd 4 * $signed(input_fmap_0[255:240]) +
	 4'sd 4 * $signed(input_fmap_0[271:256]) +
	 2'sd 1 * $signed(input_fmap_0[287:272]) +
	-4'sd 4 * $signed(input_fmap_0[303:288]) +
	-4'sd 4 * $signed(input_fmap_0[319:304]) +
	 4'sd 4 * $signed(input_fmap_0[335:320]) +
	-3'sd 2 * $signed(input_fmap_0[351:336]) +
	-4'sd 4 * $signed(input_fmap_0[367:352]) +
	-3'sd 2 * $signed(input_fmap_0[383:368]) +
	-2'sd 1 * $signed(input_fmap_1[47:32]) +
	-3'sd 2 * $signed(input_fmap_1[63:48]) +
	-3'sd 2 * $signed(input_fmap_1[79:64]) +
	-2'sd 1 * $signed(input_fmap_1[95:80]) +
	-3'sd 3 * $signed(input_fmap_1[111:96]) +
	-2'sd 1 * $signed(input_fmap_1[127:112]) +
	-2'sd 1 * $signed(input_fmap_1[143:128]) +
	 2'sd 1 * $signed(input_fmap_1[159:144]) +
	 3'sd 2 * $signed(input_fmap_1[207:192]) +
	 3'sd 2 * $signed(input_fmap_1[223:208]) +
	 2'sd 1 * $signed(input_fmap_1[239:224]) +
	 3'sd 2 * $signed(input_fmap_1[271:256]) +
	 2'sd 1 * $signed(input_fmap_1[287:272]) +
	-2'sd 1 * $signed(input_fmap_1[319:304]) +
	 2'sd 1 * $signed(input_fmap_1[351:336]) +
	-2'sd 1 * $signed(input_fmap_1[383:368]) +
	-3'sd 2 * $signed(input_fmap_1[399:384]) +
	-2'sd 1 * $signed(input_fmap_2[31:16]) +
	-2'sd 1 * $signed(input_fmap_2[47:32]) +
	-3'sd 2 * $signed(input_fmap_2[63:48]) +
	-3'sd 2 * $signed(input_fmap_2[79:64]) +
	-3'sd 2 * $signed(input_fmap_2[111:96]) +
	-3'sd 2 * $signed(input_fmap_2[127:112]) +
	-2'sd 1 * $signed(input_fmap_2[143:128]) +
	 2'sd 1 * $signed(input_fmap_2[159:144]) +
	 2'sd 1 * $signed(input_fmap_2[207:192]) +
	 3'sd 2 * $signed(input_fmap_2[223:208]) +
	 3'sd 2 * $signed(input_fmap_2[239:224]) +
	 2'sd 1 * $signed(input_fmap_2[271:256]) +
	 2'sd 1 * $signed(input_fmap_2[287:272]) +
	 2'sd 1 * $signed(input_fmap_2[303:288]) +
	 2'sd 1 * $signed(input_fmap_2[351:336]) +
	-3'sd 2 * $signed(input_fmap_2[399:384]) +
	-2'sd 1 * $signed(input_fmap_3[47:32]) +
	-3'sd 2 * $signed(input_fmap_3[63:48]) +
	-3'sd 2 * $signed(input_fmap_3[79:64]) +
	-3'sd 2 * $signed(input_fmap_3[111:96]) +
	-3'sd 2 * $signed(input_fmap_3[127:112]) +
	-2'sd 1 * $signed(input_fmap_3[143:128]) +
	-2'sd 1 * $signed(input_fmap_3[191:176]) +
	 2'sd 1 * $signed(input_fmap_3[223:208]) +
	 2'sd 1 * $signed(input_fmap_3[239:224]) +
	 2'sd 1 * $signed(input_fmap_3[287:272]) +
	 2'sd 1 * $signed(input_fmap_3[303:288]) +
	 2'sd 1 * $signed(input_fmap_3[351:336]) +
	-2'sd 1 * $signed(input_fmap_3[383:368]) +
	-3'sd 2 * $signed(input_fmap_3[399:384]) +
	-2'sd 1 * $signed(input_fmap_4[63:48]) +
	-2'sd 1 * $signed(input_fmap_4[79:64]) +
	-2'sd 1 * $signed(input_fmap_4[111:96]) +
	-2'sd 1 * $signed(input_fmap_4[127:112]) +
	-2'sd 1 * $signed(input_fmap_4[143:128]) +
	 2'sd 1 * $signed(input_fmap_4[175:160]) +
	 2'sd 1 * $signed(input_fmap_4[223:208]) +
	 2'sd 1 * $signed(input_fmap_4[239:224]) +
	 2'sd 1 * $signed(input_fmap_4[255:240]) +
	 2'sd 1 * $signed(input_fmap_4[271:256]) +
	 2'sd 1 * $signed(input_fmap_4[287:272]) +
	 2'sd 1 * $signed(input_fmap_4[303:288]) +
	-2'sd 1 * $signed(input_fmap_4[399:384]) +
	-3'sd 2 * $signed(input_fmap_5[63:48]) +
	-2'sd 1 * $signed(input_fmap_5[79:64]) +
	-3'sd 2 * $signed(input_fmap_5[111:96]) +
	-2'sd 1 * $signed(input_fmap_5[127:112]) +
	-2'sd 1 * $signed(input_fmap_5[143:128]) +
	 2'sd 1 * $signed(input_fmap_5[207:192]) +
	 2'sd 1 * $signed(input_fmap_5[223:208]) +
	 3'sd 2 * $signed(input_fmap_5[239:224]) +
	 2'sd 1 * $signed(input_fmap_5[255:240]) +
	 2'sd 1 * $signed(input_fmap_5[271:256]) +
	 2'sd 1 * $signed(input_fmap_5[287:272]) +
	 2'sd 1 * $signed(input_fmap_5[303:288]) +
	 2'sd 1 * $signed(input_fmap_5[351:336]) +
	-2'sd 1 * $signed(input_fmap_5[383:368]) +
	-2'sd 1 * $signed(input_fmap_5[399:384]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	-2'sd 1 * $signed(input_fmap_0[15:0]) +
	 2'sd 1 * $signed(input_fmap_0[79:64]) +
	-3'sd 2 * $signed(input_fmap_0[95:80]) +
	-3'sd 3 * $signed(input_fmap_0[111:96]) +
	-3'sd 2 * $signed(input_fmap_0[127:112]) +
	-2'sd 1 * $signed(input_fmap_0[143:128]) +
	-3'sd 2 * $signed(input_fmap_0[159:144]) +
	-3'sd 3 * $signed(input_fmap_0[175:160]) +
	-4'sd 6 * $signed(input_fmap_0[191:176]) +
	-2'sd 1 * $signed(input_fmap_0[207:192]) +
	 4'sd 6 * $signed(input_fmap_0[223:208]) +
	 4'sd 4 * $signed(input_fmap_0[239:224]) +
	-3'sd 3 * $signed(input_fmap_0[255:240]) +
	-4'sd 7 * $signed(input_fmap_0[271:256]) +
	-4'sd 5 * $signed(input_fmap_0[287:272]) +
	 3'sd 3 * $signed(input_fmap_0[303:288]) +
	 4'sd 4 * $signed(input_fmap_0[319:304]) +
	 2'sd 1 * $signed(input_fmap_0[335:320]) +
	-3'sd 2 * $signed(input_fmap_0[351:336]) +
	-4'sd 4 * $signed(input_fmap_0[367:352]) +
	-3'sd 3 * $signed(input_fmap_0[383:368]) +
	-2'sd 1 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[15:0]) +
	-2'sd 1 * $signed(input_fmap_1[31:16]) +
	-2'sd 1 * $signed(input_fmap_1[79:64]) +
	 2'sd 1 * $signed(input_fmap_1[95:80]) +
	 3'sd 2 * $signed(input_fmap_1[111:96]) +
	-2'sd 1 * $signed(input_fmap_1[143:128]) +
	-3'sd 2 * $signed(input_fmap_1[159:144]) +
	 3'sd 3 * $signed(input_fmap_1[191:176]) +
	 3'sd 2 * $signed(input_fmap_1[207:192]) +
	-3'sd 2 * $signed(input_fmap_1[223:208]) +
	-3'sd 3 * $signed(input_fmap_1[239:224]) +
	-3'sd 2 * $signed(input_fmap_1[255:240]) +
	 3'sd 2 * $signed(input_fmap_1[271:256]) +
	 3'sd 2 * $signed(input_fmap_1[287:272]) +
	-2'sd 1 * $signed(input_fmap_1[303:288]) +
	-3'sd 2 * $signed(input_fmap_1[319:304]) +
	-3'sd 2 * $signed(input_fmap_1[335:320]) +
	-2'sd 1 * $signed(input_fmap_1[351:336]) +
	-3'sd 2 * $signed(input_fmap_1[399:384]) +
	-2'sd 1 * $signed(input_fmap_2[47:32]) +
	-2'sd 1 * $signed(input_fmap_2[79:64]) +
	 3'sd 3 * $signed(input_fmap_2[111:96]) +
	-3'sd 3 * $signed(input_fmap_2[143:128]) +
	-3'sd 2 * $signed(input_fmap_2[159:144]) +
	 3'sd 3 * $signed(input_fmap_2[191:176]) +
	 3'sd 3 * $signed(input_fmap_2[207:192]) +
	 2'sd 1 * $signed(input_fmap_2[223:208]) +
	-3'sd 2 * $signed(input_fmap_2[239:224]) +
	-3'sd 2 * $signed(input_fmap_2[255:240]) +
	 3'sd 3 * $signed(input_fmap_2[287:272]) +
	 3'sd 2 * $signed(input_fmap_2[303:288]) +
	-2'sd 1 * $signed(input_fmap_2[335:320]) +
	-3'sd 2 * $signed(input_fmap_2[351:336]) +
	-2'sd 1 * $signed(input_fmap_2[367:352]) +
	-2'sd 1 * $signed(input_fmap_2[399:384]) +
	-2'sd 1 * $signed(input_fmap_3[15:0]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	-2'sd 1 * $signed(input_fmap_3[47:32]) +
	-2'sd 1 * $signed(input_fmap_3[79:64]) +
	-2'sd 1 * $signed(input_fmap_3[95:80]) +
	 3'sd 2 * $signed(input_fmap_3[111:96]) +
	 2'sd 1 * $signed(input_fmap_3[127:112]) +
	-3'sd 2 * $signed(input_fmap_3[143:128]) +
	-3'sd 2 * $signed(input_fmap_3[159:144]) +
	-2'sd 1 * $signed(input_fmap_3[175:160]) +
	 3'sd 3 * $signed(input_fmap_3[191:176]) +
	 3'sd 3 * $signed(input_fmap_3[207:192]) +
	-3'sd 2 * $signed(input_fmap_3[239:224]) +
	-3'sd 2 * $signed(input_fmap_3[255:240]) +
	 3'sd 3 * $signed(input_fmap_3[287:272]) +
	 2'sd 1 * $signed(input_fmap_3[303:288]) +
	-2'sd 1 * $signed(input_fmap_3[319:304]) +
	-2'sd 1 * $signed(input_fmap_3[335:320]) +
	-3'sd 2 * $signed(input_fmap_3[351:336]) +
	-2'sd 1 * $signed(input_fmap_3[367:352]) +
	-2'sd 1 * $signed(input_fmap_3[399:384]) +
	 2'sd 1 * $signed(input_fmap_4[15:0]) +
	-2'sd 1 * $signed(input_fmap_4[31:16]) +
	-3'sd 2 * $signed(input_fmap_4[47:32]) +
	-2'sd 1 * $signed(input_fmap_4[63:48]) +
	-2'sd 1 * $signed(input_fmap_4[79:64]) +
	 2'sd 1 * $signed(input_fmap_4[95:80]) +
	 3'sd 3 * $signed(input_fmap_4[111:96]) +
	-2'sd 1 * $signed(input_fmap_4[127:112]) +
	-3'sd 3 * $signed(input_fmap_4[143:128]) +
	-2'sd 1 * $signed(input_fmap_4[159:144]) +
	 4'sd 5 * $signed(input_fmap_4[191:176]) +
	 4'sd 4 * $signed(input_fmap_4[207:192]) +
	-3'sd 3 * $signed(input_fmap_4[239:224]) +
	-3'sd 2 * $signed(input_fmap_4[255:240]) +
	 2'sd 1 * $signed(input_fmap_4[271:256]) +
	 4'sd 5 * $signed(input_fmap_4[287:272]) +
	 4'sd 4 * $signed(input_fmap_4[303:288]) +
	-2'sd 1 * $signed(input_fmap_4[335:320]) +
	-3'sd 3 * $signed(input_fmap_4[351:336]) +
	 3'sd 2 * $signed(input_fmap_4[383:368]) +
	-2'sd 1 * $signed(input_fmap_5[31:16]) +
	-2'sd 1 * $signed(input_fmap_5[47:32]) +
	-2'sd 1 * $signed(input_fmap_5[79:64]) +
	 2'sd 1 * $signed(input_fmap_5[95:80]) +
	 3'sd 3 * $signed(input_fmap_5[111:96]) +
	-3'sd 2 * $signed(input_fmap_5[143:128]) +
	-2'sd 1 * $signed(input_fmap_5[159:144]) +
	 4'sd 4 * $signed(input_fmap_5[191:176]) +
	 3'sd 3 * $signed(input_fmap_5[207:192]) +
	-3'sd 3 * $signed(input_fmap_5[239:224]) +
	-2'sd 1 * $signed(input_fmap_5[255:240]) +
	 2'sd 1 * $signed(input_fmap_5[271:256]) +
	 4'sd 4 * $signed(input_fmap_5[287:272]) +
	 3'sd 3 * $signed(input_fmap_5[303:288]) +
	-2'sd 1 * $signed(input_fmap_5[319:304]) +
	-2'sd 1 * $signed(input_fmap_5[335:320]) +
	-3'sd 2 * $signed(input_fmap_5[351:336]) +
	-2'sd 1 * $signed(input_fmap_5[367:352]) +
	 2'sd 1 * $signed(input_fmap_5[383:368]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	 3'sd 2 * $signed(input_fmap_0[15:0]) +
	 3'sd 2 * $signed(input_fmap_0[31:16]) +
	-3'sd 2 * $signed(input_fmap_0[63:48]) +
	-2'sd 1 * $signed(input_fmap_0[79:64]) +
	 2'sd 1 * $signed(input_fmap_0[95:80]) +
	 3'sd 2 * $signed(input_fmap_0[111:96]) +
	-2'sd 1 * $signed(input_fmap_0[127:112]) +
	-3'sd 2 * $signed(input_fmap_0[143:128]) +
	-3'sd 3 * $signed(input_fmap_0[159:144]) +
	 3'sd 3 * $signed(input_fmap_0[175:160]) +
	-3'sd 2 * $signed(input_fmap_0[191:176]) +
	-4'sd 5 * $signed(input_fmap_0[207:192]) +
	-3'sd 2 * $signed(input_fmap_0[223:208]) +
	-2'sd 1 * $signed(input_fmap_0[239:224]) +
	-5'sd 8 * $signed(input_fmap_0[271:256]) +
	-4'sd 4 * $signed(input_fmap_0[287:272]) +
	 3'sd 2 * $signed(input_fmap_0[303:288]) +
	 4'sd 5 * $signed(input_fmap_0[319:304]) +
	-4'sd 5 * $signed(input_fmap_0[335:320]) +
	-4'sd 4 * $signed(input_fmap_0[351:336]) +
	 2'sd 1 * $signed(input_fmap_0[367:352]) +
	 4'sd 4 * $signed(input_fmap_0[383:368]) +
	 4'sd 6 * $signed(input_fmap_0[399:384]) +
	-2'sd 1 * $signed(input_fmap_1[15:0]) +
	-2'sd 1 * $signed(input_fmap_1[31:16]) +
	-2'sd 1 * $signed(input_fmap_1[47:32]) +
	 2'sd 1 * $signed(input_fmap_1[63:48]) +
	 3'sd 3 * $signed(input_fmap_1[79:64]) +
	 3'sd 2 * $signed(input_fmap_1[111:96]) +
	 2'sd 1 * $signed(input_fmap_1[143:128]) +
	 3'sd 2 * $signed(input_fmap_1[159:144]) +
	 3'sd 3 * $signed(input_fmap_1[175:160]) +
	 3'sd 2 * $signed(input_fmap_1[191:176]) +
	-2'sd 1 * $signed(input_fmap_1[207:192]) +
	 3'sd 3 * $signed(input_fmap_1[255:240]) +
	-3'sd 2 * $signed(input_fmap_1[287:272]) +
	-2'sd 1 * $signed(input_fmap_1[319:304]) +
	 2'sd 1 * $signed(input_fmap_1[335:320]) +
	-3'sd 2 * $signed(input_fmap_1[351:336]) +
	-3'sd 2 * $signed(input_fmap_1[399:384]) +
	-2'sd 1 * $signed(input_fmap_2[15:0]) +
	-2'sd 1 * $signed(input_fmap_2[31:16]) +
	-2'sd 1 * $signed(input_fmap_2[47:32]) +
	 3'sd 2 * $signed(input_fmap_2[79:64]) +
	 2'sd 1 * $signed(input_fmap_2[111:96]) +
	-2'sd 1 * $signed(input_fmap_2[143:128]) +
	 2'sd 1 * $signed(input_fmap_2[159:144]) +
	 2'sd 1 * $signed(input_fmap_2[175:160]) +
	 3'sd 2 * $signed(input_fmap_2[191:176]) +
	-2'sd 1 * $signed(input_fmap_2[223:208]) +
	 2'sd 1 * $signed(input_fmap_2[255:240]) +
	-2'sd 1 * $signed(input_fmap_2[287:272]) +
	-2'sd 1 * $signed(input_fmap_2[303:288]) +
	 2'sd 1 * $signed(input_fmap_2[335:320]) +
	-2'sd 1 * $signed(input_fmap_2[351:336]) +
	-2'sd 1 * $signed(input_fmap_2[367:352]) +
	-2'sd 1 * $signed(input_fmap_3[15:0]) +
	-2'sd 1 * $signed(input_fmap_3[31:16]) +
	-3'sd 2 * $signed(input_fmap_3[47:32]) +
	 3'sd 2 * $signed(input_fmap_3[79:64]) +
	-2'sd 1 * $signed(input_fmap_3[95:80]) +
	 2'sd 1 * $signed(input_fmap_3[111:96]) +
	-2'sd 1 * $signed(input_fmap_3[143:128]) +
	 3'sd 2 * $signed(input_fmap_3[159:144]) +
	 2'sd 1 * $signed(input_fmap_3[175:160]) +
	 3'sd 2 * $signed(input_fmap_3[191:176]) +
	-2'sd 1 * $signed(input_fmap_3[223:208]) +
	 3'sd 2 * $signed(input_fmap_3[255:240]) +
	-3'sd 2 * $signed(input_fmap_3[287:272]) +
	 2'sd 1 * $signed(input_fmap_3[335:320]) +
	-2'sd 1 * $signed(input_fmap_3[351:336]) +
	-2'sd 1 * $signed(input_fmap_3[367:352]) +
	 2'sd 1 * $signed(input_fmap_3[383:368]) +
	-2'sd 1 * $signed(input_fmap_3[399:384]) +
	 2'sd 1 * $signed(input_fmap_4[15:0]) +
	-3'sd 2 * $signed(input_fmap_4[47:32]) +
	 3'sd 2 * $signed(input_fmap_4[79:64]) +
	 2'sd 1 * $signed(input_fmap_4[95:80]) +
	-3'sd 2 * $signed(input_fmap_4[127:112]) +
	-2'sd 1 * $signed(input_fmap_4[143:128]) +
	 2'sd 1 * $signed(input_fmap_4[159:144]) +
	-2'sd 1 * $signed(input_fmap_4[207:192]) +
	-2'sd 1 * $signed(input_fmap_4[223:208]) +
	-2'sd 1 * $signed(input_fmap_4[239:224]) +
	-2'sd 1 * $signed(input_fmap_4[255:240]) +
	-2'sd 1 * $signed(input_fmap_4[287:272]) +
	-2'sd 1 * $signed(input_fmap_4[303:288]) +
	-2'sd 1 * $signed(input_fmap_4[319:304]) +
	-2'sd 1 * $signed(input_fmap_4[367:352]) +
	-2'sd 1 * $signed(input_fmap_5[31:16]) +
	-3'sd 2 * $signed(input_fmap_5[47:32]) +
	 3'sd 2 * $signed(input_fmap_5[79:64]) +
	 2'sd 1 * $signed(input_fmap_5[111:96]) +
	-2'sd 1 * $signed(input_fmap_5[127:112]) +
	-2'sd 1 * $signed(input_fmap_5[143:128]) +
	 2'sd 1 * $signed(input_fmap_5[159:144]) +
	 2'sd 1 * $signed(input_fmap_5[175:160]) +
	 2'sd 1 * $signed(input_fmap_5[191:176]) +
	 2'sd 1 * $signed(input_fmap_5[255:240]) +
	-2'sd 1 * $signed(input_fmap_5[287:272]) +
	-2'sd 1 * $signed(input_fmap_5[303:288]) +
	-2'sd 1 * $signed(input_fmap_5[319:304]) +
	 2'sd 1 * $signed(input_fmap_5[335:320]) +
	-2'sd 1 * $signed(input_fmap_5[351:336]) +
	-2'sd 1 * $signed(input_fmap_5[367:352]) +
	-2'sd 1 * $signed(input_fmap_5[399:384]);

logic [15:0] relu_0;
assign relu_0[15:0] = (conv_mac_0[31]==0) ? {{conv_mac_0[31],conv_mac_0[18:4]}} : '0;
logic [15:0] relu_1;
assign relu_1[15:0] = (conv_mac_1[31]==0) ? {{conv_mac_1[31],conv_mac_1[18:4]}} : '0;
logic [15:0] relu_2;
assign relu_2[15:0] = (conv_mac_2[31]==0) ? {{conv_mac_2[31],conv_mac_2[18:4]}} : '0;
logic [15:0] relu_3;
assign relu_3[15:0] = (conv_mac_3[31]==0) ? {{conv_mac_3[31],conv_mac_3[18:4]}} : '0;
logic [15:0] relu_4;
assign relu_4[15:0] = (conv_mac_4[31]==0) ? {{conv_mac_4[31],conv_mac_4[18:4]}} : '0;
logic [15:0] relu_5;
assign relu_5[15:0] = (conv_mac_5[31]==0) ? {{conv_mac_5[31],conv_mac_5[18:4]}} : '0;
logic [15:0] relu_6;
assign relu_6[15:0] = (conv_mac_6[31]==0) ? {{conv_mac_6[31],conv_mac_6[18:4]}} : '0;
logic [15:0] relu_7;
assign relu_7[15:0] = (conv_mac_7[31]==0) ? {{conv_mac_7[31],conv_mac_7[18:4]}} : '0;
logic [15:0] relu_8;
assign relu_8[15:0] = (conv_mac_8[31]==0) ? {{conv_mac_8[31],conv_mac_8[18:4]}} : '0;
logic [15:0] relu_9;
assign relu_9[15:0] = (conv_mac_9[31]==0) ? {{conv_mac_9[31],conv_mac_9[18:4]}} : '0;
logic [15:0] relu_10;
assign relu_10[15:0] = (conv_mac_10[31]==0) ? {{conv_mac_10[31],conv_mac_10[18:4]}} : '0;
logic [15:0] relu_11;
assign relu_11[15:0] = (conv_mac_11[31]==0) ? {{conv_mac_11[31],conv_mac_11[18:4]}} : '0;
logic [15:0] relu_12;
assign relu_12[15:0] = (conv_mac_12[31]==0) ? {{conv_mac_12[31],conv_mac_12[18:4]}} : '0;
logic [15:0] relu_13;
assign relu_13[15:0] = (conv_mac_13[31]==0) ? {{conv_mac_13[31],conv_mac_13[18:4]}} : '0;
logic [15:0] relu_14;
assign relu_14[15:0] = (conv_mac_14[31]==0) ? {{conv_mac_14[31],conv_mac_14[18:4]}} : '0;
logic [15:0] relu_15;
assign relu_15[15:0] = (conv_mac_15[31]==0) ? {{conv_mac_15[31],conv_mac_15[18:4]}} : '0;

assign output_act = {
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
