module conv14_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [2048-1:0] input_act,
    output logic [2048-1:0] output_act,
    output logic ready
);

logic [2048-1:0] input_act_ff;
always_ff @(posedge clk or negedge rstn) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
        ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
        ready <= valid;
    end
end

logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];
logic [7:0] input_fmap_64;
assign input_fmap_64 = input_act_ff[519:512];
logic [7:0] input_fmap_65;
assign input_fmap_65 = input_act_ff[527:520];
logic [7:0] input_fmap_66;
assign input_fmap_66 = input_act_ff[535:528];
logic [7:0] input_fmap_67;
assign input_fmap_67 = input_act_ff[543:536];
logic [7:0] input_fmap_68;
assign input_fmap_68 = input_act_ff[551:544];
logic [7:0] input_fmap_69;
assign input_fmap_69 = input_act_ff[559:552];
logic [7:0] input_fmap_70;
assign input_fmap_70 = input_act_ff[567:560];
logic [7:0] input_fmap_71;
assign input_fmap_71 = input_act_ff[575:568];
logic [7:0] input_fmap_72;
assign input_fmap_72 = input_act_ff[583:576];
logic [7:0] input_fmap_73;
assign input_fmap_73 = input_act_ff[591:584];
logic [7:0] input_fmap_74;
assign input_fmap_74 = input_act_ff[599:592];
logic [7:0] input_fmap_75;
assign input_fmap_75 = input_act_ff[607:600];
logic [7:0] input_fmap_76;
assign input_fmap_76 = input_act_ff[615:608];
logic [7:0] input_fmap_77;
assign input_fmap_77 = input_act_ff[623:616];
logic [7:0] input_fmap_78;
assign input_fmap_78 = input_act_ff[631:624];
logic [7:0] input_fmap_79;
assign input_fmap_79 = input_act_ff[639:632];
logic [7:0] input_fmap_80;
assign input_fmap_80 = input_act_ff[647:640];
logic [7:0] input_fmap_81;
assign input_fmap_81 = input_act_ff[655:648];
logic [7:0] input_fmap_82;
assign input_fmap_82 = input_act_ff[663:656];
logic [7:0] input_fmap_83;
assign input_fmap_83 = input_act_ff[671:664];
logic [7:0] input_fmap_84;
assign input_fmap_84 = input_act_ff[679:672];
logic [7:0] input_fmap_85;
assign input_fmap_85 = input_act_ff[687:680];
logic [7:0] input_fmap_86;
assign input_fmap_86 = input_act_ff[695:688];
logic [7:0] input_fmap_87;
assign input_fmap_87 = input_act_ff[703:696];
logic [7:0] input_fmap_88;
assign input_fmap_88 = input_act_ff[711:704];
logic [7:0] input_fmap_89;
assign input_fmap_89 = input_act_ff[719:712];
logic [7:0] input_fmap_90;
assign input_fmap_90 = input_act_ff[727:720];
logic [7:0] input_fmap_91;
assign input_fmap_91 = input_act_ff[735:728];
logic [7:0] input_fmap_92;
assign input_fmap_92 = input_act_ff[743:736];
logic [7:0] input_fmap_93;
assign input_fmap_93 = input_act_ff[751:744];
logic [7:0] input_fmap_94;
assign input_fmap_94 = input_act_ff[759:752];
logic [7:0] input_fmap_95;
assign input_fmap_95 = input_act_ff[767:760];
logic [7:0] input_fmap_96;
assign input_fmap_96 = input_act_ff[775:768];
logic [7:0] input_fmap_97;
assign input_fmap_97 = input_act_ff[783:776];
logic [7:0] input_fmap_98;
assign input_fmap_98 = input_act_ff[791:784];
logic [7:0] input_fmap_99;
assign input_fmap_99 = input_act_ff[799:792];
logic [7:0] input_fmap_100;
assign input_fmap_100 = input_act_ff[807:800];
logic [7:0] input_fmap_101;
assign input_fmap_101 = input_act_ff[815:808];
logic [7:0] input_fmap_102;
assign input_fmap_102 = input_act_ff[823:816];
logic [7:0] input_fmap_103;
assign input_fmap_103 = input_act_ff[831:824];
logic [7:0] input_fmap_104;
assign input_fmap_104 = input_act_ff[839:832];
logic [7:0] input_fmap_105;
assign input_fmap_105 = input_act_ff[847:840];
logic [7:0] input_fmap_106;
assign input_fmap_106 = input_act_ff[855:848];
logic [7:0] input_fmap_107;
assign input_fmap_107 = input_act_ff[863:856];
logic [7:0] input_fmap_108;
assign input_fmap_108 = input_act_ff[871:864];
logic [7:0] input_fmap_109;
assign input_fmap_109 = input_act_ff[879:872];
logic [7:0] input_fmap_110;
assign input_fmap_110 = input_act_ff[887:880];
logic [7:0] input_fmap_111;
assign input_fmap_111 = input_act_ff[895:888];
logic [7:0] input_fmap_112;
assign input_fmap_112 = input_act_ff[903:896];
logic [7:0] input_fmap_113;
assign input_fmap_113 = input_act_ff[911:904];
logic [7:0] input_fmap_114;
assign input_fmap_114 = input_act_ff[919:912];
logic [7:0] input_fmap_115;
assign input_fmap_115 = input_act_ff[927:920];
logic [7:0] input_fmap_116;
assign input_fmap_116 = input_act_ff[935:928];
logic [7:0] input_fmap_117;
assign input_fmap_117 = input_act_ff[943:936];
logic [7:0] input_fmap_118;
assign input_fmap_118 = input_act_ff[951:944];
logic [7:0] input_fmap_119;
assign input_fmap_119 = input_act_ff[959:952];
logic [7:0] input_fmap_120;
assign input_fmap_120 = input_act_ff[967:960];
logic [7:0] input_fmap_121;
assign input_fmap_121 = input_act_ff[975:968];
logic [7:0] input_fmap_122;
assign input_fmap_122 = input_act_ff[983:976];
logic [7:0] input_fmap_123;
assign input_fmap_123 = input_act_ff[991:984];
logic [7:0] input_fmap_124;
assign input_fmap_124 = input_act_ff[999:992];
logic [7:0] input_fmap_125;
assign input_fmap_125 = input_act_ff[1007:1000];
logic [7:0] input_fmap_126;
assign input_fmap_126 = input_act_ff[1015:1008];
logic [7:0] input_fmap_127;
assign input_fmap_127 = input_act_ff[1023:1016];
logic [7:0] input_fmap_128;
assign input_fmap_128 = input_act_ff[1031:1024];
logic [7:0] input_fmap_129;
assign input_fmap_129 = input_act_ff[1039:1032];
logic [7:0] input_fmap_130;
assign input_fmap_130 = input_act_ff[1047:1040];
logic [7:0] input_fmap_131;
assign input_fmap_131 = input_act_ff[1055:1048];
logic [7:0] input_fmap_132;
assign input_fmap_132 = input_act_ff[1063:1056];
logic [7:0] input_fmap_133;
assign input_fmap_133 = input_act_ff[1071:1064];
logic [7:0] input_fmap_134;
assign input_fmap_134 = input_act_ff[1079:1072];
logic [7:0] input_fmap_135;
assign input_fmap_135 = input_act_ff[1087:1080];
logic [7:0] input_fmap_136;
assign input_fmap_136 = input_act_ff[1095:1088];
logic [7:0] input_fmap_137;
assign input_fmap_137 = input_act_ff[1103:1096];
logic [7:0] input_fmap_138;
assign input_fmap_138 = input_act_ff[1111:1104];
logic [7:0] input_fmap_139;
assign input_fmap_139 = input_act_ff[1119:1112];
logic [7:0] input_fmap_140;
assign input_fmap_140 = input_act_ff[1127:1120];
logic [7:0] input_fmap_141;
assign input_fmap_141 = input_act_ff[1135:1128];
logic [7:0] input_fmap_142;
assign input_fmap_142 = input_act_ff[1143:1136];
logic [7:0] input_fmap_143;
assign input_fmap_143 = input_act_ff[1151:1144];
logic [7:0] input_fmap_144;
assign input_fmap_144 = input_act_ff[1159:1152];
logic [7:0] input_fmap_145;
assign input_fmap_145 = input_act_ff[1167:1160];
logic [7:0] input_fmap_146;
assign input_fmap_146 = input_act_ff[1175:1168];
logic [7:0] input_fmap_147;
assign input_fmap_147 = input_act_ff[1183:1176];
logic [7:0] input_fmap_148;
assign input_fmap_148 = input_act_ff[1191:1184];
logic [7:0] input_fmap_149;
assign input_fmap_149 = input_act_ff[1199:1192];
logic [7:0] input_fmap_150;
assign input_fmap_150 = input_act_ff[1207:1200];
logic [7:0] input_fmap_151;
assign input_fmap_151 = input_act_ff[1215:1208];
logic [7:0] input_fmap_152;
assign input_fmap_152 = input_act_ff[1223:1216];
logic [7:0] input_fmap_153;
assign input_fmap_153 = input_act_ff[1231:1224];
logic [7:0] input_fmap_154;
assign input_fmap_154 = input_act_ff[1239:1232];
logic [7:0] input_fmap_155;
assign input_fmap_155 = input_act_ff[1247:1240];
logic [7:0] input_fmap_156;
assign input_fmap_156 = input_act_ff[1255:1248];
logic [7:0] input_fmap_157;
assign input_fmap_157 = input_act_ff[1263:1256];
logic [7:0] input_fmap_158;
assign input_fmap_158 = input_act_ff[1271:1264];
logic [7:0] input_fmap_159;
assign input_fmap_159 = input_act_ff[1279:1272];
logic [7:0] input_fmap_160;
assign input_fmap_160 = input_act_ff[1287:1280];
logic [7:0] input_fmap_161;
assign input_fmap_161 = input_act_ff[1295:1288];
logic [7:0] input_fmap_162;
assign input_fmap_162 = input_act_ff[1303:1296];
logic [7:0] input_fmap_163;
assign input_fmap_163 = input_act_ff[1311:1304];
logic [7:0] input_fmap_164;
assign input_fmap_164 = input_act_ff[1319:1312];
logic [7:0] input_fmap_165;
assign input_fmap_165 = input_act_ff[1327:1320];
logic [7:0] input_fmap_166;
assign input_fmap_166 = input_act_ff[1335:1328];
logic [7:0] input_fmap_167;
assign input_fmap_167 = input_act_ff[1343:1336];
logic [7:0] input_fmap_168;
assign input_fmap_168 = input_act_ff[1351:1344];
logic [7:0] input_fmap_169;
assign input_fmap_169 = input_act_ff[1359:1352];
logic [7:0] input_fmap_170;
assign input_fmap_170 = input_act_ff[1367:1360];
logic [7:0] input_fmap_171;
assign input_fmap_171 = input_act_ff[1375:1368];
logic [7:0] input_fmap_172;
assign input_fmap_172 = input_act_ff[1383:1376];
logic [7:0] input_fmap_173;
assign input_fmap_173 = input_act_ff[1391:1384];
logic [7:0] input_fmap_174;
assign input_fmap_174 = input_act_ff[1399:1392];
logic [7:0] input_fmap_175;
assign input_fmap_175 = input_act_ff[1407:1400];
logic [7:0] input_fmap_176;
assign input_fmap_176 = input_act_ff[1415:1408];
logic [7:0] input_fmap_177;
assign input_fmap_177 = input_act_ff[1423:1416];
logic [7:0] input_fmap_178;
assign input_fmap_178 = input_act_ff[1431:1424];
logic [7:0] input_fmap_179;
assign input_fmap_179 = input_act_ff[1439:1432];
logic [7:0] input_fmap_180;
assign input_fmap_180 = input_act_ff[1447:1440];
logic [7:0] input_fmap_181;
assign input_fmap_181 = input_act_ff[1455:1448];
logic [7:0] input_fmap_182;
assign input_fmap_182 = input_act_ff[1463:1456];
logic [7:0] input_fmap_183;
assign input_fmap_183 = input_act_ff[1471:1464];
logic [7:0] input_fmap_184;
assign input_fmap_184 = input_act_ff[1479:1472];
logic [7:0] input_fmap_185;
assign input_fmap_185 = input_act_ff[1487:1480];
logic [7:0] input_fmap_186;
assign input_fmap_186 = input_act_ff[1495:1488];
logic [7:0] input_fmap_187;
assign input_fmap_187 = input_act_ff[1503:1496];
logic [7:0] input_fmap_188;
assign input_fmap_188 = input_act_ff[1511:1504];
logic [7:0] input_fmap_189;
assign input_fmap_189 = input_act_ff[1519:1512];
logic [7:0] input_fmap_190;
assign input_fmap_190 = input_act_ff[1527:1520];
logic [7:0] input_fmap_191;
assign input_fmap_191 = input_act_ff[1535:1528];
logic [7:0] input_fmap_192;
assign input_fmap_192 = input_act_ff[1543:1536];
logic [7:0] input_fmap_193;
assign input_fmap_193 = input_act_ff[1551:1544];
logic [7:0] input_fmap_194;
assign input_fmap_194 = input_act_ff[1559:1552];
logic [7:0] input_fmap_195;
assign input_fmap_195 = input_act_ff[1567:1560];
logic [7:0] input_fmap_196;
assign input_fmap_196 = input_act_ff[1575:1568];
logic [7:0] input_fmap_197;
assign input_fmap_197 = input_act_ff[1583:1576];
logic [7:0] input_fmap_198;
assign input_fmap_198 = input_act_ff[1591:1584];
logic [7:0] input_fmap_199;
assign input_fmap_199 = input_act_ff[1599:1592];
logic [7:0] input_fmap_200;
assign input_fmap_200 = input_act_ff[1607:1600];
logic [7:0] input_fmap_201;
assign input_fmap_201 = input_act_ff[1615:1608];
logic [7:0] input_fmap_202;
assign input_fmap_202 = input_act_ff[1623:1616];
logic [7:0] input_fmap_203;
assign input_fmap_203 = input_act_ff[1631:1624];
logic [7:0] input_fmap_204;
assign input_fmap_204 = input_act_ff[1639:1632];
logic [7:0] input_fmap_205;
assign input_fmap_205 = input_act_ff[1647:1640];
logic [7:0] input_fmap_206;
assign input_fmap_206 = input_act_ff[1655:1648];
logic [7:0] input_fmap_207;
assign input_fmap_207 = input_act_ff[1663:1656];
logic [7:0] input_fmap_208;
assign input_fmap_208 = input_act_ff[1671:1664];
logic [7:0] input_fmap_209;
assign input_fmap_209 = input_act_ff[1679:1672];
logic [7:0] input_fmap_210;
assign input_fmap_210 = input_act_ff[1687:1680];
logic [7:0] input_fmap_211;
assign input_fmap_211 = input_act_ff[1695:1688];
logic [7:0] input_fmap_212;
assign input_fmap_212 = input_act_ff[1703:1696];
logic [7:0] input_fmap_213;
assign input_fmap_213 = input_act_ff[1711:1704];
logic [7:0] input_fmap_214;
assign input_fmap_214 = input_act_ff[1719:1712];
logic [7:0] input_fmap_215;
assign input_fmap_215 = input_act_ff[1727:1720];
logic [7:0] input_fmap_216;
assign input_fmap_216 = input_act_ff[1735:1728];
logic [7:0] input_fmap_217;
assign input_fmap_217 = input_act_ff[1743:1736];
logic [7:0] input_fmap_218;
assign input_fmap_218 = input_act_ff[1751:1744];
logic [7:0] input_fmap_219;
assign input_fmap_219 = input_act_ff[1759:1752];
logic [7:0] input_fmap_220;
assign input_fmap_220 = input_act_ff[1767:1760];
logic [7:0] input_fmap_221;
assign input_fmap_221 = input_act_ff[1775:1768];
logic [7:0] input_fmap_222;
assign input_fmap_222 = input_act_ff[1783:1776];
logic [7:0] input_fmap_223;
assign input_fmap_223 = input_act_ff[1791:1784];
logic [7:0] input_fmap_224;
assign input_fmap_224 = input_act_ff[1799:1792];
logic [7:0] input_fmap_225;
assign input_fmap_225 = input_act_ff[1807:1800];
logic [7:0] input_fmap_226;
assign input_fmap_226 = input_act_ff[1815:1808];
logic [7:0] input_fmap_227;
assign input_fmap_227 = input_act_ff[1823:1816];
logic [7:0] input_fmap_228;
assign input_fmap_228 = input_act_ff[1831:1824];
logic [7:0] input_fmap_229;
assign input_fmap_229 = input_act_ff[1839:1832];
logic [7:0] input_fmap_230;
assign input_fmap_230 = input_act_ff[1847:1840];
logic [7:0] input_fmap_231;
assign input_fmap_231 = input_act_ff[1855:1848];
logic [7:0] input_fmap_232;
assign input_fmap_232 = input_act_ff[1863:1856];
logic [7:0] input_fmap_233;
assign input_fmap_233 = input_act_ff[1871:1864];
logic [7:0] input_fmap_234;
assign input_fmap_234 = input_act_ff[1879:1872];
logic [7:0] input_fmap_235;
assign input_fmap_235 = input_act_ff[1887:1880];
logic [7:0] input_fmap_236;
assign input_fmap_236 = input_act_ff[1895:1888];
logic [7:0] input_fmap_237;
assign input_fmap_237 = input_act_ff[1903:1896];
logic [7:0] input_fmap_238;
assign input_fmap_238 = input_act_ff[1911:1904];
logic [7:0] input_fmap_239;
assign input_fmap_239 = input_act_ff[1919:1912];
logic [7:0] input_fmap_240;
assign input_fmap_240 = input_act_ff[1927:1920];
logic [7:0] input_fmap_241;
assign input_fmap_241 = input_act_ff[1935:1928];
logic [7:0] input_fmap_242;
assign input_fmap_242 = input_act_ff[1943:1936];
logic [7:0] input_fmap_243;
assign input_fmap_243 = input_act_ff[1951:1944];
logic [7:0] input_fmap_244;
assign input_fmap_244 = input_act_ff[1959:1952];
logic [7:0] input_fmap_245;
assign input_fmap_245 = input_act_ff[1967:1960];
logic [7:0] input_fmap_246;
assign input_fmap_246 = input_act_ff[1975:1968];
logic [7:0] input_fmap_247;
assign input_fmap_247 = input_act_ff[1983:1976];
logic [7:0] input_fmap_248;
assign input_fmap_248 = input_act_ff[1991:1984];
logic [7:0] input_fmap_249;
assign input_fmap_249 = input_act_ff[1999:1992];
logic [7:0] input_fmap_250;
assign input_fmap_250 = input_act_ff[2007:2000];
logic [7:0] input_fmap_251;
assign input_fmap_251 = input_act_ff[2015:2008];
logic [7:0] input_fmap_252;
assign input_fmap_252 = input_act_ff[2023:2016];
logic [7:0] input_fmap_253;
assign input_fmap_253 = input_act_ff[2031:2024];
logic [7:0] input_fmap_254;
assign input_fmap_254 = input_act_ff[2039:2032];
logic [7:0] input_fmap_255;
assign input_fmap_255 = input_act_ff[2047:2040];

logic signed [31:0] conv_mac_0;
assign conv_mac_0 = 
	( 16'sd 31557) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8517) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26429) * $signed(input_fmap_3[7:0]) +
	( 11'sd 715) * $signed(input_fmap_4[7:0]) +
	( 10'sd 256) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8859) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29406) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24281) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19617) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11755) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30342) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5280) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1986) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6021) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13956) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19329) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31072) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28573) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7118) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12079) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25277) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16099) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7488) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15705) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17862) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3243) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31720) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29271) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16236) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_32[7:0]) +
	( 11'sd 771) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2201) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20659) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12630) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20161) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30218) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27808) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6964) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5685) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7876) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16722) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21942) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9883) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21121) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21202) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1840) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17219) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27743) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26289) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_54[7:0]) +
	( 13'sd 4017) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15256) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10133) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31111) * $signed(input_fmap_59[7:0]) +
	( 11'sd 609) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12420) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12619) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24469) * $signed(input_fmap_63[7:0]) +
	( 10'sd 441) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27907) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29962) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24501) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9944) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29415) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28273) * $signed(input_fmap_74[7:0]) +
	( 11'sd 986) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18952) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10412) * $signed(input_fmap_79[7:0]) +
	( 11'sd 969) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21652) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30773) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7358) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13785) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15478) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16177) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4517) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2049) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1039) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3757) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6555) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12167) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18157) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20927) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28110) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1694) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12645) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17673) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23171) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5602) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19639) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20345) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17407) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1640) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20652) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4774) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18218) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_110[7:0]) +
	( 9'sd 130) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3091) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15130) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8052) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20268) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8312) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23859) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4273) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4570) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23726) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8708) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25948) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17148) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12537) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29633) * $signed(input_fmap_128[7:0]) +
	( 14'sd 4204) * $signed(input_fmap_129[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_130[7:0]) +
	( 14'sd 8105) * $signed(input_fmap_131[7:0]) +
	( 16'sd 31081) * $signed(input_fmap_132[7:0]) +
	( 15'sd 14663) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11730) * $signed(input_fmap_134[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23467) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12784) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18759) * $signed(input_fmap_139[7:0]) +
	( 16'sd 19334) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10892) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14622) * $signed(input_fmap_142[7:0]) +
	( 13'sd 3679) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6690) * $signed(input_fmap_144[7:0]) +
	( 14'sd 4738) * $signed(input_fmap_145[7:0]) +
	( 15'sd 8949) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18481) * $signed(input_fmap_147[7:0]) +
	( 16'sd 24532) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23167) * $signed(input_fmap_149[7:0]) +
	( 14'sd 4101) * $signed(input_fmap_150[7:0]) +
	( 16'sd 26301) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16737) * $signed(input_fmap_152[7:0]) +
	( 15'sd 13062) * $signed(input_fmap_153[7:0]) +
	( 15'sd 13653) * $signed(input_fmap_154[7:0]) +
	( 16'sd 18266) * $signed(input_fmap_155[7:0]) +
	( 12'sd 1286) * $signed(input_fmap_156[7:0]) +
	( 15'sd 8639) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18476) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27411) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21190) * $signed(input_fmap_160[7:0]) +
	( 15'sd 10444) * $signed(input_fmap_161[7:0]) +
	( 16'sd 19100) * $signed(input_fmap_162[7:0]) +
	( 10'sd 380) * $signed(input_fmap_163[7:0]) +
	( 16'sd 17739) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22282) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9974) * $signed(input_fmap_166[7:0]) +
	( 15'sd 11535) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6829) * $signed(input_fmap_168[7:0]) +
	( 12'sd 1408) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14400) * $signed(input_fmap_170[7:0]) +
	( 15'sd 13149) * $signed(input_fmap_171[7:0]) +
	( 15'sd 13560) * $signed(input_fmap_172[7:0]) +
	( 16'sd 20983) * $signed(input_fmap_173[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_174[7:0]) +
	( 16'sd 24023) * $signed(input_fmap_175[7:0]) +
	( 16'sd 28190) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24997) * $signed(input_fmap_177[7:0]) +
	( 15'sd 12336) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5794) * $signed(input_fmap_179[7:0]) +
	( 15'sd 8949) * $signed(input_fmap_180[7:0]) +
	( 4'sd 6) * $signed(input_fmap_181[7:0]) +
	( 15'sd 14622) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12076) * $signed(input_fmap_183[7:0]) +
	( 16'sd 20496) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17113) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12177) * $signed(input_fmap_186[7:0]) +
	( 16'sd 26718) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2375) * $signed(input_fmap_188[7:0]) +
	( 16'sd 27626) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13585) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17836) * $signed(input_fmap_191[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_192[7:0]) +
	( 14'sd 4236) * $signed(input_fmap_193[7:0]) +
	( 16'sd 19059) * $signed(input_fmap_194[7:0]) +
	( 11'sd 874) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31114) * $signed(input_fmap_197[7:0]) +
	( 15'sd 8886) * $signed(input_fmap_198[7:0]) +
	( 15'sd 11968) * $signed(input_fmap_199[7:0]) +
	( 16'sd 23664) * $signed(input_fmap_200[7:0]) +
	( 15'sd 14862) * $signed(input_fmap_201[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19502) * $signed(input_fmap_204[7:0]) +
	( 16'sd 20503) * $signed(input_fmap_205[7:0]) +
	( 14'sd 4743) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28361) * $signed(input_fmap_207[7:0]) +
	( 14'sd 8062) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23599) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4357) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12062) * $signed(input_fmap_211[7:0]) +
	( 16'sd 23474) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2423) * $signed(input_fmap_213[7:0]) +
	( 14'sd 6029) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7572) * $signed(input_fmap_215[7:0]) +
	( 15'sd 10661) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10331) * $signed(input_fmap_217[7:0]) +
	( 15'sd 9297) * $signed(input_fmap_218[7:0]) +
	( 16'sd 30975) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30670) * $signed(input_fmap_220[7:0]) +
	( 16'sd 20994) * $signed(input_fmap_221[7:0]) +
	( 16'sd 20791) * $signed(input_fmap_222[7:0]) +
	( 12'sd 1369) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27564) * $signed(input_fmap_224[7:0]) +
	( 16'sd 23500) * $signed(input_fmap_225[7:0]) +
	( 15'sd 8513) * $signed(input_fmap_226[7:0]) +
	( 16'sd 30861) * $signed(input_fmap_227[7:0]) +
	( 16'sd 23467) * $signed(input_fmap_228[7:0]) +
	( 14'sd 4795) * $signed(input_fmap_229[7:0]) +
	( 15'sd 10978) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25539) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8657) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_233[7:0]) +
	( 16'sd 32206) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3425) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2915) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28296) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3953) * $signed(input_fmap_238[7:0]) +
	( 15'sd 16186) * $signed(input_fmap_239[7:0]) +
	( 16'sd 16700) * $signed(input_fmap_240[7:0]) +
	( 15'sd 12911) * $signed(input_fmap_241[7:0]) +
	( 15'sd 9817) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7025) * $signed(input_fmap_243[7:0]) +
	( 13'sd 3246) * $signed(input_fmap_244[7:0]) +
	( 16'sd 29966) * $signed(input_fmap_245[7:0]) +
	( 16'sd 26715) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17096) * $signed(input_fmap_247[7:0]) +
	( 16'sd 30000) * $signed(input_fmap_248[7:0]) +
	( 16'sd 22878) * $signed(input_fmap_249[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_250[7:0]) +
	( 16'sd 29642) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10926) * $signed(input_fmap_252[7:0]) +
	( 16'sd 23811) * $signed(input_fmap_253[7:0]) +
	( 15'sd 15453) * $signed(input_fmap_254[7:0]) +
	( 16'sd 25796) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_1;
assign conv_mac_1 = 
	( 13'sd 3941) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7972) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27228) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10091) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2153) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14417) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8945) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3839) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2788) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28625) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7952) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3298) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30186) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17530) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28572) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4505) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4804) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20405) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25134) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5345) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18701) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9039) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31581) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18517) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5469) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3644) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14845) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24293) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28880) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3255) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30003) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24878) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21494) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19050) * $signed(input_fmap_37[7:0]) +
	( 10'sd 441) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30243) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8699) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30912) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9480) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22724) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28529) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29861) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10507) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15872) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22847) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23465) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19438) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5573) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32150) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18733) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10699) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12791) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1040) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1315) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20745) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1970) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25512) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29017) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29774) * $signed(input_fmap_64[7:0]) +
	( 14'sd 8148) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21612) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19460) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25396) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19469) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30490) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28430) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23458) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22117) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2073) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31840) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10264) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2589) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26873) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3255) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11010) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11918) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23790) * $signed(input_fmap_83[7:0]) +
	( 11'sd 919) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25998) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29339) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32572) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24842) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29063) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25663) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22279) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10872) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27608) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13576) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26095) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6612) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31657) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12084) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15606) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27245) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5539) * $signed(input_fmap_104[7:0]) +
	( 9'sd 149) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6700) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13943) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28013) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4265) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30028) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7636) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14375) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6630) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19953) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14034) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20162) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26630) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17535) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17041) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10420) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31131) * $signed(input_fmap_123[7:0]) +
	( 7'sd 62) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4412) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30684) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4898) * $signed(input_fmap_128[7:0]) +
	( 15'sd 16222) * $signed(input_fmap_129[7:0]) +
	( 16'sd 32073) * $signed(input_fmap_130[7:0]) +
	( 15'sd 10043) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11531) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31492) * $signed(input_fmap_133[7:0]) +
	( 14'sd 7943) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19536) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31216) * $signed(input_fmap_136[7:0]) +
	( 15'sd 14659) * $signed(input_fmap_137[7:0]) +
	( 16'sd 25118) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20636) * $signed(input_fmap_139[7:0]) +
	( 14'sd 7490) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13265) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31146) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31953) * $signed(input_fmap_143[7:0]) +
	( 11'sd 715) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_145[7:0]) +
	( 16'sd 25838) * $signed(input_fmap_146[7:0]) +
	( 14'sd 7448) * $signed(input_fmap_147[7:0]) +
	( 16'sd 25003) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15100) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18554) * $signed(input_fmap_150[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_151[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_152[7:0]) +
	( 14'sd 5194) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31024) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_155[7:0]) +
	( 13'sd 3376) * $signed(input_fmap_156[7:0]) +
	( 16'sd 28222) * $signed(input_fmap_157[7:0]) +
	( 16'sd 27106) * $signed(input_fmap_158[7:0]) +
	( 16'sd 29107) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18527) * $signed(input_fmap_160[7:0]) +
	( 15'sd 11042) * $signed(input_fmap_161[7:0]) +
	( 15'sd 12012) * $signed(input_fmap_162[7:0]) +
	( 16'sd 19711) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24696) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9192) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_166[7:0]) +
	( 15'sd 11863) * $signed(input_fmap_167[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_168[7:0]) +
	( 14'sd 7103) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17101) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15168) * $signed(input_fmap_171[7:0]) +
	( 15'sd 13683) * $signed(input_fmap_172[7:0]) +
	( 15'sd 14548) * $signed(input_fmap_173[7:0]) +
	( 16'sd 24589) * $signed(input_fmap_174[7:0]) +
	( 15'sd 16131) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20985) * $signed(input_fmap_176[7:0]) +
	( 16'sd 20171) * $signed(input_fmap_177[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3608) * $signed(input_fmap_179[7:0]) +
	( 13'sd 2923) * $signed(input_fmap_180[7:0]) +
	( 16'sd 21934) * $signed(input_fmap_181[7:0]) +
	( 15'sd 14707) * $signed(input_fmap_182[7:0]) +
	( 13'sd 3687) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11513) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1339) * $signed(input_fmap_185[7:0]) +
	( 16'sd 21813) * $signed(input_fmap_186[7:0]) +
	( 16'sd 32107) * $signed(input_fmap_187[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2265) * $signed(input_fmap_189[7:0]) +
	( 16'sd 23051) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29953) * $signed(input_fmap_191[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6443) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14721) * $signed(input_fmap_194[7:0]) +
	( 15'sd 15927) * $signed(input_fmap_195[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21811) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9336) * $signed(input_fmap_198[7:0]) +
	( 16'sd 21417) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6788) * $signed(input_fmap_200[7:0]) +
	( 16'sd 26293) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8566) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21258) * $signed(input_fmap_203[7:0]) +
	( 14'sd 7138) * $signed(input_fmap_204[7:0]) +
	( 16'sd 16995) * $signed(input_fmap_205[7:0]) +
	( 11'sd 612) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3181) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18321) * $signed(input_fmap_208[7:0]) +
	( 15'sd 12735) * $signed(input_fmap_209[7:0]) +
	( 16'sd 16865) * $signed(input_fmap_210[7:0]) +
	( 12'sd 1334) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18091) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29935) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15548) * $signed(input_fmap_214[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_215[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_216[7:0]) +
	( 14'sd 7125) * $signed(input_fmap_217[7:0]) +
	( 12'sd 2016) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31369) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15580) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12408) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19464) * $signed(input_fmap_223[7:0]) +
	( 16'sd 23604) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14611) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_226[7:0]) +
	( 11'sd 610) * $signed(input_fmap_227[7:0]) +
	( 15'sd 9807) * $signed(input_fmap_228[7:0]) +
	( 9'sd 169) * $signed(input_fmap_229[7:0]) +
	( 15'sd 9298) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24405) * $signed(input_fmap_231[7:0]) +
	( 14'sd 5527) * $signed(input_fmap_232[7:0]) +
	( 16'sd 26373) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3157) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29306) * $signed(input_fmap_235[7:0]) +
	( 12'sd 1457) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14687) * $signed(input_fmap_237[7:0]) +
	( 16'sd 18152) * $signed(input_fmap_238[7:0]) +
	( 16'sd 30316) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9735) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7787) * $signed(input_fmap_241[7:0]) +
	( 15'sd 9641) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23514) * $signed(input_fmap_243[7:0]) +
	( 16'sd 21091) * $signed(input_fmap_244[7:0]) +
	( 15'sd 8231) * $signed(input_fmap_245[7:0]) +
	( 15'sd 8325) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_247[7:0]) +
	( 16'sd 31080) * $signed(input_fmap_248[7:0]) +
	( 15'sd 8984) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26879) * $signed(input_fmap_250[7:0]) +
	( 12'sd 1099) * $signed(input_fmap_251[7:0]) +
	( 15'sd 14725) * $signed(input_fmap_252[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13064) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14100) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_2;
assign conv_mac_2 = 
	( 16'sd 32352) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6759) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23315) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26462) * $signed(input_fmap_3[7:0]) +
	( 10'sd 378) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20673) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30824) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1881) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13938) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6987) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32433) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15157) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30732) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10690) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17975) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4348) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6871) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17199) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7382) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29273) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14321) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5199) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18181) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3822) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7085) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1963) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27791) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30027) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5133) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13135) * $signed(input_fmap_31[7:0]) +
	( 4'sd 6) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20212) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17020) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29338) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7539) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28686) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22606) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23544) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26410) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31564) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13024) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11564) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2144) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9617) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9718) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10687) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6743) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27760) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6442) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32195) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1820) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12397) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23625) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6088) * $signed(input_fmap_58[7:0]) +
	( 11'sd 626) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14321) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31927) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20689) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7528) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31174) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4380) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2422) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10145) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18455) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18748) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10867) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32185) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15167) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18139) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3825) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20096) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1601) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26974) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24572) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11356) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21326) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27356) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23962) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27721) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11955) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19429) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7940) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18371) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25634) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32373) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30951) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8630) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30493) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10914) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22627) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15108) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4440) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16908) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28789) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2612) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21035) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13115) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19093) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30670) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17049) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13609) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13952) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22361) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32525) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28300) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4634) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27457) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23735) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16965) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7402) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19235) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26228) * $signed(input_fmap_125[7:0]) +
	( 11'sd 924) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18378) * $signed(input_fmap_127[7:0]) +
	( 14'sd 5880) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10318) * $signed(input_fmap_129[7:0]) +
	( 16'sd 21211) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_131[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_132[7:0]) +
	( 16'sd 20280) * $signed(input_fmap_133[7:0]) +
	( 11'sd 687) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10743) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15034) * $signed(input_fmap_136[7:0]) +
	( 16'sd 17378) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21744) * $signed(input_fmap_139[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_140[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28425) * $signed(input_fmap_142[7:0]) +
	( 16'sd 25646) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4554) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25353) * $signed(input_fmap_145[7:0]) +
	( 14'sd 4815) * $signed(input_fmap_146[7:0]) +
	( 15'sd 10546) * $signed(input_fmap_147[7:0]) +
	( 16'sd 30842) * $signed(input_fmap_148[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_149[7:0]) +
	( 13'sd 2516) * $signed(input_fmap_150[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27142) * $signed(input_fmap_153[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27380) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7116) * $signed(input_fmap_156[7:0]) +
	( 16'sd 21769) * $signed(input_fmap_157[7:0]) +
	( 16'sd 31727) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21031) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6035) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22400) * $signed(input_fmap_161[7:0]) +
	( 16'sd 19129) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2510) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11003) * $signed(input_fmap_164[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_165[7:0]) +
	( 15'sd 11167) * $signed(input_fmap_166[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6832) * $signed(input_fmap_168[7:0]) +
	( 15'sd 15684) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24402) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20397) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3346) * $signed(input_fmap_172[7:0]) +
	( 16'sd 30103) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11682) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4513) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7880) * $signed(input_fmap_176[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15794) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18817) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27463) * $signed(input_fmap_180[7:0]) +
	( 13'sd 2988) * $signed(input_fmap_181[7:0]) +
	( 11'sd 890) * $signed(input_fmap_182[7:0]) +
	( 15'sd 11527) * $signed(input_fmap_183[7:0]) +
	( 13'sd 2097) * $signed(input_fmap_184[7:0]) +
	( 15'sd 13021) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13713) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_188[7:0]) +
	( 8'sd 102) * $signed(input_fmap_189[7:0]) +
	( 16'sd 32101) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23250) * $signed(input_fmap_191[7:0]) +
	( 16'sd 23817) * $signed(input_fmap_192[7:0]) +
	( 16'sd 24224) * $signed(input_fmap_193[7:0]) +
	( 16'sd 20026) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17363) * $signed(input_fmap_195[7:0]) +
	( 16'sd 27442) * $signed(input_fmap_196[7:0]) +
	( 14'sd 7813) * $signed(input_fmap_197[7:0]) +
	( 11'sd 883) * $signed(input_fmap_198[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_199[7:0]) +
	( 15'sd 12452) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21627) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21098) * $signed(input_fmap_202[7:0]) +
	( 16'sd 26123) * $signed(input_fmap_203[7:0]) +
	( 16'sd 18029) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24403) * $signed(input_fmap_205[7:0]) +
	( 16'sd 25862) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12763) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15165) * $signed(input_fmap_208[7:0]) +
	( 15'sd 12359) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19183) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20401) * $signed(input_fmap_211[7:0]) +
	( 16'sd 16733) * $signed(input_fmap_212[7:0]) +
	( 15'sd 15422) * $signed(input_fmap_213[7:0]) +
	( 16'sd 29954) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7065) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_216[7:0]) +
	( 12'sd 1465) * $signed(input_fmap_217[7:0]) +
	( 15'sd 11389) * $signed(input_fmap_218[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_219[7:0]) +
	( 16'sd 16800) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27998) * $signed(input_fmap_221[7:0]) +
	( 16'sd 16575) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17332) * $signed(input_fmap_223[7:0]) +
	( 16'sd 26637) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7789) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2839) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19805) * $signed(input_fmap_228[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18069) * $signed(input_fmap_230[7:0]) +
	( 15'sd 12669) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15702) * $signed(input_fmap_232[7:0]) +
	( 14'sd 7708) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19176) * $signed(input_fmap_234[7:0]) +
	( 14'sd 4914) * $signed(input_fmap_235[7:0]) +
	( 15'sd 13383) * $signed(input_fmap_236[7:0]) +
	( 11'sd 1007) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19443) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31039) * $signed(input_fmap_239[7:0]) +
	( 15'sd 11657) * $signed(input_fmap_240[7:0]) +
	( 15'sd 16280) * $signed(input_fmap_241[7:0]) +
	( 14'sd 8166) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_243[7:0]) +
	( 15'sd 11159) * $signed(input_fmap_244[7:0]) +
	( 16'sd 16506) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23021) * $signed(input_fmap_246[7:0]) +
	( 14'sd 8131) * $signed(input_fmap_247[7:0]) +
	( 16'sd 29616) * $signed(input_fmap_248[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_250[7:0]) +
	( 16'sd 24798) * $signed(input_fmap_251[7:0]) +
	( 15'sd 8904) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3274) * $signed(input_fmap_253[7:0]) +
	( 14'sd 7121) * $signed(input_fmap_254[7:0]) +
	( 10'sd 432) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_3;
assign conv_mac_3 = 
	( 13'sd 2760) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31473) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24081) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28569) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22580) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5264) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6626) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11752) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24660) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18880) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20529) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28645) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25819) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12335) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18842) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5230) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32025) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17137) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31178) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5500) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23732) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8656) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10352) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21406) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9161) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3202) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30985) * $signed(input_fmap_32[7:0]) +
	( 11'sd 694) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30013) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24308) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12290) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6326) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3472) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15937) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25040) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7004) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5064) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4408) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20892) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2608) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28808) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17338) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22109) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25286) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7439) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32758) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25524) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17237) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6232) * $signed(input_fmap_57[7:0]) +
	( 11'sd 639) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24197) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3391) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3392) * $signed(input_fmap_61[7:0]) +
	( 11'sd 538) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9473) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27119) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23079) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31938) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15277) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6687) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4997) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20139) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2828) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24848) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13949) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22211) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24470) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7010) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10125) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19980) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_80[7:0]) +
	( 13'sd 4031) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18532) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10555) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7137) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21431) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12768) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24110) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11768) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8983) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12049) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14717) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24719) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20069) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9637) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8727) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14825) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31807) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6128) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6423) * $signed(input_fmap_101[7:0]) +
	( 11'sd 758) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1924) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13338) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25588) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9156) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9430) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13677) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24780) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19552) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30031) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27521) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12328) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25512) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18583) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1540) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19525) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7272) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24958) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16174) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18988) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13716) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25116) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19288) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15495) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9581) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7471) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_130[7:0]) +
	( 14'sd 6011) * $signed(input_fmap_131[7:0]) +
	( 10'sd 306) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21820) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28331) * $signed(input_fmap_135[7:0]) +
	( 15'sd 10221) * $signed(input_fmap_136[7:0]) +
	( 15'sd 10139) * $signed(input_fmap_137[7:0]) +
	( 15'sd 14165) * $signed(input_fmap_138[7:0]) +
	( 16'sd 22714) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17573) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29263) * $signed(input_fmap_141[7:0]) +
	( 15'sd 15884) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9055) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26461) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18004) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17757) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21324) * $signed(input_fmap_148[7:0]) +
	( 16'sd 19988) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21015) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12335) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31188) * $signed(input_fmap_152[7:0]) +
	( 16'sd 32435) * $signed(input_fmap_153[7:0]) +
	( 15'sd 9064) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22279) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13249) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_158[7:0]) +
	( 16'sd 16481) * $signed(input_fmap_159[7:0]) +
	( 12'sd 1642) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4908) * $signed(input_fmap_161[7:0]) +
	( 11'sd 826) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20416) * $signed(input_fmap_163[7:0]) +
	( 16'sd 26126) * $signed(input_fmap_164[7:0]) +
	( 16'sd 25804) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22694) * $signed(input_fmap_166[7:0]) +
	( 12'sd 1622) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6360) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10259) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20693) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31247) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22384) * $signed(input_fmap_172[7:0]) +
	( 14'sd 7284) * $signed(input_fmap_173[7:0]) +
	( 15'sd 9658) * $signed(input_fmap_174[7:0]) +
	( 16'sd 22369) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29160) * $signed(input_fmap_176[7:0]) +
	( 16'sd 28969) * $signed(input_fmap_177[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25280) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29009) * $signed(input_fmap_180[7:0]) +
	( 12'sd 1747) * $signed(input_fmap_181[7:0]) +
	( 16'sd 22784) * $signed(input_fmap_182[7:0]) +
	( 16'sd 21885) * $signed(input_fmap_183[7:0]) +
	( 16'sd 20525) * $signed(input_fmap_184[7:0]) +
	( 16'sd 32269) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23101) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12154) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19529) * $signed(input_fmap_189[7:0]) +
	( 15'sd 14148) * $signed(input_fmap_190[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31633) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27934) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29711) * $signed(input_fmap_194[7:0]) +
	( 14'sd 4155) * $signed(input_fmap_195[7:0]) +
	( 13'sd 4066) * $signed(input_fmap_196[7:0]) +
	( 15'sd 9254) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18178) * $signed(input_fmap_198[7:0]) +
	( 16'sd 17720) * $signed(input_fmap_199[7:0]) +
	( 15'sd 12392) * $signed(input_fmap_200[7:0]) +
	( 15'sd 14056) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17654) * $signed(input_fmap_202[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5356) * $signed(input_fmap_204[7:0]) +
	( 16'sd 26956) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31959) * $signed(input_fmap_206[7:0]) +
	( 16'sd 22970) * $signed(input_fmap_207[7:0]) +
	( 16'sd 29783) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22933) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31680) * $signed(input_fmap_210[7:0]) +
	( 14'sd 4423) * $signed(input_fmap_211[7:0]) +
	( 15'sd 13960) * $signed(input_fmap_212[7:0]) +
	( 16'sd 16404) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7602) * $signed(input_fmap_214[7:0]) +
	( 16'sd 20860) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1573) * $signed(input_fmap_216[7:0]) +
	( 16'sd 27169) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26172) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20197) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21933) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27066) * $signed(input_fmap_221[7:0]) +
	( 16'sd 23298) * $signed(input_fmap_222[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_223[7:0]) +
	( 14'sd 5438) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26328) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22039) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3340) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22938) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_229[7:0]) +
	( 16'sd 23902) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25811) * $signed(input_fmap_231[7:0]) +
	( 11'sd 763) * $signed(input_fmap_232[7:0]) +
	( 16'sd 31975) * $signed(input_fmap_233[7:0]) +
	( 10'sd 397) * $signed(input_fmap_234[7:0]) +
	( 16'sd 20602) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_236[7:0]) +
	( 16'sd 21540) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14328) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19707) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19829) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29727) * $signed(input_fmap_241[7:0]) +
	( 14'sd 8118) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2350) * $signed(input_fmap_243[7:0]) +
	( 14'sd 5692) * $signed(input_fmap_244[7:0]) +
	( 16'sd 31612) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30330) * $signed(input_fmap_246[7:0]) +
	( 15'sd 10940) * $signed(input_fmap_247[7:0]) +
	( 15'sd 15599) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28660) * $signed(input_fmap_249[7:0]) +
	( 15'sd 14879) * $signed(input_fmap_250[7:0]) +
	( 16'sd 29681) * $signed(input_fmap_251[7:0]) +
	( 16'sd 32762) * $signed(input_fmap_252[7:0]) +
	( 16'sd 18324) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13722) * $signed(input_fmap_254[7:0]) +
	( 16'sd 17687) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_4;
assign conv_mac_4 = 
	( 15'sd 12527) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28526) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19250) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12476) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17449) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15706) * $signed(input_fmap_5[7:0]) +
	( 11'sd 793) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10654) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32166) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21646) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7362) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24326) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4182) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12718) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32060) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12681) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27162) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17540) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20936) * $signed(input_fmap_18[7:0]) +
	( 11'sd 701) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26212) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19202) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3661) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20444) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16433) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26573) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21280) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32690) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13166) * $signed(input_fmap_31[7:0]) +
	( 10'sd 490) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23177) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20060) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17422) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9448) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27429) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3136) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3882) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2439) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3052) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9213) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13537) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29779) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2886) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25253) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10828) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25062) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7188) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7149) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5102) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20671) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32021) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11120) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13771) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18064) * $signed(input_fmap_58[7:0]) +
	( 10'sd 401) * $signed(input_fmap_59[7:0]) +
	( 11'sd 876) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20750) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31866) * $signed(input_fmap_62[7:0]) +
	( 9'sd 205) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16147) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25400) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25026) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10025) * $signed(input_fmap_68[7:0]) +
	( 11'sd 970) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25459) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1887) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20997) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21634) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23391) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2188) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4625) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10495) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20199) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7771) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18286) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28010) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7550) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22080) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25721) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30820) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26496) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19929) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3131) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22786) * $signed(input_fmap_93[7:0]) +
	( 9'sd 135) * $signed(input_fmap_94[7:0]) +
	( 11'sd 744) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31048) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8523) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24003) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6761) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29190) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6327) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30660) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21649) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6051) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2575) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31835) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5985) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19472) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13133) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16708) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7009) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30162) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23393) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21593) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11092) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22543) * $signed(input_fmap_118[7:0]) +
	( 10'sd 330) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4108) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32211) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19984) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17650) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30013) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9598) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30304) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25825) * $signed(input_fmap_127[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19958) * $signed(input_fmap_129[7:0]) +
	( 15'sd 16160) * $signed(input_fmap_130[7:0]) +
	( 16'sd 30325) * $signed(input_fmap_131[7:0]) +
	( 14'sd 6693) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12081) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_134[7:0]) +
	( 15'sd 9036) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23352) * $signed(input_fmap_136[7:0]) +
	( 14'sd 7970) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31820) * $signed(input_fmap_138[7:0]) +
	( 16'sd 16883) * $signed(input_fmap_139[7:0]) +
	( 16'sd 25268) * $signed(input_fmap_140[7:0]) +
	( 14'sd 4341) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6528) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_143[7:0]) +
	( 14'sd 7325) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27737) * $signed(input_fmap_145[7:0]) +
	( 16'sd 30591) * $signed(input_fmap_146[7:0]) +
	( 16'sd 25486) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_148[7:0]) +
	( 16'sd 31390) * $signed(input_fmap_149[7:0]) +
	( 16'sd 30840) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30143) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7945) * $signed(input_fmap_152[7:0]) +
	( 16'sd 26073) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25240) * $signed(input_fmap_154[7:0]) +
	( 15'sd 8748) * $signed(input_fmap_155[7:0]) +
	( 11'sd 529) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_157[7:0]) +
	( 13'sd 2291) * $signed(input_fmap_158[7:0]) +
	( 15'sd 10309) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22583) * $signed(input_fmap_160[7:0]) +
	( 15'sd 14832) * $signed(input_fmap_161[7:0]) +
	( 15'sd 16289) * $signed(input_fmap_162[7:0]) +
	( 16'sd 18316) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8643) * $signed(input_fmap_164[7:0]) +
	( 12'sd 1768) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2406) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31338) * $signed(input_fmap_167[7:0]) +
	( 10'sd 277) * $signed(input_fmap_168[7:0]) +
	( 16'sd 29483) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11639) * $signed(input_fmap_172[7:0]) +
	( 14'sd 4340) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19704) * $signed(input_fmap_174[7:0]) +
	( 16'sd 23882) * $signed(input_fmap_175[7:0]) +
	( 16'sd 23520) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_177[7:0]) +
	( 13'sd 3515) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20091) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23922) * $signed(input_fmap_180[7:0]) +
	( 16'sd 17556) * $signed(input_fmap_181[7:0]) +
	( 15'sd 11135) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12231) * $signed(input_fmap_183[7:0]) +
	( 15'sd 16053) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25011) * $signed(input_fmap_185[7:0]) +
	( 16'sd 32700) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25233) * $signed(input_fmap_187[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3411) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28532) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29412) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31746) * $signed(input_fmap_192[7:0]) +
	( 13'sd 2881) * $signed(input_fmap_193[7:0]) +
	( 16'sd 22635) * $signed(input_fmap_194[7:0]) +
	( 13'sd 4085) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15861) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5631) * $signed(input_fmap_197[7:0]) +
	( 12'sd 1861) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20599) * $signed(input_fmap_199[7:0]) +
	( 16'sd 19578) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3874) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17513) * $signed(input_fmap_202[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_203[7:0]) +
	( 15'sd 13464) * $signed(input_fmap_204[7:0]) +
	( 16'sd 26260) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6220) * $signed(input_fmap_206[7:0]) +
	( 12'sd 2035) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25167) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13093) * $signed(input_fmap_209[7:0]) +
	( 13'sd 2809) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3640) * $signed(input_fmap_211[7:0]) +
	( 13'sd 3285) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9972) * $signed(input_fmap_213[7:0]) +
	( 16'sd 22574) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6178) * $signed(input_fmap_215[7:0]) +
	( 13'sd 2386) * $signed(input_fmap_216[7:0]) +
	( 15'sd 11269) * $signed(input_fmap_217[7:0]) +
	( 16'sd 25712) * $signed(input_fmap_218[7:0]) +
	( 16'sd 32626) * $signed(input_fmap_219[7:0]) +
	( 13'sd 3893) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28679) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19758) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12007) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27823) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14234) * $signed(input_fmap_225[7:0]) +
	( 16'sd 25922) * $signed(input_fmap_226[7:0]) +
	( 16'sd 23491) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22056) * $signed(input_fmap_228[7:0]) +
	( 16'sd 16418) * $signed(input_fmap_229[7:0]) +
	( 12'sd 1538) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31228) * $signed(input_fmap_231[7:0]) +
	( 14'sd 4736) * $signed(input_fmap_232[7:0]) +
	( 16'sd 16904) * $signed(input_fmap_233[7:0]) +
	( 16'sd 26600) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11806) * $signed(input_fmap_235[7:0]) +
	( 14'sd 6517) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29581) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22991) * $signed(input_fmap_238[7:0]) +
	( 16'sd 27109) * $signed(input_fmap_239[7:0]) +
	( 16'sd 29389) * $signed(input_fmap_240[7:0]) +
	( 15'sd 9340) * $signed(input_fmap_241[7:0]) +
	( 16'sd 18753) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28052) * $signed(input_fmap_243[7:0]) +
	( 16'sd 29601) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14845) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30945) * $signed(input_fmap_246[7:0]) +
	( 14'sd 5849) * $signed(input_fmap_247[7:0]) +
	( 16'sd 29291) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21034) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3201) * $signed(input_fmap_250[7:0]) +
	( 16'sd 28297) * $signed(input_fmap_251[7:0]) +
	( 12'sd 1906) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6280) * $signed(input_fmap_253[7:0]) +
	( 15'sd 14691) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5338) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_5;
assign conv_mac_5 = 
	( 16'sd 23652) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12473) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22285) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9426) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32059) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13379) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23680) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24309) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11605) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15710) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15098) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7093) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5424) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21376) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24887) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1323) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21596) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32156) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16838) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22996) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14988) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16993) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6736) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17751) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31609) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15134) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16258) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19342) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24896) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10553) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16199) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3253) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28198) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10724) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12444) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26621) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29735) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17124) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30337) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30612) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20429) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_46[7:0]) +
	( 8'sd 90) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21673) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21164) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16316) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14014) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23227) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30075) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14418) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18404) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16772) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4834) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28812) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2908) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32151) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24097) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4964) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5975) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12335) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8444) * $signed(input_fmap_65[7:0]) +
	( 10'sd 489) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32409) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31116) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17274) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27056) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3317) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22477) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21836) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5852) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1527) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6195) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6242) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16292) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10137) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27836) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30932) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19223) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18793) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15961) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11679) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20546) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18376) * $signed(input_fmap_96[7:0]) +
	( 14'sd 8078) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14534) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9177) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10637) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1684) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4320) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17684) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19255) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21838) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30732) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24366) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10542) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17188) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19147) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27708) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16938) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24781) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5042) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25687) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15318) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30055) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13645) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14929) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5721) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25787) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12687) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21628) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5384) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_128[7:0]) +
	( 16'sd 23389) * $signed(input_fmap_129[7:0]) +
	( 16'sd 28413) * $signed(input_fmap_130[7:0]) +
	( 11'sd 534) * $signed(input_fmap_131[7:0]) +
	( 16'sd 23944) * $signed(input_fmap_132[7:0]) +
	( 16'sd 18127) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11876) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28195) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30424) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13717) * $signed(input_fmap_137[7:0]) +
	( 16'sd 26066) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_139[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12121) * $signed(input_fmap_141[7:0]) +
	( 16'sd 32379) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17932) * $signed(input_fmap_143[7:0]) +
	( 14'sd 7809) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3795) * $signed(input_fmap_147[7:0]) +
	( 16'sd 29788) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18462) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31367) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29361) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27088) * $signed(input_fmap_153[7:0]) +
	( 12'sd 1680) * $signed(input_fmap_154[7:0]) +
	( 15'sd 8966) * $signed(input_fmap_155[7:0]) +
	( 16'sd 16648) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9050) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4198) * $signed(input_fmap_159[7:0]) +
	( 13'sd 3504) * $signed(input_fmap_160[7:0]) +
	( 16'sd 24041) * $signed(input_fmap_161[7:0]) +
	( 16'sd 32536) * $signed(input_fmap_162[7:0]) +
	( 15'sd 9203) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19102) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28588) * $signed(input_fmap_165[7:0]) +
	( 16'sd 21451) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31483) * $signed(input_fmap_167[7:0]) +
	( 16'sd 23555) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18092) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2593) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7071) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22601) * $signed(input_fmap_172[7:0]) +
	( 16'sd 16437) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27883) * $signed(input_fmap_174[7:0]) +
	( 16'sd 30914) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13204) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18473) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22469) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5594) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23004) * $signed(input_fmap_180[7:0]) +
	( 16'sd 17960) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_182[7:0]) +
	( 16'sd 31934) * $signed(input_fmap_183[7:0]) +
	( 15'sd 12916) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25806) * $signed(input_fmap_185[7:0]) +
	( 16'sd 31348) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25391) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1393) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5097) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26316) * $signed(input_fmap_191[7:0]) +
	( 16'sd 26165) * $signed(input_fmap_192[7:0]) +
	( 14'sd 7726) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_194[7:0]) +
	( 15'sd 12336) * $signed(input_fmap_195[7:0]) +
	( 16'sd 21970) * $signed(input_fmap_196[7:0]) +
	( 14'sd 6750) * $signed(input_fmap_197[7:0]) +
	( 16'sd 26135) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28113) * $signed(input_fmap_199[7:0]) +
	( 15'sd 10929) * $signed(input_fmap_200[7:0]) +
	( 13'sd 2662) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5847) * $signed(input_fmap_202[7:0]) +
	( 15'sd 10354) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19044) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15006) * $signed(input_fmap_205[7:0]) +
	( 16'sd 24724) * $signed(input_fmap_206[7:0]) +
	( 16'sd 22757) * $signed(input_fmap_207[7:0]) +
	( 16'sd 26483) * $signed(input_fmap_208[7:0]) +
	( 15'sd 9023) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31034) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15589) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_212[7:0]) +
	( 11'sd 791) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7871) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9550) * $signed(input_fmap_215[7:0]) +
	( 16'sd 26020) * $signed(input_fmap_216[7:0]) +
	( 16'sd 27078) * $signed(input_fmap_217[7:0]) +
	( 11'sd 619) * $signed(input_fmap_218[7:0]) +
	( 16'sd 31350) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26396) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25796) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10390) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28972) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19112) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_225[7:0]) +
	( 16'sd 19148) * $signed(input_fmap_226[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4258) * $signed(input_fmap_228[7:0]) +
	( 16'sd 27928) * $signed(input_fmap_229[7:0]) +
	( 14'sd 5907) * $signed(input_fmap_230[7:0]) +
	( 16'sd 26666) * $signed(input_fmap_231[7:0]) +
	( 16'sd 23482) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28248) * $signed(input_fmap_233[7:0]) +
	( 16'sd 31886) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3028) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2581) * $signed(input_fmap_236[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_237[7:0]) +
	( 16'sd 18932) * $signed(input_fmap_238[7:0]) +
	( 16'sd 29255) * $signed(input_fmap_239[7:0]) +
	( 16'sd 20146) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32042) * $signed(input_fmap_241[7:0]) +
	( 13'sd 3264) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_243[7:0]) +
	( 16'sd 32541) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22351) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17753) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27159) * $signed(input_fmap_247[7:0]) +
	( 16'sd 27878) * $signed(input_fmap_248[7:0]) +
	( 16'sd 26252) * $signed(input_fmap_249[7:0]) +
	( 7'sd 35) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12154) * $signed(input_fmap_251[7:0]) +
	( 16'sd 23698) * $signed(input_fmap_252[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_253[7:0]) +
	( 16'sd 18431) * $signed(input_fmap_254[7:0]) +
	( 15'sd 8802) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_6;
assign conv_mac_6 = 
	( 16'sd 25462) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16248) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13875) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6565) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24014) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6116) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17842) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16016) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18693) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29435) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32132) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18726) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24315) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22729) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16603) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27173) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1441) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3626) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7212) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28659) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27915) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19271) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20348) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2896) * $signed(input_fmap_23[7:0]) +
	( 9'sd 141) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13530) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2348) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16527) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18023) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27668) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16592) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2196) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1646) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4463) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9884) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26120) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26111) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29215) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4355) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6674) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27099) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25445) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22047) * $signed(input_fmap_45[7:0]) +
	( 11'sd 705) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15661) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21693) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11917) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13236) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5229) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3172) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24552) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4784) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24900) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7706) * $signed(input_fmap_56[7:0]) +
	( 11'sd 534) * $signed(input_fmap_57[7:0]) +
	( 12'sd 2024) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20664) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17177) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15010) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22927) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13978) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19083) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2481) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22645) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29640) * $signed(input_fmap_69[7:0]) +
	( 7'sd 62) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24708) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23754) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5871) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22401) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22145) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16787) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16789) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30208) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31418) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28180) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16103) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15430) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27927) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5788) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31697) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7592) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19750) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1462) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8542) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3792) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10562) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9304) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19365) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26792) * $signed(input_fmap_97[7:0]) +
	( 10'sd 437) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23226) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24898) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7254) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3591) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14340) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10263) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12283) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14030) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8943) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10717) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21859) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26468) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18232) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30342) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19985) * $signed(input_fmap_114[7:0]) +
	( 11'sd 571) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19287) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13261) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32494) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5598) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19774) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19061) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21264) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5565) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4710) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24361) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8839) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7305) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25401) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20797) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14056) * $signed(input_fmap_132[7:0]) +
	( 15'sd 9969) * $signed(input_fmap_133[7:0]) +
	( 16'sd 30063) * $signed(input_fmap_134[7:0]) +
	( 13'sd 2425) * $signed(input_fmap_135[7:0]) +
	( 14'sd 8020) * $signed(input_fmap_136[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9974) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31418) * $signed(input_fmap_139[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_140[7:0]) +
	( 12'sd 1101) * $signed(input_fmap_141[7:0]) +
	( 15'sd 15871) * $signed(input_fmap_142[7:0]) +
	( 15'sd 15106) * $signed(input_fmap_143[7:0]) +
	( 15'sd 14430) * $signed(input_fmap_144[7:0]) +
	( 15'sd 11221) * $signed(input_fmap_145[7:0]) +
	( 15'sd 8546) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9365) * $signed(input_fmap_147[7:0]) +
	( 15'sd 8777) * $signed(input_fmap_148[7:0]) +
	( 16'sd 26987) * $signed(input_fmap_149[7:0]) +
	( 15'sd 14649) * $signed(input_fmap_150[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2741) * $signed(input_fmap_152[7:0]) +
	( 16'sd 28310) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30889) * $signed(input_fmap_154[7:0]) +
	( 14'sd 6603) * $signed(input_fmap_155[7:0]) +
	( 14'sd 4216) * $signed(input_fmap_156[7:0]) +
	( 14'sd 4475) * $signed(input_fmap_157[7:0]) +
	( 16'sd 16870) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32435) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18972) * $signed(input_fmap_160[7:0]) +
	( 13'sd 2524) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27785) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20446) * $signed(input_fmap_163[7:0]) +
	( 15'sd 15783) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9384) * $signed(input_fmap_165[7:0]) +
	( 16'sd 28808) * $signed(input_fmap_166[7:0]) +
	( 16'sd 28329) * $signed(input_fmap_167[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_168[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_169[7:0]) +
	( 16'sd 26679) * $signed(input_fmap_170[7:0]) +
	( 16'sd 23073) * $signed(input_fmap_171[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_172[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11130) * $signed(input_fmap_174[7:0]) +
	( 16'sd 20380) * $signed(input_fmap_175[7:0]) +
	( 16'sd 31055) * $signed(input_fmap_176[7:0]) +
	( 16'sd 23782) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31540) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18393) * $signed(input_fmap_179[7:0]) +
	( 15'sd 14773) * $signed(input_fmap_180[7:0]) +
	( 14'sd 7388) * $signed(input_fmap_181[7:0]) +
	( 15'sd 11868) * $signed(input_fmap_182[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24452) * $signed(input_fmap_184[7:0]) +
	( 15'sd 13934) * $signed(input_fmap_185[7:0]) +
	( 16'sd 19132) * $signed(input_fmap_186[7:0]) +
	( 16'sd 31597) * $signed(input_fmap_187[7:0]) +
	( 16'sd 30982) * $signed(input_fmap_188[7:0]) +
	( 15'sd 12887) * $signed(input_fmap_189[7:0]) +
	( 16'sd 18365) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5639) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15674) * $signed(input_fmap_192[7:0]) +
	( 16'sd 32198) * $signed(input_fmap_193[7:0]) +
	( 16'sd 17990) * $signed(input_fmap_194[7:0]) +
	( 16'sd 23460) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20345) * $signed(input_fmap_196[7:0]) +
	( 16'sd 30892) * $signed(input_fmap_197[7:0]) +
	( 14'sd 4903) * $signed(input_fmap_198[7:0]) +
	( 15'sd 13630) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_200[7:0]) +
	( 16'sd 19814) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7219) * $signed(input_fmap_202[7:0]) +
	( 14'sd 4158) * $signed(input_fmap_203[7:0]) +
	( 16'sd 18983) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11280) * $signed(input_fmap_205[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_206[7:0]) +
	( 16'sd 31012) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12135) * $signed(input_fmap_208[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_209[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_210[7:0]) +
	( 16'sd 16689) * $signed(input_fmap_211[7:0]) +
	( 16'sd 32234) * $signed(input_fmap_212[7:0]) +
	( 15'sd 10897) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_214[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_215[7:0]) +
	( 14'sd 8181) * $signed(input_fmap_216[7:0]) +
	( 14'sd 6536) * $signed(input_fmap_217[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15549) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_220[7:0]) +
	( 16'sd 29034) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14060) * $signed(input_fmap_222[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_223[7:0]) +
	( 16'sd 18025) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2567) * $signed(input_fmap_225[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_226[7:0]) +
	( 15'sd 10758) * $signed(input_fmap_227[7:0]) +
	( 16'sd 27176) * $signed(input_fmap_228[7:0]) +
	( 16'sd 27602) * $signed(input_fmap_229[7:0]) +
	( 9'sd 141) * $signed(input_fmap_230[7:0]) +
	( 16'sd 23306) * $signed(input_fmap_231[7:0]) +
	( 16'sd 19356) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11739) * $signed(input_fmap_233[7:0]) +
	( 16'sd 28652) * $signed(input_fmap_234[7:0]) +
	( 16'sd 24263) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25383) * $signed(input_fmap_236[7:0]) +
	( 16'sd 31885) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19344) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23657) * $signed(input_fmap_239[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_240[7:0]) +
	( 16'sd 22721) * $signed(input_fmap_241[7:0]) +
	( 16'sd 30181) * $signed(input_fmap_242[7:0]) +
	( 16'sd 27914) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6269) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5912) * $signed(input_fmap_245[7:0]) +
	( 15'sd 13918) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3837) * $signed(input_fmap_247[7:0]) +
	( 13'sd 2640) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15769) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24605) * $signed(input_fmap_250[7:0]) +
	( 14'sd 5714) * $signed(input_fmap_251[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13959) * $signed(input_fmap_253[7:0]) +
	( 16'sd 29873) * $signed(input_fmap_254[7:0]) +
	( 16'sd 25661) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_7;
assign conv_mac_7 = 
	( 16'sd 28599) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8400) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6959) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12478) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25760) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9072) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20658) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26417) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22444) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7298) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19280) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20060) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17539) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17076) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32763) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31661) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32282) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11692) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19676) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31741) * $signed(input_fmap_22[7:0]) +
	( 13'sd 4061) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11016) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12522) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1271) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31074) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12081) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29290) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11404) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3939) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8428) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17941) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15730) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1515) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3474) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26650) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16308) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15307) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16628) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25223) * $signed(input_fmap_43[7:0]) +
	( 7'sd 55) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8533) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30887) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17737) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11922) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20206) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11272) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10649) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14265) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18582) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25829) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12915) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21112) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30512) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31754) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2125) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15875) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10802) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32187) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28342) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26460) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25993) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1837) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16003) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30503) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5731) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23470) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9065) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16915) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5698) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18385) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1704) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30345) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28219) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17501) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21728) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10873) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29606) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10226) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12833) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15009) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19448) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25679) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31003) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17724) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7294) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13495) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27819) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26346) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13912) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21879) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2754) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30507) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23958) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26314) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21365) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19163) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29283) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22164) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28158) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26834) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11971) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23120) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15416) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11090) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13059) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8237) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27203) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14852) * $signed(input_fmap_130[7:0]) +
	( 15'sd 11523) * $signed(input_fmap_131[7:0]) +
	( 15'sd 9505) * $signed(input_fmap_132[7:0]) +
	( 12'sd 1932) * $signed(input_fmap_133[7:0]) +
	( 16'sd 29151) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18039) * $signed(input_fmap_135[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24839) * $signed(input_fmap_137[7:0]) +
	( 13'sd 3018) * $signed(input_fmap_138[7:0]) +
	( 15'sd 12990) * $signed(input_fmap_139[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14152) * $signed(input_fmap_142[7:0]) +
	( 15'sd 16116) * $signed(input_fmap_143[7:0]) +
	( 16'sd 25216) * $signed(input_fmap_144[7:0]) +
	( 15'sd 9981) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24968) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_147[7:0]) +
	( 16'sd 25830) * $signed(input_fmap_148[7:0]) +
	( 16'sd 26299) * $signed(input_fmap_149[7:0]) +
	( 16'sd 20850) * $signed(input_fmap_150[7:0]) +
	( 16'sd 22237) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20857) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31869) * $signed(input_fmap_153[7:0]) +
	( 15'sd 9962) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27428) * $signed(input_fmap_155[7:0]) +
	( 15'sd 11543) * $signed(input_fmap_156[7:0]) +
	( 13'sd 2477) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1453) * $signed(input_fmap_158[7:0]) +
	( 16'sd 29813) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24544) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4269) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2961) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8336) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3790) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9656) * $signed(input_fmap_165[7:0]) +
	( 16'sd 25532) * $signed(input_fmap_166[7:0]) +
	( 13'sd 2979) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20679) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21642) * $signed(input_fmap_169[7:0]) +
	( 11'sd 718) * $signed(input_fmap_170[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_171[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_172[7:0]) +
	( 13'sd 2155) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16859) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25320) * $signed(input_fmap_175[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1776) * $signed(input_fmap_177[7:0]) +
	( 16'sd 29666) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28568) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21902) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18046) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10408) * $signed(input_fmap_182[7:0]) +
	( 16'sd 28197) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30566) * $signed(input_fmap_184[7:0]) +
	( 14'sd 4102) * $signed(input_fmap_185[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_186[7:0]) +
	( 16'sd 23489) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21923) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11089) * $signed(input_fmap_189[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20624) * $signed(input_fmap_192[7:0]) +
	( 16'sd 25846) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30164) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24418) * $signed(input_fmap_195[7:0]) +
	( 16'sd 18495) * $signed(input_fmap_196[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24716) * $signed(input_fmap_198[7:0]) +
	( 15'sd 13506) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31963) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21659) * $signed(input_fmap_201[7:0]) +
	( 16'sd 23000) * $signed(input_fmap_202[7:0]) +
	( 16'sd 20301) * $signed(input_fmap_203[7:0]) +
	( 13'sd 3838) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1545) * $signed(input_fmap_205[7:0]) +
	( 12'sd 1294) * $signed(input_fmap_206[7:0]) +
	( 16'sd 31789) * $signed(input_fmap_207[7:0]) +
	( 11'sd 629) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19675) * $signed(input_fmap_209[7:0]) +
	( 14'sd 6099) * $signed(input_fmap_210[7:0]) +
	( 16'sd 21405) * $signed(input_fmap_211[7:0]) +
	( 11'sd 660) * $signed(input_fmap_212[7:0]) +
	( 15'sd 10628) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20218) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17293) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19148) * $signed(input_fmap_216[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_217[7:0]) +
	( 16'sd 18652) * $signed(input_fmap_218[7:0]) +
	( 16'sd 27802) * $signed(input_fmap_219[7:0]) +
	( 15'sd 11393) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19827) * $signed(input_fmap_221[7:0]) +
	( 16'sd 22916) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22938) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1238) * $signed(input_fmap_224[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_225[7:0]) +
	( 15'sd 16051) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5721) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2083) * $signed(input_fmap_228[7:0]) +
	( 14'sd 7409) * $signed(input_fmap_229[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_230[7:0]) +
	( 14'sd 6342) * $signed(input_fmap_231[7:0]) +
	( 16'sd 23550) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5759) * $signed(input_fmap_233[7:0]) +
	( 16'sd 21733) * $signed(input_fmap_234[7:0]) +
	( 15'sd 15094) * $signed(input_fmap_235[7:0]) +
	( 16'sd 19939) * $signed(input_fmap_236[7:0]) +
	( 16'sd 32687) * $signed(input_fmap_237[7:0]) +
	( 13'sd 2331) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_239[7:0]) +
	( 13'sd 2563) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18376) * $signed(input_fmap_241[7:0]) +
	( 16'sd 18691) * $signed(input_fmap_242[7:0]) +
	( 16'sd 26422) * $signed(input_fmap_243[7:0]) +
	( 14'sd 5049) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30913) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23230) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27993) * $signed(input_fmap_247[7:0]) +
	( 15'sd 12246) * $signed(input_fmap_248[7:0]) +
	( 14'sd 7901) * $signed(input_fmap_249[7:0]) +
	( 15'sd 11087) * $signed(input_fmap_250[7:0]) +
	( 16'sd 24497) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20633) * $signed(input_fmap_254[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_8;
assign conv_mac_8 = 
	( 16'sd 24188) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11331) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1330) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2400) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11437) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22253) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22141) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16729) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5740) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29892) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2079) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18919) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19474) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21336) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30960) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28975) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16201) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10372) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15496) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14678) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7266) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8687) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13040) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23306) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27997) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14589) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17167) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26256) * $signed(input_fmap_31[7:0]) +
	( 11'sd 538) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19750) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8989) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29877) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8768) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9962) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21683) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15767) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32592) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27182) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23049) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12959) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29935) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26880) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9645) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2654) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22809) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4582) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6871) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5764) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9134) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30078) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30219) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30197) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9097) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14523) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5288) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20645) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25064) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12812) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8621) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31710) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17648) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21932) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11815) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1553) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30309) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26787) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1522) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14095) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25866) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18318) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32723) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1062) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5210) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30683) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23725) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19086) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9057) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3378) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27846) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22253) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4312) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27570) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5254) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24993) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31184) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23221) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10341) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9865) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20949) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22203) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24751) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12965) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29875) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1889) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4830) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29592) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32265) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30153) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29942) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3616) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27954) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17386) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21704) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29926) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3205) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23471) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18159) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23456) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21837) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32098) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21917) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24394) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32102) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20030) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_127[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_128[7:0]) +
	( 14'sd 4592) * $signed(input_fmap_129[7:0]) +
	( 16'sd 17645) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23256) * $signed(input_fmap_131[7:0]) +
	( 16'sd 21584) * $signed(input_fmap_132[7:0]) +
	( 13'sd 3514) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32344) * $signed(input_fmap_134[7:0]) +
	( 16'sd 30127) * $signed(input_fmap_135[7:0]) +
	( 16'sd 24212) * $signed(input_fmap_136[7:0]) +
	( 11'sd 881) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31621) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24075) * $signed(input_fmap_139[7:0]) +
	( 16'sd 27207) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5989) * $signed(input_fmap_141[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5498) * $signed(input_fmap_143[7:0]) +
	( 16'sd 27821) * $signed(input_fmap_144[7:0]) +
	( 12'sd 1650) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19014) * $signed(input_fmap_146[7:0]) +
	( 15'sd 16201) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26200) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17921) * $signed(input_fmap_149[7:0]) +
	( 13'sd 3919) * $signed(input_fmap_150[7:0]) +
	( 16'sd 31547) * $signed(input_fmap_151[7:0]) +
	( 16'sd 32284) * $signed(input_fmap_152[7:0]) +
	( 11'sd 624) * $signed(input_fmap_153[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30805) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28435) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25076) * $signed(input_fmap_157[7:0]) +
	( 16'sd 22668) * $signed(input_fmap_158[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_159[7:0]) +
	( 16'sd 30259) * $signed(input_fmap_160[7:0]) +
	( 16'sd 29452) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3622) * $signed(input_fmap_163[7:0]) +
	( 15'sd 14615) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22638) * $signed(input_fmap_165[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_166[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_167[7:0]) +
	( 16'sd 22995) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18723) * $signed(input_fmap_170[7:0]) +
	( 14'sd 5401) * $signed(input_fmap_171[7:0]) +
	( 15'sd 10306) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18061) * $signed(input_fmap_173[7:0]) +
	( 16'sd 21917) * $signed(input_fmap_174[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_175[7:0]) +
	( 16'sd 30439) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1627) * $signed(input_fmap_177[7:0]) +
	( 16'sd 21402) * $signed(input_fmap_178[7:0]) +
	( 15'sd 12269) * $signed(input_fmap_179[7:0]) +
	( 15'sd 14718) * $signed(input_fmap_180[7:0]) +
	( 16'sd 21018) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6317) * $signed(input_fmap_182[7:0]) +
	( 16'sd 18782) * $signed(input_fmap_183[7:0]) +
	( 16'sd 16545) * $signed(input_fmap_184[7:0]) +
	( 11'sd 650) * $signed(input_fmap_185[7:0]) +
	( 15'sd 16027) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18422) * $signed(input_fmap_187[7:0]) +
	( 16'sd 28249) * $signed(input_fmap_188[7:0]) +
	( 16'sd 24603) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4289) * $signed(input_fmap_190[7:0]) +
	( 16'sd 21660) * $signed(input_fmap_191[7:0]) +
	( 16'sd 25924) * $signed(input_fmap_192[7:0]) +
	( 15'sd 16047) * $signed(input_fmap_193[7:0]) +
	( 16'sd 32611) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19054) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24739) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1392) * $signed(input_fmap_197[7:0]) +
	( 8'sd 103) * $signed(input_fmap_198[7:0]) +
	( 16'sd 17302) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5121) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_201[7:0]) +
	( 16'sd 25580) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25338) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4564) * $signed(input_fmap_204[7:0]) +
	( 15'sd 16187) * $signed(input_fmap_205[7:0]) +
	( 15'sd 16252) * $signed(input_fmap_206[7:0]) +
	( 15'sd 8399) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7614) * $signed(input_fmap_209[7:0]) +
	( 15'sd 12731) * $signed(input_fmap_210[7:0]) +
	( 14'sd 8007) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11750) * $signed(input_fmap_212[7:0]) +
	( 16'sd 27192) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1489) * $signed(input_fmap_214[7:0]) +
	( 14'sd 4910) * $signed(input_fmap_215[7:0]) +
	( 15'sd 15698) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_217[7:0]) +
	( 16'sd 32465) * $signed(input_fmap_218[7:0]) +
	( 16'sd 27793) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25333) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28400) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15327) * $signed(input_fmap_222[7:0]) +
	( 15'sd 10672) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7176) * $signed(input_fmap_224[7:0]) +
	( 16'sd 22157) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6451) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24351) * $signed(input_fmap_227[7:0]) +
	( 16'sd 27133) * $signed(input_fmap_228[7:0]) +
	( 15'sd 9833) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18194) * $signed(input_fmap_230[7:0]) +
	( 13'sd 2556) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29526) * $signed(input_fmap_232[7:0]) +
	( 14'sd 4906) * $signed(input_fmap_233[7:0]) +
	( 16'sd 32742) * $signed(input_fmap_234[7:0]) +
	( 15'sd 9883) * $signed(input_fmap_235[7:0]) +
	( 15'sd 8969) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2940) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12960) * $signed(input_fmap_238[7:0]) +
	( 15'sd 14159) * $signed(input_fmap_239[7:0]) +
	( 16'sd 24589) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23065) * $signed(input_fmap_241[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22960) * $signed(input_fmap_244[7:0]) +
	( 16'sd 16957) * $signed(input_fmap_245[7:0]) +
	( 13'sd 2295) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3735) * $signed(input_fmap_247[7:0]) +
	( 16'sd 29781) * $signed(input_fmap_248[7:0]) +
	( 12'sd 1977) * $signed(input_fmap_249[7:0]) +
	( 13'sd 2578) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22801) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30161) * $signed(input_fmap_252[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_253[7:0]) +
	( 14'sd 7359) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5197) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_9;
assign conv_mac_9 = 
	( 16'sd 26831) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22303) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26573) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8299) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26240) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2793) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25742) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14286) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6298) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15095) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21393) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21095) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27772) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16415) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5163) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16175) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27286) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17780) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_22[7:0]) +
	( 11'sd 729) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2424) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4540) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15391) * $signed(input_fmap_26[7:0]) +
	( 8'sd 72) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1265) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29931) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8443) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12997) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32527) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31034) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5168) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21361) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11768) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6913) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30386) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31649) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14905) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4163) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15420) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32004) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18781) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24462) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3810) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6078) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24528) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9112) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2431) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30094) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32069) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17105) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29000) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29480) * $signed(input_fmap_58[7:0]) +
	( 7'sd 63) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27800) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26543) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4836) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1760) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11684) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15229) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12075) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9624) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4255) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7644) * $signed(input_fmap_70[7:0]) +
	( 10'sd 429) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19505) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29176) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2701) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32735) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4825) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23342) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5728) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22285) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19680) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8502) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30019) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10353) * $signed(input_fmap_87[7:0]) +
	( 8'sd 106) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23376) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22649) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28931) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25606) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14531) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13503) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17046) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12792) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14512) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13720) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5495) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15182) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15602) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7134) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9739) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6018) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7974) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10540) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17559) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19849) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30699) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21170) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24238) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31340) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5676) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5050) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27879) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16944) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16837) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3569) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29885) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20991) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31158) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6742) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3529) * $signed(input_fmap_127[7:0]) +
	( 15'sd 12906) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_129[7:0]) +
	( 15'sd 8242) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15979) * $signed(input_fmap_131[7:0]) +
	( 16'sd 30043) * $signed(input_fmap_132[7:0]) +
	( 16'sd 32503) * $signed(input_fmap_133[7:0]) +
	( 15'sd 15332) * $signed(input_fmap_134[7:0]) +
	( 14'sd 5070) * $signed(input_fmap_135[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_137[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18324) * $signed(input_fmap_139[7:0]) +
	( 16'sd 20221) * $signed(input_fmap_140[7:0]) +
	( 16'sd 32338) * $signed(input_fmap_141[7:0]) +
	( 15'sd 13581) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10661) * $signed(input_fmap_143[7:0]) +
	( 16'sd 32633) * $signed(input_fmap_144[7:0]) +
	( 15'sd 15240) * $signed(input_fmap_145[7:0]) +
	( 16'sd 26848) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_147[7:0]) +
	( 15'sd 14935) * $signed(input_fmap_148[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_149[7:0]) +
	( 16'sd 19492) * $signed(input_fmap_150[7:0]) +
	( 14'sd 5694) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29648) * $signed(input_fmap_152[7:0]) +
	( 15'sd 15923) * $signed(input_fmap_153[7:0]) +
	( 16'sd 27111) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_155[7:0]) +
	( 14'sd 4303) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31006) * $signed(input_fmap_157[7:0]) +
	( 15'sd 14486) * $signed(input_fmap_158[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_159[7:0]) +
	( 7'sd 59) * $signed(input_fmap_160[7:0]) +
	( 15'sd 9252) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4867) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32439) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3505) * $signed(input_fmap_164[7:0]) +
	( 14'sd 7225) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_166[7:0]) +
	( 16'sd 18942) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29148) * $signed(input_fmap_168[7:0]) +
	( 15'sd 15186) * $signed(input_fmap_169[7:0]) +
	( 12'sd 1484) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_171[7:0]) +
	( 16'sd 25798) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12914) * $signed(input_fmap_173[7:0]) +
	( 16'sd 17300) * $signed(input_fmap_174[7:0]) +
	( 15'sd 14683) * $signed(input_fmap_175[7:0]) +
	( 14'sd 4873) * $signed(input_fmap_176[7:0]) +
	( 14'sd 4377) * $signed(input_fmap_177[7:0]) +
	( 16'sd 21860) * $signed(input_fmap_178[7:0]) +
	( 15'sd 8688) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26687) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15660) * $signed(input_fmap_181[7:0]) +
	( 16'sd 27163) * $signed(input_fmap_182[7:0]) +
	( 15'sd 14336) * $signed(input_fmap_183[7:0]) +
	( 16'sd 25137) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27519) * $signed(input_fmap_185[7:0]) +
	( 12'sd 1383) * $signed(input_fmap_186[7:0]) +
	( 16'sd 29064) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17770) * $signed(input_fmap_188[7:0]) +
	( 16'sd 28130) * $signed(input_fmap_189[7:0]) +
	( 15'sd 12670) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29450) * $signed(input_fmap_191[7:0]) +
	( 16'sd 26736) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6584) * $signed(input_fmap_193[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_194[7:0]) +
	( 15'sd 11608) * $signed(input_fmap_195[7:0]) +
	( 16'sd 23668) * $signed(input_fmap_196[7:0]) +
	( 13'sd 3382) * $signed(input_fmap_197[7:0]) +
	( 16'sd 16675) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14363) * $signed(input_fmap_199[7:0]) +
	( 16'sd 24670) * $signed(input_fmap_200[7:0]) +
	( 14'sd 7638) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21670) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15566) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30600) * $signed(input_fmap_205[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7740) * $signed(input_fmap_207[7:0]) +
	( 12'sd 1825) * $signed(input_fmap_208[7:0]) +
	( 11'sd 779) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30262) * $signed(input_fmap_210[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_211[7:0]) +
	( 16'sd 32510) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23838) * $signed(input_fmap_213[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9233) * $signed(input_fmap_215[7:0]) +
	( 15'sd 12950) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30110) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10090) * $signed(input_fmap_218[7:0]) +
	( 15'sd 9500) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25973) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22737) * $signed(input_fmap_223[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_225[7:0]) +
	( 10'sd 383) * $signed(input_fmap_226[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_227[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_228[7:0]) +
	( 12'sd 1109) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15604) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7277) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_232[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_233[7:0]) +
	( 15'sd 10095) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3119) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31277) * $signed(input_fmap_236[7:0]) +
	( 16'sd 26105) * $signed(input_fmap_237[7:0]) +
	( 14'sd 7866) * $signed(input_fmap_238[7:0]) +
	( 16'sd 25064) * $signed(input_fmap_239[7:0]) +
	( 15'sd 8389) * $signed(input_fmap_240[7:0]) +
	( 16'sd 24943) * $signed(input_fmap_241[7:0]) +
	( 13'sd 2304) * $signed(input_fmap_242[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_243[7:0]) +
	( 16'sd 26282) * $signed(input_fmap_244[7:0]) +
	( 16'sd 29858) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15971) * $signed(input_fmap_246[7:0]) +
	( 10'sd 382) * $signed(input_fmap_247[7:0]) +
	( 15'sd 9740) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2870) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3816) * $signed(input_fmap_250[7:0]) +
	( 16'sd 23541) * $signed(input_fmap_251[7:0]) +
	( 16'sd 24890) * $signed(input_fmap_252[7:0]) +
	( 9'sd 152) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5699) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5275) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_10;
assign conv_mac_10 = 
	( 14'sd 4509) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26027) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20295) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28578) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3973) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1569) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1747) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19735) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4907) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12516) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5026) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17182) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10102) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28418) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29877) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13219) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25871) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14002) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29947) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14783) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3018) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16736) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11596) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18196) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21932) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2141) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5701) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8407) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19449) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13003) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20064) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18642) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2453) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18342) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26581) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12918) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4593) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15861) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21772) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20083) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13713) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13516) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27918) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26844) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9668) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8790) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28781) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2588) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7823) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20580) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6955) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14692) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20115) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9026) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15943) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18333) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24396) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28212) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6629) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9693) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15029) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26890) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3373) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16263) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7984) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27334) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27957) * $signed(input_fmap_71[7:0]) +
	( 11'sd 997) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7574) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26433) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11946) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24631) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19227) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24279) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18769) * $signed(input_fmap_81[7:0]) +
	( 10'sd 382) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9181) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17484) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18097) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6620) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9874) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4715) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2761) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29559) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7387) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32020) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1488) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28301) * $signed(input_fmap_95[7:0]) +
	( 10'sd 438) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17668) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24647) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28445) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5221) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29964) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22159) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18974) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2058) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22256) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6098) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10412) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26022) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1077) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31820) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18162) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1340) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7785) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23423) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12465) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21997) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32391) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3838) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7960) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21504) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9588) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22527) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7975) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32447) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32073) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7505) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23872) * $signed(input_fmap_128[7:0]) +
	( 16'sd 21025) * $signed(input_fmap_129[7:0]) +
	( 13'sd 2337) * $signed(input_fmap_130[7:0]) +
	( 16'sd 17395) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11596) * $signed(input_fmap_132[7:0]) +
	( 13'sd 2938) * $signed(input_fmap_133[7:0]) +
	( 16'sd 27390) * $signed(input_fmap_134[7:0]) +
	( 14'sd 7390) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2467) * $signed(input_fmap_136[7:0]) +
	( 16'sd 17481) * $signed(input_fmap_137[7:0]) +
	( 16'sd 26964) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2399) * $signed(input_fmap_139[7:0]) +
	( 16'sd 21964) * $signed(input_fmap_140[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21166) * $signed(input_fmap_142[7:0]) +
	( 16'sd 16795) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13368) * $signed(input_fmap_144[7:0]) +
	( 15'sd 12132) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3083) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18241) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21616) * $signed(input_fmap_148[7:0]) +
	( 15'sd 8714) * $signed(input_fmap_149[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24775) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14524) * $signed(input_fmap_152[7:0]) +
	( 16'sd 18784) * $signed(input_fmap_153[7:0]) +
	( 11'sd 987) * $signed(input_fmap_154[7:0]) +
	( 16'sd 25702) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_157[7:0]) +
	( 16'sd 24535) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4720) * $signed(input_fmap_159[7:0]) +
	( 15'sd 8260) * $signed(input_fmap_160[7:0]) +
	( 15'sd 8800) * $signed(input_fmap_161[7:0]) +
	( 14'sd 7272) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20564) * $signed(input_fmap_163[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10254) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8449) * $signed(input_fmap_166[7:0]) +
	( 15'sd 12759) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17681) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18478) * $signed(input_fmap_169[7:0]) +
	( 16'sd 30178) * $signed(input_fmap_170[7:0]) +
	( 12'sd 1506) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7257) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23935) * $signed(input_fmap_173[7:0]) +
	( 13'sd 2809) * $signed(input_fmap_174[7:0]) +
	( 15'sd 11523) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10866) * $signed(input_fmap_176[7:0]) +
	( 16'sd 17599) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32309) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18616) * $signed(input_fmap_179[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_180[7:0]) +
	( 16'sd 24900) * $signed(input_fmap_181[7:0]) +
	( 16'sd 23763) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5015) * $signed(input_fmap_183[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27883) * $signed(input_fmap_185[7:0]) +
	( 16'sd 19194) * $signed(input_fmap_186[7:0]) +
	( 16'sd 20208) * $signed(input_fmap_187[7:0]) +
	( 15'sd 8704) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11028) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31098) * $signed(input_fmap_190[7:0]) +
	( 16'sd 16523) * $signed(input_fmap_191[7:0]) +
	( 11'sd 972) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11315) * $signed(input_fmap_193[7:0]) +
	( 15'sd 11236) * $signed(input_fmap_194[7:0]) +
	( 16'sd 18716) * $signed(input_fmap_195[7:0]) +
	( 12'sd 1199) * $signed(input_fmap_196[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2758) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12085) * $signed(input_fmap_199[7:0]) +
	( 16'sd 16744) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13249) * $signed(input_fmap_201[7:0]) +
	( 16'sd 28634) * $signed(input_fmap_202[7:0]) +
	( 16'sd 17819) * $signed(input_fmap_203[7:0]) +
	( 16'sd 21294) * $signed(input_fmap_204[7:0]) +
	( 15'sd 13302) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27799) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13763) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30335) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7900) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10543) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3037) * $signed(input_fmap_211[7:0]) +
	( 16'sd 22658) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2647) * $signed(input_fmap_213[7:0]) +
	( 15'sd 16314) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2216) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11976) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17345) * $signed(input_fmap_217[7:0]) +
	( 16'sd 32503) * $signed(input_fmap_218[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_219[7:0]) +
	( 15'sd 10258) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27640) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18822) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17434) * $signed(input_fmap_223[7:0]) +
	( 16'sd 20502) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14002) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20357) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8764) * $signed(input_fmap_228[7:0]) +
	( 16'sd 25733) * $signed(input_fmap_229[7:0]) +
	( 15'sd 13985) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7532) * $signed(input_fmap_231[7:0]) +
	( 10'sd 374) * $signed(input_fmap_232[7:0]) +
	( 11'sd 824) * $signed(input_fmap_233[7:0]) +
	( 16'sd 31964) * $signed(input_fmap_234[7:0]) +
	( 15'sd 15497) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28986) * $signed(input_fmap_236[7:0]) +
	( 16'sd 17310) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5669) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_239[7:0]) +
	( 15'sd 14623) * $signed(input_fmap_240[7:0]) +
	( 16'sd 19539) * $signed(input_fmap_241[7:0]) +
	( 16'sd 20700) * $signed(input_fmap_242[7:0]) +
	( 15'sd 11026) * $signed(input_fmap_243[7:0]) +
	( 16'sd 16929) * $signed(input_fmap_244[7:0]) +
	( 16'sd 18370) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22864) * $signed(input_fmap_246[7:0]) +
	( 16'sd 24928) * $signed(input_fmap_247[7:0]) +
	( 13'sd 2984) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14030) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24831) * $signed(input_fmap_250[7:0]) +
	( 15'sd 10915) * $signed(input_fmap_251[7:0]) +
	( 13'sd 3916) * $signed(input_fmap_252[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_253[7:0]) +
	( 15'sd 16309) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5669) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_11;
assign conv_mac_11 = 
	( 16'sd 24633) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29977) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17081) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4886) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3070) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17032) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13283) * $signed(input_fmap_9[7:0]) +
	( 11'sd 938) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16560) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28974) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30745) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30399) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23249) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19815) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29426) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32619) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27573) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11631) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23525) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14394) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21861) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28610) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1299) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4494) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21632) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32103) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25669) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16697) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1954) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3481) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27611) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9774) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15511) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12237) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25426) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22031) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10633) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28898) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20913) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4977) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2837) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11480) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15578) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1907) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3061) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31758) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28020) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24875) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1304) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29856) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22666) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20297) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19276) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22889) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8715) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29148) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17782) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30083) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20406) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9346) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28145) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2067) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28427) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18004) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28150) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10389) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4754) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11500) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8106) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22020) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10075) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3727) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1921) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5828) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6974) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2461) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10908) * $signed(input_fmap_90[7:0]) +
	( 12'sd 2008) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6439) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21930) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14592) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29010) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4796) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31035) * $signed(input_fmap_97[7:0]) +
	( 11'sd 997) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24557) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16840) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10281) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31341) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14423) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12935) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2734) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27455) * $signed(input_fmap_109[7:0]) +
	( 11'sd 693) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11221) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12004) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10626) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7216) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15768) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18571) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12704) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31101) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31677) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8641) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8428) * $signed(input_fmap_123[7:0]) +
	( 8'sd 120) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_125[7:0]) +
	( 10'sd 400) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4659) * $signed(input_fmap_127[7:0]) +
	( 16'sd 32334) * $signed(input_fmap_128[7:0]) +
	( 11'sd 876) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14609) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23763) * $signed(input_fmap_131[7:0]) +
	( 16'sd 17590) * $signed(input_fmap_132[7:0]) +
	( 16'sd 32013) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31329) * $signed(input_fmap_134[7:0]) +
	( 16'sd 29222) * $signed(input_fmap_135[7:0]) +
	( 13'sd 3930) * $signed(input_fmap_136[7:0]) +
	( 14'sd 7632) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2097) * $signed(input_fmap_139[7:0]) +
	( 15'sd 12576) * $signed(input_fmap_140[7:0]) +
	( 14'sd 6715) * $signed(input_fmap_141[7:0]) +
	( 10'sd 450) * $signed(input_fmap_142[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28889) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24774) * $signed(input_fmap_146[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_147[7:0]) +
	( 15'sd 9074) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7283) * $signed(input_fmap_149[7:0]) +
	( 16'sd 32712) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19348) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6633) * $signed(input_fmap_152[7:0]) +
	( 16'sd 16822) * $signed(input_fmap_153[7:0]) +
	( 12'sd 1864) * $signed(input_fmap_154[7:0]) +
	( 16'sd 21265) * $signed(input_fmap_155[7:0]) +
	( 12'sd 1802) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23525) * $signed(input_fmap_157[7:0]) +
	( 16'sd 31908) * $signed(input_fmap_158[7:0]) +
	( 15'sd 11412) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11649) * $signed(input_fmap_160[7:0]) +
	( 16'sd 25692) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30705) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24615) * $signed(input_fmap_163[7:0]) +
	( 14'sd 7822) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23770) * $signed(input_fmap_165[7:0]) +
	( 15'sd 16349) * $signed(input_fmap_166[7:0]) +
	( 16'sd 16401) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17590) * $signed(input_fmap_168[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17586) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20224) * $signed(input_fmap_171[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27734) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16499) * $signed(input_fmap_174[7:0]) +
	( 16'sd 18331) * $signed(input_fmap_175[7:0]) +
	( 14'sd 4285) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19936) * $signed(input_fmap_177[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_178[7:0]) +
	( 10'sd 385) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32490) * $signed(input_fmap_180[7:0]) +
	( 12'sd 1165) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16635) * $signed(input_fmap_182[7:0]) +
	( 16'sd 31538) * $signed(input_fmap_183[7:0]) +
	( 15'sd 15737) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22523) * $signed(input_fmap_185[7:0]) +
	( 16'sd 32146) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4536) * $signed(input_fmap_187[7:0]) +
	( 15'sd 8374) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25360) * $signed(input_fmap_189[7:0]) +
	( 16'sd 29268) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24546) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29652) * $signed(input_fmap_192[7:0]) +
	( 15'sd 14737) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9672) * $signed(input_fmap_194[7:0]) +
	( 13'sd 2442) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24921) * $signed(input_fmap_196[7:0]) +
	( 14'sd 6708) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27969) * $signed(input_fmap_198[7:0]) +
	( 16'sd 27836) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_200[7:0]) +
	( 16'sd 17209) * $signed(input_fmap_201[7:0]) +
	( 16'sd 20453) * $signed(input_fmap_202[7:0]) +
	( 16'sd 27459) * $signed(input_fmap_203[7:0]) +
	( 16'sd 20155) * $signed(input_fmap_204[7:0]) +
	( 16'sd 19665) * $signed(input_fmap_205[7:0]) +
	( 16'sd 24091) * $signed(input_fmap_206[7:0]) +
	( 16'sd 32290) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6741) * $signed(input_fmap_208[7:0]) +
	( 16'sd 21786) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18330) * $signed(input_fmap_210[7:0]) +
	( 16'sd 21955) * $signed(input_fmap_211[7:0]) +
	( 14'sd 5168) * $signed(input_fmap_212[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30117) * $signed(input_fmap_214[7:0]) +
	( 15'sd 14566) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23967) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24732) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7278) * $signed(input_fmap_218[7:0]) +
	( 15'sd 11616) * $signed(input_fmap_219[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_220[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2664) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25318) * $signed(input_fmap_223[7:0]) +
	( 13'sd 4061) * $signed(input_fmap_224[7:0]) +
	( 14'sd 4986) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7550) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9946) * $signed(input_fmap_227[7:0]) +
	( 16'sd 16872) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24990) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27996) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10580) * $signed(input_fmap_231[7:0]) +
	( 16'sd 19758) * $signed(input_fmap_232[7:0]) +
	( 13'sd 2189) * $signed(input_fmap_233[7:0]) +
	( 15'sd 10694) * $signed(input_fmap_234[7:0]) +
	( 16'sd 25958) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31623) * $signed(input_fmap_236[7:0]) +
	( 10'sd 275) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13070) * $signed(input_fmap_238[7:0]) +
	( 14'sd 6422) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26824) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32160) * $signed(input_fmap_241[7:0]) +
	( 14'sd 6259) * $signed(input_fmap_242[7:0]) +
	( 15'sd 12987) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22315) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19814) * $signed(input_fmap_245[7:0]) +
	( 16'sd 27220) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21376) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10285) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28973) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22929) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2676) * $signed(input_fmap_251[7:0]) +
	( 11'sd 771) * $signed(input_fmap_252[7:0]) +
	( 15'sd 14025) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26001) * $signed(input_fmap_254[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_12;
assign conv_mac_12 = 
	( 16'sd 22467) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1825) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30688) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9164) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4383) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11020) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12624) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16289) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13743) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21939) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30596) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9800) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24816) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4872) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24537) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15950) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25706) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20129) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21058) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19569) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18587) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18415) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32475) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32738) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26973) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17072) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2965) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8685) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15669) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10546) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5687) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7682) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9226) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20288) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15427) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30392) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27915) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2826) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20569) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2271) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13302) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16634) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5994) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31780) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16324) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2432) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14414) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31280) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20248) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30007) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31411) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19624) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30161) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14452) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24855) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18532) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20099) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30268) * $signed(input_fmap_67[7:0]) +
	( 10'sd 272) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28136) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14915) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2391) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19562) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9032) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12507) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22027) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16157) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13306) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19657) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15006) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17278) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6389) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2184) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27983) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29098) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13212) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5274) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2831) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32514) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7664) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9305) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3720) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26625) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30307) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21033) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13476) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17265) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3507) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17726) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10488) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2165) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12943) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28002) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8615) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22800) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7646) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15308) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18436) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3727) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14902) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2747) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30245) * $signed(input_fmap_117[7:0]) +
	( 11'sd 736) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8839) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25228) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20142) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9473) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16645) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1333) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28003) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24052) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_127[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13395) * $signed(input_fmap_129[7:0]) +
	( 13'sd 2668) * $signed(input_fmap_130[7:0]) +
	( 15'sd 12739) * $signed(input_fmap_131[7:0]) +
	( 16'sd 23922) * $signed(input_fmap_132[7:0]) +
	( 16'sd 30681) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5294) * $signed(input_fmap_134[7:0]) +
	( 16'sd 30340) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31155) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25903) * $signed(input_fmap_137[7:0]) +
	( 16'sd 24987) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_139[7:0]) +
	( 14'sd 6688) * $signed(input_fmap_140[7:0]) +
	( 16'sd 28749) * $signed(input_fmap_141[7:0]) +
	( 16'sd 18319) * $signed(input_fmap_142[7:0]) +
	( 16'sd 30090) * $signed(input_fmap_143[7:0]) +
	( 15'sd 10067) * $signed(input_fmap_144[7:0]) +
	( 12'sd 1998) * $signed(input_fmap_145[7:0]) +
	( 15'sd 12150) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3636) * $signed(input_fmap_147[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17176) * $signed(input_fmap_149[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3494) * $signed(input_fmap_151[7:0]) +
	( 14'sd 8144) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2613) * $signed(input_fmap_153[7:0]) +
	( 16'sd 28330) * $signed(input_fmap_154[7:0]) +
	( 16'sd 18238) * $signed(input_fmap_155[7:0]) +
	( 16'sd 16441) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18386) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28995) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5887) * $signed(input_fmap_159[7:0]) +
	( 14'sd 4456) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22854) * $signed(input_fmap_161[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32441) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1722) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30319) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13550) * $signed(input_fmap_166[7:0]) +
	( 16'sd 25482) * $signed(input_fmap_167[7:0]) +
	( 15'sd 11786) * $signed(input_fmap_168[7:0]) +
	( 13'sd 2970) * $signed(input_fmap_169[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19146) * $signed(input_fmap_171[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18730) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16568) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25327) * $signed(input_fmap_175[7:0]) +
	( 15'sd 12963) * $signed(input_fmap_176[7:0]) +
	( 16'sd 26355) * $signed(input_fmap_177[7:0]) +
	( 16'sd 20693) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_179[7:0]) +
	( 16'sd 19196) * $signed(input_fmap_180[7:0]) +
	( 14'sd 4497) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19777) * $signed(input_fmap_182[7:0]) +
	( 12'sd 1755) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26869) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3550) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4779) * $signed(input_fmap_186[7:0]) +
	( 16'sd 26282) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4187) * $signed(input_fmap_188[7:0]) +
	( 16'sd 18418) * $signed(input_fmap_189[7:0]) +
	( 15'sd 11321) * $signed(input_fmap_190[7:0]) +
	( 16'sd 16853) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22616) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5821) * $signed(input_fmap_193[7:0]) +
	( 16'sd 32527) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19525) * $signed(input_fmap_195[7:0]) +
	( 16'sd 23617) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14124) * $signed(input_fmap_197[7:0]) +
	( 15'sd 14621) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15523) * $signed(input_fmap_200[7:0]) +
	( 11'sd 783) * $signed(input_fmap_201[7:0]) +
	( 9'sd 169) * $signed(input_fmap_202[7:0]) +
	( 16'sd 31489) * $signed(input_fmap_203[7:0]) +
	( 16'sd 23768) * $signed(input_fmap_204[7:0]) +
	( 14'sd 7145) * $signed(input_fmap_205[7:0]) +
	( 15'sd 10798) * $signed(input_fmap_206[7:0]) +
	( 16'sd 31177) * $signed(input_fmap_207[7:0]) +
	( 16'sd 27413) * $signed(input_fmap_208[7:0]) +
	( 15'sd 16177) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31141) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30708) * $signed(input_fmap_211[7:0]) +
	( 16'sd 25915) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6444) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7249) * $signed(input_fmap_214[7:0]) +
	( 16'sd 26388) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19869) * $signed(input_fmap_216[7:0]) +
	( 15'sd 12977) * $signed(input_fmap_217[7:0]) +
	( 14'sd 8105) * $signed(input_fmap_218[7:0]) +
	( 14'sd 6186) * $signed(input_fmap_219[7:0]) +
	( 15'sd 9395) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5648) * $signed(input_fmap_221[7:0]) +
	( 16'sd 31993) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14225) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30922) * $signed(input_fmap_224[7:0]) +
	( 11'sd 834) * $signed(input_fmap_225[7:0]) +
	( 16'sd 24866) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19387) * $signed(input_fmap_228[7:0]) +
	( 16'sd 30497) * $signed(input_fmap_229[7:0]) +
	( 16'sd 19847) * $signed(input_fmap_230[7:0]) +
	( 16'sd 30985) * $signed(input_fmap_231[7:0]) +
	( 16'sd 17541) * $signed(input_fmap_232[7:0]) +
	( 15'sd 12012) * $signed(input_fmap_233[7:0]) +
	( 16'sd 20935) * $signed(input_fmap_234[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_235[7:0]) +
	( 12'sd 1300) * $signed(input_fmap_236[7:0]) +
	( 16'sd 16445) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17020) * $signed(input_fmap_238[7:0]) +
	( 12'sd 1995) * $signed(input_fmap_239[7:0]) +
	( 11'sd 752) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30439) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26487) * $signed(input_fmap_242[7:0]) +
	( 16'sd 27494) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13584) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12347) * $signed(input_fmap_245[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_246[7:0]) +
	( 14'sd 6941) * $signed(input_fmap_247[7:0]) +
	( 16'sd 19316) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14225) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26014) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2243) * $signed(input_fmap_251[7:0]) +
	( 12'sd 1873) * $signed(input_fmap_252[7:0]) +
	( 15'sd 14499) * $signed(input_fmap_253[7:0]) +
	( 16'sd 18377) * $signed(input_fmap_254[7:0]) +
	( 13'sd 3590) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_13;
assign conv_mac_13 = 
	( 14'sd 4236) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24969) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28876) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25054) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18622) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7092) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29975) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7936) * $signed(input_fmap_8[7:0]) +
	( 14'sd 8187) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13044) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9372) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25128) * $signed(input_fmap_12[7:0]) +
	( 11'sd 820) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15991) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13457) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21292) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30535) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26560) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27553) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19756) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1880) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15342) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21558) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9857) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12348) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30080) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14644) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14348) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4592) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26951) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14768) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13497) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20907) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15597) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28303) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30197) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11497) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3867) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19900) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19821) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13491) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17906) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32098) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6371) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23197) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16457) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5028) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31727) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23290) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1276) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20075) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3356) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4247) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21459) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27526) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28969) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25126) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10515) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30289) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2332) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14777) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11345) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29184) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3722) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9387) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9841) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30103) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2915) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17117) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7309) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8704) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29521) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27730) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4871) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27175) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5260) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29553) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27226) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19200) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20537) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10373) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21653) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9930) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1589) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3993) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7100) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12447) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23209) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16879) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13364) * $signed(input_fmap_101[7:0]) +
	( 14'sd 8159) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22483) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12877) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16896) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25109) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8571) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7623) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21900) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1035) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12320) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27039) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10683) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24478) * $signed(input_fmap_114[7:0]) +
	( 10'sd 471) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17106) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5833) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15675) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9150) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23266) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10491) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13022) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3434) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29359) * $signed(input_fmap_127[7:0]) +
	( 16'sd 32470) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14303) * $signed(input_fmap_129[7:0]) +
	( 14'sd 4442) * $signed(input_fmap_130[7:0]) +
	( 15'sd 16246) * $signed(input_fmap_131[7:0]) +
	( 16'sd 24965) * $signed(input_fmap_132[7:0]) +
	( 16'sd 27343) * $signed(input_fmap_133[7:0]) +
	( 16'sd 26322) * $signed(input_fmap_134[7:0]) +
	( 12'sd 1096) * $signed(input_fmap_135[7:0]) +
	( 15'sd 9988) * $signed(input_fmap_136[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_137[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2241) * $signed(input_fmap_139[7:0]) +
	( 13'sd 2355) * $signed(input_fmap_140[7:0]) +
	( 16'sd 27633) * $signed(input_fmap_141[7:0]) +
	( 14'sd 7109) * $signed(input_fmap_142[7:0]) +
	( 15'sd 11852) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2483) * $signed(input_fmap_144[7:0]) +
	( 15'sd 14304) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7014) * $signed(input_fmap_146[7:0]) +
	( 16'sd 23949) * $signed(input_fmap_147[7:0]) +
	( 16'sd 32653) * $signed(input_fmap_148[7:0]) +
	( 15'sd 16017) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21687) * $signed(input_fmap_150[7:0]) +
	( 9'sd 195) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7672) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31849) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10209) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27742) * $signed(input_fmap_155[7:0]) +
	( 16'sd 19167) * $signed(input_fmap_156[7:0]) +
	( 15'sd 12651) * $signed(input_fmap_157[7:0]) +
	( 13'sd 3850) * $signed(input_fmap_158[7:0]) +
	( 16'sd 19575) * $signed(input_fmap_159[7:0]) +
	( 15'sd 8429) * $signed(input_fmap_160[7:0]) +
	( 15'sd 14700) * $signed(input_fmap_161[7:0]) +
	( 16'sd 20335) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_163[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_164[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30316) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20915) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26410) * $signed(input_fmap_168[7:0]) +
	( 15'sd 9590) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11695) * $signed(input_fmap_170[7:0]) +
	( 16'sd 17730) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7582) * $signed(input_fmap_172[7:0]) +
	( 14'sd 6596) * $signed(input_fmap_173[7:0]) +
	( 14'sd 4855) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3358) * $signed(input_fmap_175[7:0]) +
	( 15'sd 9230) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18031) * $signed(input_fmap_177[7:0]) +
	( 16'sd 16919) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5064) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15618) * $signed(input_fmap_180[7:0]) +
	( 16'sd 20165) * $signed(input_fmap_181[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_182[7:0]) +
	( 15'sd 13557) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8216) * $signed(input_fmap_184[7:0]) +
	( 11'sd 819) * $signed(input_fmap_185[7:0]) +
	( 16'sd 24281) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22129) * $signed(input_fmap_187[7:0]) +
	( 16'sd 19956) * $signed(input_fmap_188[7:0]) +
	( 16'sd 21031) * $signed(input_fmap_189[7:0]) +
	( 10'sd 349) * $signed(input_fmap_190[7:0]) +
	( 16'sd 27424) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20028) * $signed(input_fmap_193[7:0]) +
	( 16'sd 25582) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19916) * $signed(input_fmap_195[7:0]) +
	( 16'sd 18680) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31436) * $signed(input_fmap_197[7:0]) +
	( 15'sd 15331) * $signed(input_fmap_198[7:0]) +
	( 16'sd 32182) * $signed(input_fmap_199[7:0]) +
	( 16'sd 17667) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3092) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5268) * $signed(input_fmap_202[7:0]) +
	( 15'sd 10704) * $signed(input_fmap_203[7:0]) +
	( 16'sd 31009) * $signed(input_fmap_204[7:0]) +
	( 15'sd 8503) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21062) * $signed(input_fmap_206[7:0]) +
	( 16'sd 24036) * $signed(input_fmap_207[7:0]) +
	( 15'sd 14597) * $signed(input_fmap_208[7:0]) +
	( 16'sd 27260) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5244) * $signed(input_fmap_211[7:0]) +
	( 14'sd 5425) * $signed(input_fmap_212[7:0]) +
	( 16'sd 17051) * $signed(input_fmap_213[7:0]) +
	( 16'sd 32549) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23485) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24718) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24550) * $signed(input_fmap_217[7:0]) +
	( 16'sd 25373) * $signed(input_fmap_218[7:0]) +
	( 16'sd 32280) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19692) * $signed(input_fmap_220[7:0]) +
	( 16'sd 18551) * $signed(input_fmap_221[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_222[7:0]) +
	( 15'sd 16051) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19915) * $signed(input_fmap_224[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30697) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6353) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6141) * $signed(input_fmap_229[7:0]) +
	( 15'sd 8724) * $signed(input_fmap_230[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_231[7:0]) +
	( 11'sd 561) * $signed(input_fmap_232[7:0]) +
	( 16'sd 16751) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3099) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26543) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10100) * $signed(input_fmap_236[7:0]) +
	( 16'sd 23664) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16721) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20874) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10156) * $signed(input_fmap_240[7:0]) +
	( 14'sd 4304) * $signed(input_fmap_241[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_243[7:0]) +
	( 16'sd 23604) * $signed(input_fmap_244[7:0]) +
	( 15'sd 9735) * $signed(input_fmap_245[7:0]) +
	( 16'sd 25357) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12549) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26137) * $signed(input_fmap_248[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7037) * $signed(input_fmap_250[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_251[7:0]) +
	( 16'sd 31826) * $signed(input_fmap_252[7:0]) +
	( 15'sd 12135) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1417) * $signed(input_fmap_254[7:0]) +
	( 16'sd 28986) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_14;
assign conv_mac_14 = 
	( 15'sd 10686) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6034) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1728) * $signed(input_fmap_3[7:0]) +
	( 11'sd 759) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4953) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1872) * $signed(input_fmap_6[7:0]) +
	( 10'sd 458) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27534) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28301) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3975) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28668) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32480) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16807) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18164) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14360) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20349) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2656) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23876) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15825) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6898) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14420) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22699) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23380) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26761) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20456) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28262) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9025) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23021) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4727) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22706) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25687) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10095) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1836) * $signed(input_fmap_40[7:0]) +
	( 12'sd 2010) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23573) * $signed(input_fmap_42[7:0]) +
	( 11'sd 644) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13654) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25154) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12948) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13091) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12246) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7111) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4161) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29390) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12221) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31284) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31993) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1983) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26510) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1529) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23495) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31597) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12817) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26725) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1464) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31444) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23114) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29181) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24019) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9036) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9884) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17112) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21571) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9806) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14111) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7411) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16521) * $signed(input_fmap_78[7:0]) +
	( 11'sd 549) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22267) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26854) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2446) * $signed(input_fmap_82[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29481) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24588) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13545) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16103) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21063) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6163) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29324) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28604) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26764) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31514) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18053) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21096) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7962) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14979) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31627) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26172) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23800) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26366) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5981) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9245) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13958) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11479) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30725) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4919) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7011) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7087) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6471) * $signed(input_fmap_112[7:0]) +
	( 9'sd 194) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9428) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6879) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15390) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15377) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17576) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32018) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1441) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17273) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16452) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4195) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29001) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3676) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16043) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9243) * $signed(input_fmap_128[7:0]) +
	( 16'sd 22309) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_130[7:0]) +
	( 16'sd 28628) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18444) * $signed(input_fmap_132[7:0]) +
	( 16'sd 24867) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32331) * $signed(input_fmap_134[7:0]) +
	( 13'sd 3299) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15154) * $signed(input_fmap_136[7:0]) +
	( 16'sd 16731) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11918) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21216) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_140[7:0]) +
	( 16'sd 16818) * $signed(input_fmap_141[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20582) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_144[7:0]) +
	( 16'sd 30939) * $signed(input_fmap_145[7:0]) +
	( 16'sd 20757) * $signed(input_fmap_146[7:0]) +
	( 15'sd 15307) * $signed(input_fmap_147[7:0]) +
	( 15'sd 9681) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27179) * $signed(input_fmap_149[7:0]) +
	( 12'sd 1352) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19793) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2542) * $signed(input_fmap_152[7:0]) +
	( 14'sd 6538) * $signed(input_fmap_153[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13462) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25241) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20469) * $signed(input_fmap_157[7:0]) +
	( 15'sd 14813) * $signed(input_fmap_158[7:0]) +
	( 16'sd 31164) * $signed(input_fmap_159[7:0]) +
	( 15'sd 12333) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19559) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30744) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3707) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28761) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9261) * $signed(input_fmap_166[7:0]) +
	( 14'sd 4196) * $signed(input_fmap_167[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27343) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18371) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15605) * $signed(input_fmap_172[7:0]) +
	( 14'sd 4303) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11857) * $signed(input_fmap_174[7:0]) +
	( 16'sd 19873) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29909) * $signed(input_fmap_176[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32001) * $signed(input_fmap_178[7:0]) +
	( 8'sd 78) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21526) * $signed(input_fmap_180[7:0]) +
	( 16'sd 20415) * $signed(input_fmap_181[7:0]) +
	( 16'sd 28133) * $signed(input_fmap_182[7:0]) +
	( 14'sd 7297) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9574) * $signed(input_fmap_184[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_185[7:0]) +
	( 16'sd 27780) * $signed(input_fmap_186[7:0]) +
	( 15'sd 15095) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1999) * $signed(input_fmap_188[7:0]) +
	( 16'sd 29462) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28431) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24024) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28353) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27882) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17405) * $signed(input_fmap_196[7:0]) +
	( 14'sd 4993) * $signed(input_fmap_197[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20989) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18503) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13682) * $signed(input_fmap_201[7:0]) +
	( 14'sd 6249) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13169) * $signed(input_fmap_203[7:0]) +
	( 16'sd 31290) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6168) * $signed(input_fmap_205[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_206[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17411) * $signed(input_fmap_208[7:0]) +
	( 14'sd 6921) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11493) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28480) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26368) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1203) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17924) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23778) * $signed(input_fmap_215[7:0]) +
	( 15'sd 15222) * $signed(input_fmap_216[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_217[7:0]) +
	( 13'sd 3575) * $signed(input_fmap_218[7:0]) +
	( 14'sd 8181) * $signed(input_fmap_219[7:0]) +
	( 14'sd 6884) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1718) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10089) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19703) * $signed(input_fmap_224[7:0]) +
	( 14'sd 7735) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29604) * $signed(input_fmap_226[7:0]) +
	( 16'sd 21693) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24572) * $signed(input_fmap_228[7:0]) +
	( 16'sd 32042) * $signed(input_fmap_229[7:0]) +
	( 15'sd 11071) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3718) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18530) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11267) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18815) * $signed(input_fmap_234[7:0]) +
	( 13'sd 2311) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27488) * $signed(input_fmap_236[7:0]) +
	( 16'sd 22594) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22797) * $signed(input_fmap_238[7:0]) +
	( 16'sd 24139) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1269) * $signed(input_fmap_240[7:0]) +
	( 16'sd 16911) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26916) * $signed(input_fmap_242[7:0]) +
	( 16'sd 30648) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28470) * $signed(input_fmap_244[7:0]) +
	( 16'sd 17075) * $signed(input_fmap_245[7:0]) +
	( 14'sd 4272) * $signed(input_fmap_246[7:0]) +
	( 15'sd 16374) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32595) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12978) * $signed(input_fmap_249[7:0]) +
	( 14'sd 4199) * $signed(input_fmap_250[7:0]) +
	( 15'sd 9242) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26982) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27766) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1534) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10702) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_15;
assign conv_mac_15 = 
	( 11'sd 561) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11397) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10357) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16460) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28223) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12421) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11157) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27641) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18401) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6862) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26542) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14842) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30306) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19297) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30131) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1202) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3906) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4221) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26493) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20371) * $signed(input_fmap_23[7:0]) +
	( 8'sd 72) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26519) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9369) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15487) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13387) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25139) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20846) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29577) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19790) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2806) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3030) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32687) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9689) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1226) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17575) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3491) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9545) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20825) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26963) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22116) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1653) * $signed(input_fmap_48[7:0]) +
	( 12'sd 2008) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7081) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18486) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21104) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28626) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27399) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21699) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25014) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26892) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16242) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19801) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10180) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8332) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17667) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13703) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20113) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6389) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28407) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1932) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12611) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8680) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26589) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5732) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32282) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15477) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31315) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1958) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15861) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20666) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16253) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20096) * $signed(input_fmap_86[7:0]) +
	( 11'sd 542) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2815) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26534) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14621) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21376) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27939) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17699) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20722) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31198) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16075) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4593) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10140) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25088) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13497) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27915) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4746) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20547) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11967) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22670) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24705) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29304) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17224) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21368) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26841) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13670) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1959) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11329) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20866) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22523) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8235) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16545) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20380) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22681) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30049) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1273) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11121) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12716) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8146) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29080) * $signed(input_fmap_128[7:0]) +
	( 15'sd 11319) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6375) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20525) * $signed(input_fmap_131[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_132[7:0]) +
	( 10'sd 403) * $signed(input_fmap_133[7:0]) +
	( 16'sd 20564) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18682) * $signed(input_fmap_135[7:0]) +
	( 16'sd 29530) * $signed(input_fmap_136[7:0]) +
	( 15'sd 16146) * $signed(input_fmap_137[7:0]) +
	( 14'sd 4743) * $signed(input_fmap_138[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_139[7:0]) +
	( 15'sd 16199) * $signed(input_fmap_140[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21316) * $signed(input_fmap_142[7:0]) +
	( 15'sd 11627) * $signed(input_fmap_143[7:0]) +
	( 16'sd 25888) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25071) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27075) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24866) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21872) * $signed(input_fmap_148[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_149[7:0]) +
	( 16'sd 32717) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6378) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31889) * $signed(input_fmap_152[7:0]) +
	( 14'sd 5979) * $signed(input_fmap_153[7:0]) +
	( 16'sd 29989) * $signed(input_fmap_154[7:0]) +
	( 16'sd 21640) * $signed(input_fmap_155[7:0]) +
	( 16'sd 27235) * $signed(input_fmap_156[7:0]) +
	( 13'sd 2518) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9934) * $signed(input_fmap_158[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27808) * $signed(input_fmap_160[7:0]) +
	( 15'sd 15454) * $signed(input_fmap_161[7:0]) +
	( 16'sd 28565) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24330) * $signed(input_fmap_163[7:0]) +
	( 16'sd 23845) * $signed(input_fmap_164[7:0]) +
	( 14'sd 6002) * $signed(input_fmap_165[7:0]) +
	( 16'sd 27334) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30579) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4807) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3484) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23927) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11452) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_172[7:0]) +
	( 10'sd 401) * $signed(input_fmap_173[7:0]) +
	( 15'sd 13126) * $signed(input_fmap_174[7:0]) +
	( 13'sd 2851) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27157) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24262) * $signed(input_fmap_177[7:0]) +
	( 11'sd 742) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15629) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4449) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25482) * $signed(input_fmap_181[7:0]) +
	( 12'sd 1043) * $signed(input_fmap_182[7:0]) +
	( 15'sd 14048) * $signed(input_fmap_183[7:0]) +
	( 15'sd 12080) * $signed(input_fmap_184[7:0]) +
	( 11'sd 619) * $signed(input_fmap_185[7:0]) +
	( 15'sd 14517) * $signed(input_fmap_186[7:0]) +
	( 14'sd 7012) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4754) * $signed(input_fmap_188[7:0]) +
	( 14'sd 4164) * $signed(input_fmap_189[7:0]) +
	( 13'sd 4077) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31613) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29560) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27057) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29307) * $signed(input_fmap_194[7:0]) +
	( 16'sd 31733) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15834) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11958) * $signed(input_fmap_197[7:0]) +
	( 16'sd 16821) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12818) * $signed(input_fmap_199[7:0]) +
	( 16'sd 27832) * $signed(input_fmap_200[7:0]) +
	( 13'sd 2621) * $signed(input_fmap_201[7:0]) +
	( 14'sd 6968) * $signed(input_fmap_202[7:0]) +
	( 15'sd 9191) * $signed(input_fmap_203[7:0]) +
	( 15'sd 8653) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30964) * $signed(input_fmap_205[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13323) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25666) * $signed(input_fmap_208[7:0]) +
	( 14'sd 6019) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19221) * $signed(input_fmap_210[7:0]) +
	( 16'sd 22920) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29549) * $signed(input_fmap_212[7:0]) +
	( 16'sd 19050) * $signed(input_fmap_213[7:0]) +
	( 16'sd 25553) * $signed(input_fmap_214[7:0]) +
	( 16'sd 19722) * $signed(input_fmap_215[7:0]) +
	( 16'sd 27691) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24454) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13899) * $signed(input_fmap_218[7:0]) +
	( 16'sd 31651) * $signed(input_fmap_219[7:0]) +
	( 11'sd 527) * $signed(input_fmap_220[7:0]) +
	( 16'sd 24982) * $signed(input_fmap_221[7:0]) +
	( 16'sd 16721) * $signed(input_fmap_222[7:0]) +
	( 12'sd 1318) * $signed(input_fmap_223[7:0]) +
	( 15'sd 10774) * $signed(input_fmap_224[7:0]) +
	( 15'sd 11443) * $signed(input_fmap_225[7:0]) +
	( 15'sd 9814) * $signed(input_fmap_226[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_227[7:0]) +
	( 16'sd 20687) * $signed(input_fmap_228[7:0]) +
	( 15'sd 11960) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7978) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20021) * $signed(input_fmap_232[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_234[7:0]) +
	( 16'sd 23084) * $signed(input_fmap_235[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_236[7:0]) +
	( 16'sd 23874) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23779) * $signed(input_fmap_238[7:0]) +
	( 16'sd 27447) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18520) * $signed(input_fmap_240[7:0]) +
	( 16'sd 24172) * $signed(input_fmap_241[7:0]) +
	( 8'sd 93) * $signed(input_fmap_242[7:0]) +
	( 16'sd 30738) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12124) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10031) * $signed(input_fmap_245[7:0]) +
	( 13'sd 3507) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3432) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28669) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12387) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12325) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17093) * $signed(input_fmap_252[7:0]) +
	( 16'sd 18906) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31431) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5706) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_16;
assign conv_mac_16 = 
	( 16'sd 16476) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5251) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24585) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29487) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12258) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8548) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5086) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14389) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11717) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25810) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30377) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9317) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16982) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3627) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3963) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31756) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21453) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2613) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19915) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14706) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15296) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20679) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18111) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31007) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22977) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23774) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30773) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28479) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21349) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7628) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7237) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7142) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9903) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24278) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4148) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31275) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6203) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22413) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30805) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16143) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28836) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8493) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31329) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7949) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13642) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17720) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14207) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1061) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19146) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19093) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11146) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28823) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4723) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6617) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17703) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19570) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12981) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14332) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17765) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7395) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21809) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30570) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24451) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30026) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4727) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9236) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6521) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1058) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29321) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22175) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12850) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3367) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11738) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20932) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1682) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32746) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18283) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7284) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28473) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7496) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24254) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4836) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18875) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1565) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2150) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8774) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31422) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23930) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23068) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29682) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20971) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28464) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23118) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11594) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9665) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24193) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14539) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24127) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2986) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2636) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12773) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18991) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10433) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9364) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17923) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12561) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4974) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17164) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1186) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15495) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15199) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4256) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_127[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_128[7:0]) +
	( 15'sd 11142) * $signed(input_fmap_129[7:0]) +
	( 14'sd 4173) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5959) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14443) * $signed(input_fmap_132[7:0]) +
	( 16'sd 24655) * $signed(input_fmap_133[7:0]) +
	( 16'sd 30028) * $signed(input_fmap_134[7:0]) +
	( 14'sd 5416) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8977) * $signed(input_fmap_136[7:0]) +
	( 16'sd 21124) * $signed(input_fmap_137[7:0]) +
	( 15'sd 13767) * $signed(input_fmap_138[7:0]) +
	( 16'sd 22231) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19112) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31734) * $signed(input_fmap_143[7:0]) +
	( 16'sd 25863) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23541) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9743) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19770) * $signed(input_fmap_147[7:0]) +
	( 15'sd 8814) * $signed(input_fmap_148[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_149[7:0]) +
	( 16'sd 19208) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18651) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16389) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_153[7:0]) +
	( 16'sd 29492) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15325) * $signed(input_fmap_156[7:0]) +
	( 13'sd 3745) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25760) * $signed(input_fmap_158[7:0]) +
	( 11'sd 809) * $signed(input_fmap_159[7:0]) +
	( 16'sd 28162) * $signed(input_fmap_160[7:0]) +
	( 16'sd 18278) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13644) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32237) * $signed(input_fmap_163[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9230) * $signed(input_fmap_165[7:0]) +
	( 16'sd 25923) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23059) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1790) * $signed(input_fmap_168[7:0]) +
	( 16'sd 24246) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24787) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30061) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9470) * $signed(input_fmap_172[7:0]) +
	( 16'sd 22783) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19117) * $signed(input_fmap_174[7:0]) +
	( 16'sd 22605) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1881) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19587) * $signed(input_fmap_177[7:0]) +
	( 16'sd 19249) * $signed(input_fmap_178[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6328) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30676) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_182[7:0]) +
	( 10'sd 338) * $signed(input_fmap_183[7:0]) +
	( 16'sd 28622) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27875) * $signed(input_fmap_185[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11710) * $signed(input_fmap_187[7:0]) +
	( 11'sd 757) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3727) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17788) * $signed(input_fmap_191[7:0]) +
	( 16'sd 30184) * $signed(input_fmap_192[7:0]) +
	( 14'sd 4880) * $signed(input_fmap_193[7:0]) +
	( 14'sd 6141) * $signed(input_fmap_194[7:0]) +
	( 15'sd 10799) * $signed(input_fmap_195[7:0]) +
	( 16'sd 26657) * $signed(input_fmap_196[7:0]) +
	( 16'sd 27167) * $signed(input_fmap_197[7:0]) +
	( 16'sd 23644) * $signed(input_fmap_198[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_200[7:0]) +
	( 16'sd 28569) * $signed(input_fmap_201[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19539) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_204[7:0]) +
	( 16'sd 22364) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29417) * $signed(input_fmap_206[7:0]) +
	( 15'sd 10278) * $signed(input_fmap_207[7:0]) +
	( 16'sd 29292) * $signed(input_fmap_208[7:0]) +
	( 11'sd 667) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4788) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23205) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17814) * $signed(input_fmap_212[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30897) * $signed(input_fmap_214[7:0]) +
	( 16'sd 32548) * $signed(input_fmap_215[7:0]) +
	( 15'sd 9971) * $signed(input_fmap_216[7:0]) +
	( 16'sd 27831) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31727) * $signed(input_fmap_218[7:0]) +
	( 15'sd 13148) * $signed(input_fmap_219[7:0]) +
	( 14'sd 5202) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6312) * $signed(input_fmap_221[7:0]) +
	( 16'sd 20817) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17647) * $signed(input_fmap_223[7:0]) +
	( 14'sd 5533) * $signed(input_fmap_224[7:0]) +
	( 16'sd 16395) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14772) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3388) * $signed(input_fmap_227[7:0]) +
	( 16'sd 28944) * $signed(input_fmap_228[7:0]) +
	( 16'sd 31002) * $signed(input_fmap_229[7:0]) +
	( 16'sd 20331) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13811) * $signed(input_fmap_231[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3170) * $signed(input_fmap_233[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_234[7:0]) +
	( 16'sd 28411) * $signed(input_fmap_235[7:0]) +
	( 15'sd 8694) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11328) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12911) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19397) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25412) * $signed(input_fmap_240[7:0]) +
	( 16'sd 24105) * $signed(input_fmap_241[7:0]) +
	( 16'sd 24868) * $signed(input_fmap_242[7:0]) +
	( 11'sd 741) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24453) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10902) * $signed(input_fmap_246[7:0]) +
	( 14'sd 5349) * $signed(input_fmap_247[7:0]) +
	( 15'sd 11378) * $signed(input_fmap_248[7:0]) +
	( 14'sd 7754) * $signed(input_fmap_249[7:0]) +
	( 15'sd 15503) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27676) * $signed(input_fmap_251[7:0]) +
	( 16'sd 19515) * $signed(input_fmap_252[7:0]) +
	( 16'sd 18774) * $signed(input_fmap_253[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_254[7:0]) +
	( 13'sd 3669) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_17;
assign conv_mac_17 = 
	( 15'sd 9112) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31697) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32062) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25557) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28507) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14092) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3077) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13563) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28450) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4170) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17570) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26283) * $signed(input_fmap_14[7:0]) +
	( 11'sd 893) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20372) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18216) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31816) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17340) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1674) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23792) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2511) * $signed(input_fmap_22[7:0]) +
	( 11'sd 685) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23002) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15636) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24954) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14977) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9892) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19983) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3798) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15589) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22383) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5586) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1040) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13493) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3606) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17309) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29258) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21203) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23224) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31363) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31069) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17080) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22070) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8918) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14190) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14009) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6350) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11725) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12500) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5788) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20688) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12478) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26743) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28691) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12396) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18985) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20685) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7245) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19437) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28199) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4258) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20231) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13381) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13052) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5512) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21103) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16429) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8421) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6138) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28393) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20111) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31970) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23119) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31268) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20160) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27301) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13196) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28492) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13300) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7665) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16252) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2181) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12358) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12592) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30708) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27519) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3377) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25821) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30054) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19114) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18461) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24960) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16851) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29500) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13261) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14658) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4218) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23068) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8551) * $signed(input_fmap_106[7:0]) +
	( 9'sd 242) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21439) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31337) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15792) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25261) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17781) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28600) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20319) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17797) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22235) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10070) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21213) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7396) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6947) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22275) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27207) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17638) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20585) * $signed(input_fmap_127[7:0]) +
	( 16'sd 24109) * $signed(input_fmap_128[7:0]) +
	( 16'sd 29154) * $signed(input_fmap_129[7:0]) +
	( 11'sd 864) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24622) * $signed(input_fmap_131[7:0]) +
	( 16'sd 27770) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10536) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1309) * $signed(input_fmap_134[7:0]) +
	( 14'sd 6471) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2717) * $signed(input_fmap_136[7:0]) +
	( 16'sd 28487) * $signed(input_fmap_137[7:0]) +
	( 14'sd 6284) * $signed(input_fmap_138[7:0]) +
	( 12'sd 1340) * $signed(input_fmap_139[7:0]) +
	( 11'sd 942) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3797) * $signed(input_fmap_141[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_142[7:0]) +
	( 15'sd 14800) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4592) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23505) * $signed(input_fmap_145[7:0]) +
	( 16'sd 30023) * $signed(input_fmap_146[7:0]) +
	( 10'sd 494) * $signed(input_fmap_147[7:0]) +
	( 16'sd 19144) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4768) * $signed(input_fmap_149[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_150[7:0]) +
	( 16'sd 27988) * $signed(input_fmap_151[7:0]) +
	( 15'sd 15526) * $signed(input_fmap_152[7:0]) +
	( 16'sd 16405) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25839) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_155[7:0]) +
	( 15'sd 11930) * $signed(input_fmap_156[7:0]) +
	( 14'sd 4770) * $signed(input_fmap_157[7:0]) +
	( 10'sd 291) * $signed(input_fmap_158[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_159[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_160[7:0]) +
	( 16'sd 21428) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10571) * $signed(input_fmap_162[7:0]) +
	( 16'sd 16948) * $signed(input_fmap_163[7:0]) +
	( 15'sd 15613) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22761) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31118) * $signed(input_fmap_166[7:0]) +
	( 16'sd 16440) * $signed(input_fmap_167[7:0]) +
	( 16'sd 21949) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30838) * $signed(input_fmap_169[7:0]) +
	( 15'sd 15143) * $signed(input_fmap_170[7:0]) +
	( 16'sd 28547) * $signed(input_fmap_171[7:0]) +
	( 15'sd 8232) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27522) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27406) * $signed(input_fmap_174[7:0]) +
	( 15'sd 12447) * $signed(input_fmap_175[7:0]) +
	( 15'sd 8814) * $signed(input_fmap_176[7:0]) +
	( 15'sd 14150) * $signed(input_fmap_177[7:0]) +
	( 14'sd 4990) * $signed(input_fmap_178[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11045) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4130) * $signed(input_fmap_182[7:0]) +
	( 15'sd 16099) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13967) * $signed(input_fmap_184[7:0]) +
	( 13'sd 2551) * $signed(input_fmap_185[7:0]) +
	( 16'sd 20646) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25557) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12858) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19514) * $signed(input_fmap_189[7:0]) +
	( 14'sd 7433) * $signed(input_fmap_190[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_191[7:0]) +
	( 15'sd 8462) * $signed(input_fmap_192[7:0]) +
	( 16'sd 18728) * $signed(input_fmap_193[7:0]) +
	( 16'sd 19266) * $signed(input_fmap_194[7:0]) +
	( 9'sd 236) * $signed(input_fmap_195[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32469) * $signed(input_fmap_197[7:0]) +
	( 14'sd 4723) * $signed(input_fmap_198[7:0]) +
	( 16'sd 17773) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_200[7:0]) +
	( 16'sd 19915) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8951) * $signed(input_fmap_202[7:0]) +
	( 15'sd 14294) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15907) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28814) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12483) * $signed(input_fmap_206[7:0]) +
	( 10'sd 258) * $signed(input_fmap_207[7:0]) +
	( 16'sd 19829) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23718) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30695) * $signed(input_fmap_210[7:0]) +
	( 15'sd 13075) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24924) * $signed(input_fmap_212[7:0]) +
	( 14'sd 8085) * $signed(input_fmap_213[7:0]) +
	( 16'sd 27290) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5017) * $signed(input_fmap_215[7:0]) +
	( 16'sd 31436) * $signed(input_fmap_216[7:0]) +
	( 15'sd 8481) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_218[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13284) * $signed(input_fmap_220[7:0]) +
	( 16'sd 32275) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19273) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8753) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1035) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13252) * $signed(input_fmap_225[7:0]) +
	( 15'sd 12198) * $signed(input_fmap_226[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_227[7:0]) +
	( 13'sd 3188) * $signed(input_fmap_228[7:0]) +
	( 12'sd 1505) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7886) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28521) * $signed(input_fmap_231[7:0]) +
	( 16'sd 32152) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11204) * $signed(input_fmap_233[7:0]) +
	( 16'sd 32096) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3840) * $signed(input_fmap_235[7:0]) +
	( 15'sd 16054) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2531) * $signed(input_fmap_237[7:0]) +
	( 16'sd 24339) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9055) * $signed(input_fmap_239[7:0]) +
	( 13'sd 2841) * $signed(input_fmap_240[7:0]) +
	( 12'sd 1922) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29184) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28239) * $signed(input_fmap_243[7:0]) +
	( 15'sd 11074) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12417) * $signed(input_fmap_245[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_246[7:0]) +
	( 14'sd 6271) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10364) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4882) * $signed(input_fmap_249[7:0]) +
	( 16'sd 21802) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19548) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4541) * $signed(input_fmap_252[7:0]) +
	( 16'sd 30196) * $signed(input_fmap_253[7:0]) +
	( 14'sd 6326) * $signed(input_fmap_254[7:0]) +
	( 16'sd 17966) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_18;
assign conv_mac_18 = 
	( 16'sd 26362) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6774) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_2[7:0]) +
	( 14'sd 8033) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24855) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3901) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7906) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18649) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15530) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28135) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30312) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2457) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7154) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7104) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4730) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16730) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8868) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11169) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2359) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24886) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22356) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11529) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17363) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17290) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27257) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14133) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29224) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9385) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27879) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25430) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29482) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24330) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24318) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20729) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26607) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22551) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8989) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23393) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26753) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8195) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2201) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13202) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12103) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6867) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11532) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20238) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8944) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21621) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8511) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31185) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8631) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23267) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1996) * $signed(input_fmap_59[7:0]) +
	( 10'sd 365) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29589) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15938) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19176) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30962) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19103) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16674) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31097) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6983) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7989) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7714) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3594) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4389) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11513) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18764) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4786) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19501) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31140) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4190) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13546) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30770) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10493) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2475) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18238) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7463) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12651) * $signed(input_fmap_87[7:0]) +
	( 9'sd 255) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9637) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32318) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26526) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2426) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23631) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16771) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21407) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5922) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19246) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23784) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17348) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17521) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25164) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15240) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1625) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12560) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18371) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21205) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4975) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14245) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29063) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22936) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20545) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23015) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24366) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2629) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5229) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9322) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31005) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29546) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9092) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3490) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14173) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9203) * $signed(input_fmap_128[7:0]) +
	( 15'sd 12559) * $signed(input_fmap_129[7:0]) +
	( 15'sd 11158) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23250) * $signed(input_fmap_131[7:0]) +
	( 15'sd 12706) * $signed(input_fmap_132[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19292) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10517) * $signed(input_fmap_135[7:0]) +
	( 16'sd 22219) * $signed(input_fmap_136[7:0]) +
	( 16'sd 16896) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11681) * $signed(input_fmap_138[7:0]) +
	( 12'sd 1918) * $signed(input_fmap_139[7:0]) +
	( 15'sd 13567) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5465) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25122) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23169) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27726) * $signed(input_fmap_145[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9895) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23920) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27818) * $signed(input_fmap_149[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_150[7:0]) +
	( 15'sd 11667) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3267) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24156) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5603) * $signed(input_fmap_155[7:0]) +
	( 16'sd 21907) * $signed(input_fmap_156[7:0]) +
	( 11'sd 1003) * $signed(input_fmap_157[7:0]) +
	( 14'sd 5441) * $signed(input_fmap_158[7:0]) +
	( 15'sd 9239) * $signed(input_fmap_159[7:0]) +
	( 15'sd 12795) * $signed(input_fmap_160[7:0]) +
	( 16'sd 24556) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14735) * $signed(input_fmap_162[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1102) * $signed(input_fmap_164[7:0]) +
	( 16'sd 17310) * $signed(input_fmap_165[7:0]) +
	( 14'sd 5146) * $signed(input_fmap_166[7:0]) +
	( 16'sd 29301) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29031) * $signed(input_fmap_168[7:0]) +
	( 15'sd 8682) * $signed(input_fmap_169[7:0]) +
	( 14'sd 4659) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18548) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7455) * $signed(input_fmap_172[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_173[7:0]) +
	( 15'sd 9796) * $signed(input_fmap_174[7:0]) +
	( 16'sd 23028) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13129) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15792) * $signed(input_fmap_177[7:0]) +
	( 16'sd 24653) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6191) * $signed(input_fmap_179[7:0]) +
	( 16'sd 22308) * $signed(input_fmap_180[7:0]) +
	( 16'sd 31162) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30388) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27810) * $signed(input_fmap_183[7:0]) +
	( 12'sd 1813) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22058) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12086) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4248) * $signed(input_fmap_187[7:0]) +
	( 15'sd 11193) * $signed(input_fmap_188[7:0]) +
	( 16'sd 27405) * $signed(input_fmap_189[7:0]) +
	( 13'sd 2499) * $signed(input_fmap_190[7:0]) +
	( 16'sd 28320) * $signed(input_fmap_191[7:0]) +
	( 15'sd 10602) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22328) * $signed(input_fmap_193[7:0]) +
	( 14'sd 5149) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27250) * $signed(input_fmap_195[7:0]) +
	( 10'sd 417) * $signed(input_fmap_196[7:0]) +
	( 13'sd 3861) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10656) * $signed(input_fmap_199[7:0]) +
	( 15'sd 12748) * $signed(input_fmap_200[7:0]) +
	( 16'sd 23004) * $signed(input_fmap_201[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_202[7:0]) +
	( 14'sd 4686) * $signed(input_fmap_203[7:0]) +
	( 16'sd 22708) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12078) * $signed(input_fmap_205[7:0]) +
	( 15'sd 13829) * $signed(input_fmap_206[7:0]) +
	( 15'sd 16359) * $signed(input_fmap_207[7:0]) +
	( 15'sd 13866) * $signed(input_fmap_208[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_209[7:0]) +
	( 16'sd 16841) * $signed(input_fmap_210[7:0]) +
	( 16'sd 18607) * $signed(input_fmap_211[7:0]) +
	( 15'sd 16028) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12225) * $signed(input_fmap_213[7:0]) +
	( 15'sd 8386) * $signed(input_fmap_214[7:0]) +
	( 16'sd 32684) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18165) * $signed(input_fmap_216[7:0]) +
	( 15'sd 15027) * $signed(input_fmap_217[7:0]) +
	( 15'sd 9372) * $signed(input_fmap_218[7:0]) +
	( 13'sd 2324) * $signed(input_fmap_219[7:0]) +
	( 16'sd 27171) * $signed(input_fmap_220[7:0]) +
	( 15'sd 11353) * $signed(input_fmap_221[7:0]) +
	( 16'sd 17708) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12779) * $signed(input_fmap_223[7:0]) +
	( 16'sd 22555) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3611) * $signed(input_fmap_225[7:0]) +
	( 16'sd 19563) * $signed(input_fmap_226[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10820) * $signed(input_fmap_228[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_229[7:0]) +
	( 12'sd 1660) * $signed(input_fmap_230[7:0]) +
	( 15'sd 11216) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12222) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_233[7:0]) +
	( 16'sd 20597) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11579) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28468) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17584) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6867) * $signed(input_fmap_240[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1859) * $signed(input_fmap_242[7:0]) +
	( 16'sd 27979) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12132) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6623) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31571) * $signed(input_fmap_246[7:0]) +
	( 16'sd 25724) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4255) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3614) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30252) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20907) * $signed(input_fmap_254[7:0]) +
	( 12'sd 1658) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_19;
assign conv_mac_19 = 
	( 16'sd 28995) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28292) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11246) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24391) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15055) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5114) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7106) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26762) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29572) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21032) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19372) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4564) * $signed(input_fmap_14[7:0]) +
	( 11'sd 541) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10198) * $signed(input_fmap_16[7:0]) +
	( 10'sd 288) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30625) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5066) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29255) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24879) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12730) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1882) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11024) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1943) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21305) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27983) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16072) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14245) * $signed(input_fmap_31[7:0]) +
	( 11'sd 924) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13951) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5353) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16799) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2313) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2138) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24457) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18577) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20211) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22685) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22361) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18271) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6783) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22746) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7788) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14784) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5155) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29121) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27142) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25221) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9724) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23879) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3398) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28217) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9263) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16398) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29265) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6994) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18352) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20405) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22864) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19049) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3454) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31087) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3308) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_72[7:0]) +
	( 6'sd 24) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30702) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7593) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13764) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9923) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29519) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28398) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22720) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17469) * $signed(input_fmap_81[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_82[7:0]) +
	( 11'sd 881) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4973) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10376) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3937) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4502) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28601) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31824) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22788) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8971) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31378) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8657) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18040) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26201) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18054) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14173) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6295) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5980) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19445) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23030) * $signed(input_fmap_101[7:0]) +
	( 14'sd 8045) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18121) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28354) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14789) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24146) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4833) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31799) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27788) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21246) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6020) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26317) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10524) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2209) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14725) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6071) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17823) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22945) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27778) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19795) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4819) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13239) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15829) * $signed(input_fmap_128[7:0]) +
	( 16'sd 16854) * $signed(input_fmap_129[7:0]) +
	( 16'sd 21549) * $signed(input_fmap_130[7:0]) +
	( 16'sd 28961) * $signed(input_fmap_131[7:0]) +
	( 16'sd 19768) * $signed(input_fmap_132[7:0]) +
	( 16'sd 17231) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25814) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26635) * $signed(input_fmap_135[7:0]) +
	( 16'sd 16908) * $signed(input_fmap_136[7:0]) +
	( 16'sd 19303) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29495) * $signed(input_fmap_138[7:0]) +
	( 15'sd 10742) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15397) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3080) * $signed(input_fmap_141[7:0]) +
	( 14'sd 5079) * $signed(input_fmap_142[7:0]) +
	( 13'sd 3521) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11871) * $signed(input_fmap_144[7:0]) +
	( 11'sd 897) * $signed(input_fmap_145[7:0]) +
	( 7'sd 35) * $signed(input_fmap_146[7:0]) +
	( 15'sd 10098) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6995) * $signed(input_fmap_148[7:0]) +
	( 16'sd 21586) * $signed(input_fmap_149[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_150[7:0]) +
	( 15'sd 9286) * $signed(input_fmap_151[7:0]) +
	( 14'sd 5576) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14326) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23007) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13105) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28442) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23153) * $signed(input_fmap_157[7:0]) +
	( 16'sd 24348) * $signed(input_fmap_158[7:0]) +
	( 16'sd 19213) * $signed(input_fmap_159[7:0]) +
	( 16'sd 29349) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19435) * $signed(input_fmap_161[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28864) * $signed(input_fmap_163[7:0]) +
	( 16'sd 21024) * $signed(input_fmap_164[7:0]) +
	( 15'sd 8841) * $signed(input_fmap_165[7:0]) +
	( 16'sd 23870) * $signed(input_fmap_166[7:0]) +
	( 16'sd 27512) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17402) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10922) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14467) * $signed(input_fmap_170[7:0]) +
	( 16'sd 28286) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7737) * $signed(input_fmap_172[7:0]) +
	( 16'sd 22467) * $signed(input_fmap_173[7:0]) +
	( 14'sd 5623) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25070) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1123) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22181) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27253) * $signed(input_fmap_178[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_179[7:0]) +
	( 14'sd 5569) * $signed(input_fmap_180[7:0]) +
	( 15'sd 14382) * $signed(input_fmap_181[7:0]) +
	( 16'sd 25637) * $signed(input_fmap_182[7:0]) +
	( 15'sd 9989) * $signed(input_fmap_183[7:0]) +
	( 15'sd 16055) * $signed(input_fmap_184[7:0]) +
	( 16'sd 16420) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_186[7:0]) +
	( 16'sd 19834) * $signed(input_fmap_187[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_189[7:0]) +
	( 13'sd 2215) * $signed(input_fmap_190[7:0]) +
	( 16'sd 22624) * $signed(input_fmap_191[7:0]) +
	( 15'sd 10023) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27996) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30751) * $signed(input_fmap_194[7:0]) +
	( 15'sd 11628) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22679) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15176) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29797) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12165) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_200[7:0]) +
	( 14'sd 4200) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7257) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2271) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2278) * $signed(input_fmap_204[7:0]) +
	( 15'sd 14971) * $signed(input_fmap_205[7:0]) +
	( 16'sd 32427) * $signed(input_fmap_206[7:0]) +
	( 16'sd 24573) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_208[7:0]) +
	( 14'sd 6115) * $signed(input_fmap_209[7:0]) +
	( 16'sd 24076) * $signed(input_fmap_210[7:0]) +
	( 10'sd 306) * $signed(input_fmap_211[7:0]) +
	( 16'sd 20718) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_213[7:0]) +
	( 16'sd 22207) * $signed(input_fmap_214[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_215[7:0]) +
	( 15'sd 12238) * $signed(input_fmap_216[7:0]) +
	( 16'sd 29897) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5445) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15354) * $signed(input_fmap_219[7:0]) +
	( 16'sd 23845) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15931) * $signed(input_fmap_221[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_222[7:0]) +
	( 14'sd 6144) * $signed(input_fmap_223[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_224[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29756) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2825) * $signed(input_fmap_228[7:0]) +
	( 16'sd 28849) * $signed(input_fmap_229[7:0]) +
	( 16'sd 19091) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_231[7:0]) +
	( 16'sd 25659) * $signed(input_fmap_232[7:0]) +
	( 16'sd 19321) * $signed(input_fmap_233[7:0]) +
	( 16'sd 20741) * $signed(input_fmap_234[7:0]) +
	( 16'sd 27124) * $signed(input_fmap_235[7:0]) +
	( 15'sd 15489) * $signed(input_fmap_236[7:0]) +
	( 16'sd 30041) * $signed(input_fmap_237[7:0]) +
	( 16'sd 26536) * $signed(input_fmap_238[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26433) * $signed(input_fmap_240[7:0]) +
	( 14'sd 8168) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17608) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2436) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22725) * $signed(input_fmap_245[7:0]) +
	( 16'sd 29954) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18755) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3002) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_249[7:0]) +
	( 16'sd 19663) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18227) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5616) * $signed(input_fmap_252[7:0]) +
	( 16'sd 32385) * $signed(input_fmap_253[7:0]) +
	( 16'sd 18846) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23886) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_20;
assign conv_mac_20 = 
	( 15'sd 12757) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28116) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26166) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23146) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32140) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17451) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2585) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2636) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2061) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30431) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9680) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7094) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11043) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15135) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11900) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13710) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22651) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12549) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23215) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17578) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29279) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24359) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29792) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7210) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17689) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1913) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11448) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3636) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11298) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28388) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31933) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2870) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7785) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12355) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11509) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7550) * $signed(input_fmap_38[7:0]) +
	( 14'sd 8114) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1597) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15497) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9530) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2065) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17490) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30489) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5804) * $signed(input_fmap_46[7:0]) +
	( 10'sd 388) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9300) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32059) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30796) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10861) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22481) * $signed(input_fmap_52[7:0]) +
	( 9'sd 181) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24567) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25130) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13014) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24759) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19515) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3679) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2375) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27043) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23296) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13387) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11846) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3747) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27892) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29982) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21282) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19140) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13813) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7241) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4550) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21930) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20259) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16070) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17890) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19861) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28126) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15980) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21856) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21328) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26960) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13805) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21981) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31446) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13775) * $signed(input_fmap_92[7:0]) +
	( 11'sd 953) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18584) * $signed(input_fmap_94[7:0]) +
	( 11'sd 797) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8599) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4181) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31182) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1804) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26373) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2519) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3647) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11733) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2212) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9200) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21487) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17073) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19772) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25202) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18958) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5540) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5914) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4666) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15060) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12382) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1617) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9967) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6446) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17294) * $signed(input_fmap_123[7:0]) +
	( 13'sd 4011) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27900) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30463) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_127[7:0]) +
	( 16'sd 28134) * $signed(input_fmap_128[7:0]) +
	( 16'sd 22651) * $signed(input_fmap_129[7:0]) +
	( 16'sd 21934) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24652) * $signed(input_fmap_131[7:0]) +
	( 16'sd 20234) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_133[7:0]) +
	( 16'sd 22681) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32351) * $signed(input_fmap_135[7:0]) +
	( 16'sd 26671) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25643) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22271) * $signed(input_fmap_138[7:0]) +
	( 15'sd 15139) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15232) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31772) * $signed(input_fmap_141[7:0]) +
	( 12'sd 1210) * $signed(input_fmap_142[7:0]) +
	( 15'sd 8252) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22631) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19838) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13767) * $signed(input_fmap_147[7:0]) +
	( 11'sd 586) * $signed(input_fmap_148[7:0]) +
	( 15'sd 13124) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9599) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12642) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31277) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17183) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6816) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13174) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18591) * $signed(input_fmap_157[7:0]) +
	( 16'sd 32648) * $signed(input_fmap_158[7:0]) +
	( 16'sd 19146) * $signed(input_fmap_159[7:0]) +
	( 15'sd 9147) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4581) * $signed(input_fmap_161[7:0]) +
	( 15'sd 9881) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28561) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9506) * $signed(input_fmap_164[7:0]) +
	( 12'sd 1127) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3687) * $signed(input_fmap_166[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_167[7:0]) +
	( 16'sd 22516) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10644) * $signed(input_fmap_169[7:0]) +
	( 16'sd 32009) * $signed(input_fmap_170[7:0]) +
	( 16'sd 28039) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19679) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18868) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3527) * $signed(input_fmap_175[7:0]) +
	( 16'sd 31352) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31756) * $signed(input_fmap_177[7:0]) +
	( 16'sd 24530) * $signed(input_fmap_178[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_179[7:0]) +
	( 16'sd 20452) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18956) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5421) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29787) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8966) * $signed(input_fmap_184[7:0]) +
	( 15'sd 8430) * $signed(input_fmap_185[7:0]) +
	( 16'sd 20158) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9057) * $signed(input_fmap_187[7:0]) +
	( 15'sd 11527) * $signed(input_fmap_188[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30154) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_191[7:0]) +
	( 16'sd 32463) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12083) * $signed(input_fmap_193[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_194[7:0]) +
	( 13'sd 2499) * $signed(input_fmap_195[7:0]) +
	( 11'sd 701) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18601) * $signed(input_fmap_198[7:0]) +
	( 6'sd 31) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29843) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_201[7:0]) +
	( 15'sd 10468) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12384) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15192) * $signed(input_fmap_204[7:0]) +
	( 16'sd 27502) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_206[7:0]) +
	( 15'sd 14381) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22400) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22329) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30133) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1904) * $signed(input_fmap_212[7:0]) +
	( 16'sd 18965) * $signed(input_fmap_213[7:0]) +
	( 11'sd 563) * $signed(input_fmap_214[7:0]) +
	( 11'sd 660) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_216[7:0]) +
	( 16'sd 27303) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28294) * $signed(input_fmap_218[7:0]) +
	( 15'sd 9635) * $signed(input_fmap_219[7:0]) +
	( 16'sd 27354) * $signed(input_fmap_220[7:0]) +
	( 16'sd 17626) * $signed(input_fmap_221[7:0]) +
	( 16'sd 27930) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24875) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7985) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5100) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7891) * $signed(input_fmap_226[7:0]) +
	( 16'sd 25606) * $signed(input_fmap_227[7:0]) +
	( 15'sd 16261) * $signed(input_fmap_228[7:0]) +
	( 16'sd 19405) * $signed(input_fmap_229[7:0]) +
	( 16'sd 19595) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1213) * $signed(input_fmap_231[7:0]) +
	( 14'sd 4868) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18937) * $signed(input_fmap_233[7:0]) +
	( 16'sd 26787) * $signed(input_fmap_234[7:0]) +
	( 15'sd 13938) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25616) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2639) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16490) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23787) * $signed(input_fmap_239[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_240[7:0]) +
	( 13'sd 2451) * $signed(input_fmap_241[7:0]) +
	( 14'sd 4140) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7114) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13810) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15470) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9616) * $signed(input_fmap_247[7:0]) +
	( 15'sd 15200) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9064) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_250[7:0]) +
	( 16'sd 30026) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26237) * $signed(input_fmap_252[7:0]) +
	( 16'sd 23442) * $signed(input_fmap_253[7:0]) +
	( 14'sd 4699) * $signed(input_fmap_254[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_21;
assign conv_mac_21 = 
	( 16'sd 29762) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12594) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6422) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10051) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12634) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10217) * $signed(input_fmap_5[7:0]) +
	( 11'sd 707) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12318) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28607) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10774) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24633) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23470) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5975) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32617) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10161) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19164) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30444) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24614) * $signed(input_fmap_18[7:0]) +
	( 7'sd 37) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18143) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32543) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17865) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32190) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3972) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20843) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25198) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13372) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20122) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18300) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19098) * $signed(input_fmap_31[7:0]) +
	( 6'sd 25) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3789) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11309) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6707) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2794) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1924) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18315) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11767) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11967) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10840) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5371) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13515) * $signed(input_fmap_43[7:0]) +
	( 11'sd 947) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32262) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17365) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14755) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10145) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20459) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12238) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28412) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22269) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18692) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11538) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25625) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24221) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8467) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29401) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29028) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12131) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7967) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24947) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22417) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30934) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22496) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25863) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6505) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11451) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27129) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31565) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27644) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27002) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14837) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18337) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30384) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16765) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20328) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21088) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17742) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12539) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31156) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11649) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8399) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6977) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16913) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7714) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29162) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2437) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26836) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14298) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30888) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7322) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15902) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31690) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13060) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13305) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15876) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31193) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4891) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25755) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26889) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2494) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21029) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12479) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25793) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10554) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32591) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14257) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5347) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3719) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14423) * $signed(input_fmap_124[7:0]) +
	( 15'sd 15985) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30938) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6052) * $signed(input_fmap_127[7:0]) +
	( 16'sd 22749) * $signed(input_fmap_128[7:0]) +
	( 15'sd 8964) * $signed(input_fmap_129[7:0]) +
	( 13'sd 3822) * $signed(input_fmap_130[7:0]) +
	( 11'sd 977) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18820) * $signed(input_fmap_132[7:0]) +
	( 15'sd 9900) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5135) * $signed(input_fmap_134[7:0]) +
	( 15'sd 12075) * $signed(input_fmap_135[7:0]) +
	( 16'sd 26135) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13129) * $signed(input_fmap_137[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27644) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30376) * $signed(input_fmap_140[7:0]) +
	( 16'sd 17664) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27572) * $signed(input_fmap_142[7:0]) +
	( 13'sd 3638) * $signed(input_fmap_143[7:0]) +
	( 15'sd 16054) * $signed(input_fmap_144[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_145[7:0]) +
	( 14'sd 6711) * $signed(input_fmap_146[7:0]) +
	( 16'sd 20690) * $signed(input_fmap_147[7:0]) +
	( 8'sd 72) * $signed(input_fmap_148[7:0]) +
	( 14'sd 5801) * $signed(input_fmap_149[7:0]) +
	( 16'sd 22195) * $signed(input_fmap_150[7:0]) +
	( 15'sd 11047) * $signed(input_fmap_151[7:0]) +
	( 16'sd 32186) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24717) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6393) * $signed(input_fmap_154[7:0]) +
	( 13'sd 3372) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25279) * $signed(input_fmap_157[7:0]) +
	( 14'sd 6567) * $signed(input_fmap_158[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_159[7:0]) +
	( 13'sd 3315) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31051) * $signed(input_fmap_161[7:0]) +
	( 16'sd 22040) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30729) * $signed(input_fmap_163[7:0]) +
	( 16'sd 23176) * $signed(input_fmap_164[7:0]) +
	( 13'sd 3862) * $signed(input_fmap_165[7:0]) +
	( 14'sd 7639) * $signed(input_fmap_166[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6737) * $signed(input_fmap_168[7:0]) +
	( 16'sd 32136) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24851) * $signed(input_fmap_170[7:0]) +
	( 15'sd 8335) * $signed(input_fmap_171[7:0]) +
	( 14'sd 5287) * $signed(input_fmap_172[7:0]) +
	( 16'sd 32095) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26192) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3571) * $signed(input_fmap_175[7:0]) +
	( 16'sd 23204) * $signed(input_fmap_176[7:0]) +
	( 15'sd 11444) * $signed(input_fmap_177[7:0]) +
	( 16'sd 18833) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5202) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24342) * $signed(input_fmap_180[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_181[7:0]) +
	( 15'sd 9455) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27684) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11617) * $signed(input_fmap_184[7:0]) +
	( 14'sd 4904) * $signed(input_fmap_185[7:0]) +
	( 16'sd 19447) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5983) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31950) * $signed(input_fmap_188[7:0]) +
	( 15'sd 13997) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20462) * $signed(input_fmap_190[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_191[7:0]) +
	( 15'sd 16154) * $signed(input_fmap_192[7:0]) +
	( 14'sd 4876) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27763) * $signed(input_fmap_194[7:0]) +
	( 11'sd 738) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15171) * $signed(input_fmap_196[7:0]) +
	( 9'sd 253) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9004) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29990) * $signed(input_fmap_199[7:0]) +
	( 11'sd 615) * $signed(input_fmap_200[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_201[7:0]) +
	( 16'sd 16485) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2698) * $signed(input_fmap_203[7:0]) +
	( 14'sd 8159) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15870) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20561) * $signed(input_fmap_206[7:0]) +
	( 14'sd 4401) * $signed(input_fmap_207[7:0]) +
	( 16'sd 23075) * $signed(input_fmap_208[7:0]) +
	( 15'sd 16319) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1707) * $signed(input_fmap_210[7:0]) +
	( 15'sd 14080) * $signed(input_fmap_211[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6483) * $signed(input_fmap_213[7:0]) +
	( 16'sd 26413) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10598) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4164) * $signed(input_fmap_216[7:0]) +
	( 14'sd 4199) * $signed(input_fmap_217[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12786) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24951) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15233) * $signed(input_fmap_222[7:0]) +
	( 14'sd 7627) * $signed(input_fmap_223[7:0]) +
	( 15'sd 11207) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1229) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31541) * $signed(input_fmap_226[7:0]) +
	( 16'sd 18952) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24638) * $signed(input_fmap_228[7:0]) +
	( 15'sd 11274) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14782) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28260) * $signed(input_fmap_231[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_232[7:0]) +
	( 16'sd 17710) * $signed(input_fmap_233[7:0]) +
	( 10'sd 382) * $signed(input_fmap_234[7:0]) +
	( 15'sd 8685) * $signed(input_fmap_235[7:0]) +
	( 16'sd 20685) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19581) * $signed(input_fmap_237[7:0]) +
	( 16'sd 31336) * $signed(input_fmap_238[7:0]) +
	( 16'sd 30534) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6546) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26218) * $signed(input_fmap_241[7:0]) +
	( 16'sd 22017) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30806) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14129) * $signed(input_fmap_246[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_247[7:0]) +
	( 13'sd 2584) * $signed(input_fmap_248[7:0]) +
	( 14'sd 6879) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25354) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27289) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27750) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9392) * $signed(input_fmap_254[7:0]) +
	( 11'sd 680) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_22;
assign conv_mac_22 = 
	( 12'sd 1605) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25972) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24166) * $signed(input_fmap_2[7:0]) +
	( 11'sd 682) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29686) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27955) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29606) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23566) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16612) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14471) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31447) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26883) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20432) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13002) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19445) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27468) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24875) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20943) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4841) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7411) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3343) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_21[7:0]) +
	( 10'sd 498) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21667) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32009) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19794) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19271) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28863) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20852) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30258) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29893) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13899) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7156) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30178) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17539) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23971) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22167) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18133) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27349) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11816) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10105) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14029) * $signed(input_fmap_43[7:0]) +
	( 11'sd 568) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31245) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29889) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5662) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29760) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23832) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28270) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24765) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29070) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18782) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2618) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31327) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4510) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13298) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2068) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_61[7:0]) +
	( 11'sd 867) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16305) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4802) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11850) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11236) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32255) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13435) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23457) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17931) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24409) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20515) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28439) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20400) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30768) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25873) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6911) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16217) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27977) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16161) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20041) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14992) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15979) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14438) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11255) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28323) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22463) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29509) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11461) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15274) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17484) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12415) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32151) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20452) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7632) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29080) * $signed(input_fmap_100[7:0]) +
	( 13'sd 4067) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6130) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13202) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13268) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10270) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5616) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26854) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28434) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16270) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20697) * $signed(input_fmap_110[7:0]) +
	( 11'sd 670) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15676) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15776) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2304) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20874) * $signed(input_fmap_116[7:0]) +
	( 7'sd 34) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20616) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15770) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18436) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9582) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22547) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2602) * $signed(input_fmap_124[7:0]) +
	( 10'sd 395) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30737) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32111) * $signed(input_fmap_127[7:0]) +
	( 16'sd 26616) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17777) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_130[7:0]) +
	( 16'sd 16959) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10422) * $signed(input_fmap_132[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_133[7:0]) +
	( 16'sd 29886) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23990) * $signed(input_fmap_135[7:0]) +
	( 16'sd 18413) * $signed(input_fmap_136[7:0]) +
	( 16'sd 30357) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9174) * $signed(input_fmap_138[7:0]) +
	( 15'sd 15251) * $signed(input_fmap_139[7:0]) +
	( 16'sd 31780) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3009) * $signed(input_fmap_141[7:0]) +
	( 16'sd 20142) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23196) * $signed(input_fmap_143[7:0]) +
	( 12'sd 1368) * $signed(input_fmap_144[7:0]) +
	( 16'sd 24875) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19518) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17481) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21181) * $signed(input_fmap_148[7:0]) +
	( 14'sd 6786) * $signed(input_fmap_149[7:0]) +
	( 16'sd 29003) * $signed(input_fmap_150[7:0]) +
	( 14'sd 7654) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30220) * $signed(input_fmap_152[7:0]) +
	( 16'sd 32315) * $signed(input_fmap_153[7:0]) +
	( 16'sd 17283) * $signed(input_fmap_154[7:0]) +
	( 15'sd 14113) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_157[7:0]) +
	( 14'sd 7188) * $signed(input_fmap_158[7:0]) +
	( 16'sd 19847) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18420) * $signed(input_fmap_160[7:0]) +
	( 16'sd 25765) * $signed(input_fmap_161[7:0]) +
	( 16'sd 23058) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32495) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6840) * $signed(input_fmap_164[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_165[7:0]) +
	( 10'sd 377) * $signed(input_fmap_166[7:0]) +
	( 11'sd 615) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14599) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_169[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11716) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19416) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29244) * $signed(input_fmap_173[7:0]) +
	( 16'sd 24118) * $signed(input_fmap_174[7:0]) +
	( 16'sd 22578) * $signed(input_fmap_175[7:0]) +
	( 16'sd 16386) * $signed(input_fmap_176[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_177[7:0]) +
	( 9'sd 154) * $signed(input_fmap_178[7:0]) +
	( 16'sd 29891) * $signed(input_fmap_179[7:0]) +
	( 16'sd 18371) * $signed(input_fmap_180[7:0]) +
	( 15'sd 12995) * $signed(input_fmap_181[7:0]) +
	( 15'sd 14841) * $signed(input_fmap_182[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11450) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3680) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3861) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1631) * $signed(input_fmap_187[7:0]) +
	( 16'sd 26287) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7609) * $signed(input_fmap_189[7:0]) +
	( 15'sd 12119) * $signed(input_fmap_190[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_191[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_192[7:0]) +
	( 16'sd 23251) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_194[7:0]) +
	( 11'sd 668) * $signed(input_fmap_195[7:0]) +
	( 16'sd 30838) * $signed(input_fmap_196[7:0]) +
	( 15'sd 12794) * $signed(input_fmap_197[7:0]) +
	( 14'sd 6462) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12192) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20918) * $signed(input_fmap_200[7:0]) +
	( 14'sd 5001) * $signed(input_fmap_201[7:0]) +
	( 16'sd 28758) * $signed(input_fmap_202[7:0]) +
	( 13'sd 3622) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5252) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31962) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28959) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12802) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12197) * $signed(input_fmap_208[7:0]) +
	( 14'sd 8018) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5127) * $signed(input_fmap_210[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1210) * $signed(input_fmap_212[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_213[7:0]) +
	( 16'sd 25317) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_216[7:0]) +
	( 12'sd 1180) * $signed(input_fmap_217[7:0]) +
	( 16'sd 20603) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_219[7:0]) +
	( 15'sd 15557) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28864) * $signed(input_fmap_221[7:0]) +
	( 15'sd 9157) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24404) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1429) * $signed(input_fmap_224[7:0]) +
	( 11'sd 630) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14240) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24625) * $signed(input_fmap_227[7:0]) +
	( 16'sd 27304) * $signed(input_fmap_228[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_229[7:0]) +
	( 16'sd 31717) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28250) * $signed(input_fmap_231[7:0]) +
	( 11'sd 677) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14354) * $signed(input_fmap_233[7:0]) +
	( 16'sd 27888) * $signed(input_fmap_234[7:0]) +
	( 14'sd 4647) * $signed(input_fmap_235[7:0]) +
	( 16'sd 19347) * $signed(input_fmap_236[7:0]) +
	( 16'sd 30352) * $signed(input_fmap_237[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_238[7:0]) +
	( 12'sd 1106) * $signed(input_fmap_239[7:0]) +
	( 15'sd 13285) * $signed(input_fmap_240[7:0]) +
	( 16'sd 28702) * $signed(input_fmap_241[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31482) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24737) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30408) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23069) * $signed(input_fmap_246[7:0]) +
	( 15'sd 14794) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4844) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24705) * $signed(input_fmap_249[7:0]) +
	( 14'sd 6053) * $signed(input_fmap_250[7:0]) +
	( 16'sd 28477) * $signed(input_fmap_251[7:0]) +
	( 16'sd 21516) * $signed(input_fmap_252[7:0]) +
	( 12'sd 1792) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19697) * $signed(input_fmap_254[7:0]) +
	( 16'sd 28697) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_23;
assign conv_mac_23 = 
	( 16'sd 29222) * $signed(input_fmap_0[7:0]) +
	( 11'sd 565) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18310) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26544) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26201) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17315) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11606) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1157) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11916) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27158) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14696) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25049) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29682) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3973) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16855) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24567) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16507) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8862) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1704) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5956) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28198) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12749) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27001) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6861) * $signed(input_fmap_29[7:0]) +
	( 8'sd 122) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3224) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18778) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1285) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6939) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10158) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17821) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9556) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1221) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12942) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26263) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30953) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24377) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9050) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7302) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32555) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21844) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22071) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6190) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4320) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19625) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26299) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14549) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1059) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7501) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29758) * $signed(input_fmap_57[7:0]) +
	( 11'sd 635) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8417) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31033) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29802) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2064) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27984) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5887) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14266) * $signed(input_fmap_65[7:0]) +
	( 11'sd 952) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28744) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8565) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23899) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26629) * $signed(input_fmap_70[7:0]) +
	( 11'sd 687) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21545) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31844) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25622) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12576) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4475) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28017) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29052) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3918) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10936) * $signed(input_fmap_80[7:0]) +
	( 11'sd 530) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19804) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10244) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6464) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2416) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23419) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17958) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21765) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31169) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6584) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3868) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1396) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31142) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31503) * $signed(input_fmap_97[7:0]) +
	( 10'sd 483) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32019) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27018) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26454) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10546) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1913) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18275) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11966) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10555) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20230) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24272) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30372) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2908) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6526) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28345) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4771) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12149) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30132) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6044) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7561) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20059) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13326) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24499) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7748) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5615) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22016) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31457) * $signed(input_fmap_128[7:0]) +
	( 15'sd 16305) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_130[7:0]) +
	( 16'sd 32670) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8736) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28943) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18632) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23548) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1636) * $signed(input_fmap_136[7:0]) +
	( 15'sd 10240) * $signed(input_fmap_137[7:0]) +
	( 15'sd 14139) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2843) * $signed(input_fmap_139[7:0]) +
	( 16'sd 19154) * $signed(input_fmap_140[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6198) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23766) * $signed(input_fmap_143[7:0]) +
	( 15'sd 15917) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8979) * $signed(input_fmap_145[7:0]) +
	( 16'sd 32593) * $signed(input_fmap_146[7:0]) +
	( 16'sd 23451) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23487) * $signed(input_fmap_148[7:0]) +
	( 14'sd 6368) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15671) * $signed(input_fmap_150[7:0]) +
	( 16'sd 27491) * $signed(input_fmap_151[7:0]) +
	( 15'sd 13187) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23860) * $signed(input_fmap_153[7:0]) +
	( 10'sd 347) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23022) * $signed(input_fmap_155[7:0]) +
	( 15'sd 16132) * $signed(input_fmap_156[7:0]) +
	( 14'sd 7798) * $signed(input_fmap_157[7:0]) +
	( 13'sd 2174) * $signed(input_fmap_158[7:0]) +
	( 14'sd 7189) * $signed(input_fmap_159[7:0]) +
	( 15'sd 9290) * $signed(input_fmap_160[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29882) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3619) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12521) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20392) * $signed(input_fmap_167[7:0]) +
	( 15'sd 16004) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28715) * $signed(input_fmap_170[7:0]) +
	( 16'sd 26380) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19628) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1971) * $signed(input_fmap_173[7:0]) +
	( 16'sd 30223) * $signed(input_fmap_174[7:0]) +
	( 15'sd 9998) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_176[7:0]) +
	( 11'sd 523) * $signed(input_fmap_177[7:0]) +
	( 15'sd 11740) * $signed(input_fmap_178[7:0]) +
	( 16'sd 21804) * $signed(input_fmap_179[7:0]) +
	( 15'sd 12480) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11796) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12286) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5284) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22672) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15151) * $signed(input_fmap_185[7:0]) +
	( 8'sd 92) * $signed(input_fmap_186[7:0]) +
	( 15'sd 13198) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23998) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9430) * $signed(input_fmap_190[7:0]) +
	( 15'sd 15492) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22496) * $signed(input_fmap_192[7:0]) +
	( 15'sd 14642) * $signed(input_fmap_193[7:0]) +
	( 16'sd 20643) * $signed(input_fmap_194[7:0]) +
	( 15'sd 12832) * $signed(input_fmap_195[7:0]) +
	( 14'sd 4870) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18369) * $signed(input_fmap_198[7:0]) +
	( 16'sd 32735) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8212) * $signed(input_fmap_200[7:0]) +
	( 16'sd 30229) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8625) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6415) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15850) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2588) * $signed(input_fmap_206[7:0]) +
	( 13'sd 2680) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30723) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10352) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26193) * $signed(input_fmap_211[7:0]) +
	( 14'sd 4322) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12645) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14331) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10956) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28630) * $signed(input_fmap_216[7:0]) +
	( 14'sd 8020) * $signed(input_fmap_217[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21457) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28449) * $signed(input_fmap_220[7:0]) +
	( 15'sd 11684) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_222[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13443) * $signed(input_fmap_224[7:0]) +
	( 5'sd 13) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6858) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13625) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18018) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24626) * $signed(input_fmap_229[7:0]) +
	( 15'sd 13032) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_231[7:0]) +
	( 13'sd 2703) * $signed(input_fmap_232[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_233[7:0]) +
	( 16'sd 31433) * $signed(input_fmap_234[7:0]) +
	( 13'sd 2560) * $signed(input_fmap_235[7:0]) +
	( 16'sd 29764) * $signed(input_fmap_236[7:0]) +
	( 14'sd 4737) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23801) * $signed(input_fmap_238[7:0]) +
	( 11'sd 760) * $signed(input_fmap_239[7:0]) +
	( 16'sd 30137) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32501) * $signed(input_fmap_241[7:0]) +
	( 16'sd 21190) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10954) * $signed(input_fmap_243[7:0]) +
	( 15'sd 14342) * $signed(input_fmap_244[7:0]) +
	( 16'sd 17225) * $signed(input_fmap_245[7:0]) +
	( 16'sd 29910) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9964) * $signed(input_fmap_247[7:0]) +
	( 14'sd 7162) * $signed(input_fmap_248[7:0]) +
	( 15'sd 8977) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24878) * $signed(input_fmap_250[7:0]) +
	( 16'sd 25207) * $signed(input_fmap_251[7:0]) +
	( 8'sd 82) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2258) * $signed(input_fmap_253[7:0]) +
	( 16'sd 17388) * $signed(input_fmap_254[7:0]) +
	( 14'sd 6833) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_24;
assign conv_mac_24 = 
	( 16'sd 22875) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3738) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31052) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13390) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27190) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12015) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23889) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7642) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20308) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20918) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20848) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6461) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21361) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13291) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12237) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3295) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24282) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19246) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_18[7:0]) +
	( 11'sd 924) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3995) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3024) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23309) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18919) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4213) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31980) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2867) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24370) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3887) * $signed(input_fmap_30[7:0]) +
	( 10'sd 354) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31669) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6260) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1208) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4602) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11563) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12365) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22445) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3258) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7027) * $signed(input_fmap_40[7:0]) +
	( 14'sd 8093) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16774) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11854) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10455) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17948) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13968) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29192) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25330) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26797) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24522) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7808) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16779) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12290) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12390) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28196) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29167) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2377) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24108) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24923) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9752) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21740) * $signed(input_fmap_64[7:0]) +
	( 11'sd 905) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25198) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22500) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25404) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20145) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24604) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14923) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2351) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18247) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24893) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3053) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12893) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12176) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6268) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18558) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29260) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21834) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1839) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6441) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2545) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30915) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15291) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20980) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15164) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31581) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24848) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20476) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15663) * $signed(input_fmap_96[7:0]) +
	( 9'sd 169) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3601) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4097) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13464) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18384) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2331) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26849) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13692) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16196) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29790) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3687) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31911) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30124) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11844) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19863) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2766) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10086) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15760) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26689) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13353) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7726) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5935) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18270) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15901) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31381) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5007) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23645) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21524) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1026) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_127[7:0]) +
	( 16'sd 19070) * $signed(input_fmap_128[7:0]) +
	( 16'sd 16653) * $signed(input_fmap_129[7:0]) +
	( 15'sd 11343) * $signed(input_fmap_130[7:0]) +
	( 15'sd 16194) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18924) * $signed(input_fmap_132[7:0]) +
	( 11'sd 799) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_134[7:0]) +
	( 13'sd 2477) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_136[7:0]) +
	( 15'sd 8294) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17510) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21070) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17238) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31187) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21881) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26778) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28832) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7807) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24974) * $signed(input_fmap_146[7:0]) +
	( 14'sd 7590) * $signed(input_fmap_147[7:0]) +
	( 14'sd 5781) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15257) * $signed(input_fmap_149[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3002) * $signed(input_fmap_151[7:0]) +
	( 12'sd 2031) * $signed(input_fmap_152[7:0]) +
	( 16'sd 29098) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7186) * $signed(input_fmap_154[7:0]) +
	( 16'sd 29035) * $signed(input_fmap_155[7:0]) +
	( 16'sd 16523) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5641) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9262) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12462) * $signed(input_fmap_159[7:0]) +
	( 15'sd 9770) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4382) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_162[7:0]) +
	( 14'sd 6885) * $signed(input_fmap_163[7:0]) +
	( 16'sd 18130) * $signed(input_fmap_164[7:0]) +
	( 16'sd 25993) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30092) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31979) * $signed(input_fmap_167[7:0]) +
	( 13'sd 3338) * $signed(input_fmap_168[7:0]) +
	( 16'sd 28040) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14929) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7828) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7870) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23712) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26949) * $signed(input_fmap_174[7:0]) +
	( 15'sd 8959) * $signed(input_fmap_175[7:0]) +
	( 16'sd 24501) * $signed(input_fmap_176[7:0]) +
	( 15'sd 10415) * $signed(input_fmap_177[7:0]) +
	( 14'sd 6013) * $signed(input_fmap_178[7:0]) +
	( 16'sd 27636) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3301) * $signed(input_fmap_180[7:0]) +
	( 10'sd 290) * $signed(input_fmap_181[7:0]) +
	( 15'sd 16228) * $signed(input_fmap_182[7:0]) +
	( 14'sd 4877) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9496) * $signed(input_fmap_184[7:0]) +
	( 16'sd 23245) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18596) * $signed(input_fmap_186[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_187[7:0]) +
	( 16'sd 25132) * $signed(input_fmap_188[7:0]) +
	( 15'sd 12719) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27351) * $signed(input_fmap_190[7:0]) +
	( 15'sd 8365) * $signed(input_fmap_191[7:0]) +
	( 16'sd 26012) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15176) * $signed(input_fmap_193[7:0]) +
	( 15'sd 15709) * $signed(input_fmap_194[7:0]) +
	( 16'sd 21170) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17728) * $signed(input_fmap_196[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_197[7:0]) +
	( 15'sd 14881) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10117) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_200[7:0]) +
	( 16'sd 32128) * $signed(input_fmap_201[7:0]) +
	( 16'sd 16428) * $signed(input_fmap_202[7:0]) +
	( 16'sd 18367) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17661) * $signed(input_fmap_204[7:0]) +
	( 16'sd 25013) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5311) * $signed(input_fmap_207[7:0]) +
	( 16'sd 32182) * $signed(input_fmap_208[7:0]) +
	( 16'sd 16428) * $signed(input_fmap_209[7:0]) +
	( 16'sd 21388) * $signed(input_fmap_210[7:0]) +
	( 16'sd 19658) * $signed(input_fmap_211[7:0]) +
	( 15'sd 8699) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29875) * $signed(input_fmap_213[7:0]) +
	( 13'sd 2616) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9038) * $signed(input_fmap_215[7:0]) +
	( 16'sd 21434) * $signed(input_fmap_216[7:0]) +
	( 14'sd 5539) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10724) * $signed(input_fmap_218[7:0]) +
	( 14'sd 6502) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28845) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25278) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12281) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_223[7:0]) +
	( 11'sd 1001) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1184) * $signed(input_fmap_225[7:0]) +
	( 16'sd 26248) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14340) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24263) * $signed(input_fmap_228[7:0]) +
	( 16'sd 28168) * $signed(input_fmap_229[7:0]) +
	( 11'sd 524) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20399) * $signed(input_fmap_231[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23508) * $signed(input_fmap_233[7:0]) +
	( 9'sd 191) * $signed(input_fmap_234[7:0]) +
	( 16'sd 27592) * $signed(input_fmap_235[7:0]) +
	( 16'sd 26108) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2452) * $signed(input_fmap_237[7:0]) +
	( 15'sd 11178) * $signed(input_fmap_238[7:0]) +
	( 16'sd 27824) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22038) * $signed(input_fmap_240[7:0]) +
	( 14'sd 4158) * $signed(input_fmap_241[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20175) * $signed(input_fmap_244[7:0]) +
	( 15'sd 15487) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11822) * $signed(input_fmap_246[7:0]) +
	( 16'sd 26776) * $signed(input_fmap_247[7:0]) +
	( 16'sd 23132) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24483) * $signed(input_fmap_249[7:0]) +
	( 10'sd 505) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7628) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20812) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2896) * $signed(input_fmap_253[7:0]) +
	( 14'sd 6161) * $signed(input_fmap_254[7:0]) +
	( 16'sd 27861) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_25;
assign conv_mac_25 = 
	( 16'sd 26117) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18558) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22559) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29649) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21304) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15116) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9352) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4751) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19692) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20900) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22111) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15026) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2158) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1585) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31803) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28361) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15069) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15040) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5615) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27851) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22698) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10238) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8295) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6464) * $signed(input_fmap_24[7:0]) +
	( 15'sd 16172) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27378) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29896) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14271) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24496) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23719) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2437) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22269) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25798) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6965) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13132) * $signed(input_fmap_37[7:0]) +
	( 10'sd 440) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19486) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21360) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16777) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24917) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22105) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27927) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16175) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22808) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10816) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24432) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21352) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21614) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10120) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31698) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25139) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30526) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15145) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_58[7:0]) +
	( 11'sd 992) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31882) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23198) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5505) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24024) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17571) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25467) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5094) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2460) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25608) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15682) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19108) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14671) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1119) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30329) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20494) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14669) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7960) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9557) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12441) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21617) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26928) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5517) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20147) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6308) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23481) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22050) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27535) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28985) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9697) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31822) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5979) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15995) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19354) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12838) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1557) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1042) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29103) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23836) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21563) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32148) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6123) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30333) * $signed(input_fmap_104[7:0]) +
	( 13'sd 4043) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10622) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11241) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10313) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21161) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7551) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26149) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18760) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6991) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30576) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14160) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16786) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5632) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6073) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1361) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7673) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21611) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14563) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32353) * $signed(input_fmap_127[7:0]) +
	( 14'sd 6514) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1861) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19068) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31557) * $signed(input_fmap_131[7:0]) +
	( 11'sd 847) * $signed(input_fmap_132[7:0]) +
	( 14'sd 6415) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10121) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23979) * $signed(input_fmap_136[7:0]) +
	( 16'sd 29147) * $signed(input_fmap_137[7:0]) +
	( 16'sd 30074) * $signed(input_fmap_138[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_139[7:0]) +
	( 16'sd 32664) * $signed(input_fmap_140[7:0]) +
	( 14'sd 8136) * $signed(input_fmap_141[7:0]) +
	( 16'sd 23798) * $signed(input_fmap_142[7:0]) +
	( 15'sd 13855) * $signed(input_fmap_143[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21844) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15630) * $signed(input_fmap_146[7:0]) +
	( 13'sd 2790) * $signed(input_fmap_147[7:0]) +
	( 16'sd 30599) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15992) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18638) * $signed(input_fmap_150[7:0]) +
	( 16'sd 20660) * $signed(input_fmap_151[7:0]) +
	( 14'sd 4234) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12208) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23376) * $signed(input_fmap_154[7:0]) +
	( 16'sd 29240) * $signed(input_fmap_155[7:0]) +
	( 14'sd 5924) * $signed(input_fmap_156[7:0]) +
	( 13'sd 3774) * $signed(input_fmap_157[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_158[7:0]) +
	( 15'sd 11120) * $signed(input_fmap_159[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4571) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2068) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1126) * $signed(input_fmap_164[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_165[7:0]) +
	( 8'sd 66) * $signed(input_fmap_166[7:0]) +
	( 16'sd 19004) * $signed(input_fmap_167[7:0]) +
	( 16'sd 22149) * $signed(input_fmap_168[7:0]) +
	( 16'sd 24551) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31631) * $signed(input_fmap_170[7:0]) +
	( 16'sd 23803) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31213) * $signed(input_fmap_172[7:0]) +
	( 16'sd 22757) * $signed(input_fmap_173[7:0]) +
	( 15'sd 9459) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17960) * $signed(input_fmap_175[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27792) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9716) * $signed(input_fmap_178[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_179[7:0]) +
	( 15'sd 9190) * $signed(input_fmap_180[7:0]) +
	( 16'sd 19019) * $signed(input_fmap_181[7:0]) +
	( 16'sd 17222) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30360) * $signed(input_fmap_183[7:0]) +
	( 16'sd 18455) * $signed(input_fmap_184[7:0]) +
	( 16'sd 30904) * $signed(input_fmap_185[7:0]) +
	( 16'sd 32139) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28261) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21851) * $signed(input_fmap_188[7:0]) +
	( 16'sd 28531) * $signed(input_fmap_189[7:0]) +
	( 14'sd 8042) * $signed(input_fmap_190[7:0]) +
	( 14'sd 7170) * $signed(input_fmap_191[7:0]) +
	( 15'sd 13488) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12454) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23881) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24722) * $signed(input_fmap_195[7:0]) +
	( 16'sd 30142) * $signed(input_fmap_196[7:0]) +
	( 15'sd 12374) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_198[7:0]) +
	( 16'sd 16942) * $signed(input_fmap_199[7:0]) +
	( 11'sd 653) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9127) * $signed(input_fmap_201[7:0]) +
	( 16'sd 30574) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13941) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12222) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30602) * $signed(input_fmap_205[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15416) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22416) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3882) * $signed(input_fmap_210[7:0]) +
	( 14'sd 4471) * $signed(input_fmap_211[7:0]) +
	( 16'sd 27071) * $signed(input_fmap_212[7:0]) +
	( 16'sd 30915) * $signed(input_fmap_213[7:0]) +
	( 16'sd 25518) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6641) * $signed(input_fmap_215[7:0]) +
	( 16'sd 26688) * $signed(input_fmap_216[7:0]) +
	( 16'sd 29596) * $signed(input_fmap_217[7:0]) +
	( 14'sd 4720) * $signed(input_fmap_218[7:0]) +
	( 15'sd 13895) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28277) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28717) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25039) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12742) * $signed(input_fmap_223[7:0]) +
	( 14'sd 4441) * $signed(input_fmap_224[7:0]) +
	( 16'sd 21305) * $signed(input_fmap_225[7:0]) +
	( 14'sd 5706) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24544) * $signed(input_fmap_228[7:0]) +
	( 16'sd 28844) * $signed(input_fmap_229[7:0]) +
	( 6'sd 23) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20821) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21521) * $signed(input_fmap_233[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11214) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23737) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20985) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23060) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5631) * $signed(input_fmap_239[7:0]) +
	( 13'sd 3545) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23205) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29804) * $signed(input_fmap_242[7:0]) +
	( 15'sd 14996) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24338) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12446) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31898) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_247[7:0]) +
	( 16'sd 20333) * $signed(input_fmap_248[7:0]) +
	( 15'sd 13139) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26018) * $signed(input_fmap_251[7:0]) +
	( 12'sd 1622) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2448) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19052) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20586) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_26;
assign conv_mac_26 = 
	( 15'sd 15101) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32736) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16973) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3955) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27401) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2206) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30028) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2179) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5704) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16979) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15773) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5744) * $signed(input_fmap_12[7:0]) +
	( 9'sd 244) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18470) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25365) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5068) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31677) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31076) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19754) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27324) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12379) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13747) * $signed(input_fmap_22[7:0]) +
	( 9'sd 173) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26672) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8128) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13815) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31388) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7256) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32551) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4728) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7129) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32364) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13396) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26864) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11729) * $signed(input_fmap_36[7:0]) +
	( 11'sd 966) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22310) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11541) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22406) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6031) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8630) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21169) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30351) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22320) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7377) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28981) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7725) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12307) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13928) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2394) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6037) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16820) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3267) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20707) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14594) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12419) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20770) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17674) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5720) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32709) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16223) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29075) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1879) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30361) * $signed(input_fmap_66[7:0]) +
	( 14'sd 4975) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9009) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4439) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18198) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9320) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12451) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14796) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5652) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12627) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7218) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8860) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12665) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14211) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16159) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32621) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4317) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7150) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13493) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13274) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31539) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18024) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6244) * $signed(input_fmap_89[7:0]) +
	( 14'sd 8050) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13776) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30719) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26658) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22320) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23640) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21182) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13144) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10652) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15781) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1809) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15679) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3260) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3661) * $signed(input_fmap_103[7:0]) +
	( 10'sd 283) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7667) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14876) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27944) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13336) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20628) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18331) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2649) * $signed(input_fmap_111[7:0]) +
	( 10'sd 406) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9210) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32391) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18627) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31708) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24563) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25422) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5066) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10957) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20035) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14412) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15200) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14319) * $signed(input_fmap_129[7:0]) +
	( 16'sd 26679) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19341) * $signed(input_fmap_131[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21968) * $signed(input_fmap_133[7:0]) +
	( 14'sd 7708) * $signed(input_fmap_134[7:0]) +
	( 12'sd 1070) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17264) * $signed(input_fmap_136[7:0]) +
	( 16'sd 22620) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7779) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_139[7:0]) +
	( 14'sd 4917) * $signed(input_fmap_140[7:0]) +
	( 15'sd 11729) * $signed(input_fmap_141[7:0]) +
	( 14'sd 7626) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6796) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26253) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24418) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19228) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31142) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6115) * $signed(input_fmap_151[7:0]) +
	( 14'sd 8143) * $signed(input_fmap_152[7:0]) +
	( 16'sd 22823) * $signed(input_fmap_153[7:0]) +
	( 15'sd 15378) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22165) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24887) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18620) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21639) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26324) * $signed(input_fmap_160[7:0]) +
	( 16'sd 25757) * $signed(input_fmap_161[7:0]) +
	( 16'sd 17704) * $signed(input_fmap_162[7:0]) +
	( 16'sd 31295) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1137) * $signed(input_fmap_164[7:0]) +
	( 16'sd 25998) * $signed(input_fmap_165[7:0]) +
	( 15'sd 15920) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9674) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4981) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3716) * $signed(input_fmap_169[7:0]) +
	( 16'sd 25747) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20961) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6657) * $signed(input_fmap_172[7:0]) +
	( 15'sd 13295) * $signed(input_fmap_173[7:0]) +
	( 16'sd 31200) * $signed(input_fmap_174[7:0]) +
	( 16'sd 20518) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27844) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_177[7:0]) +
	( 14'sd 6713) * $signed(input_fmap_178[7:0]) +
	( 15'sd 11841) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3017) * $signed(input_fmap_180[7:0]) +
	( 15'sd 10951) * $signed(input_fmap_181[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_182[7:0]) +
	( 15'sd 10770) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30731) * $signed(input_fmap_184[7:0]) +
	( 16'sd 28483) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6888) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9086) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23403) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11831) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13231) * $signed(input_fmap_190[7:0]) +
	( 15'sd 16170) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12406) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11345) * $signed(input_fmap_193[7:0]) +
	( 15'sd 13587) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25046) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1047) * $signed(input_fmap_197[7:0]) +
	( 16'sd 30975) * $signed(input_fmap_198[7:0]) +
	( 14'sd 8084) * $signed(input_fmap_199[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27330) * $signed(input_fmap_201[7:0]) +
	( 8'sd 95) * $signed(input_fmap_202[7:0]) +
	( 16'sd 23022) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17898) * $signed(input_fmap_204[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_205[7:0]) +
	( 16'sd 16846) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1588) * $signed(input_fmap_207[7:0]) +
	( 16'sd 21014) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20136) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31616) * $signed(input_fmap_210[7:0]) +
	( 14'sd 7831) * $signed(input_fmap_211[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_212[7:0]) +
	( 16'sd 30795) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7993) * $signed(input_fmap_214[7:0]) +
	( 15'sd 14602) * $signed(input_fmap_215[7:0]) +
	( 15'sd 8753) * $signed(input_fmap_216[7:0]) +
	( 16'sd 23612) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13413) * $signed(input_fmap_218[7:0]) +
	( 16'sd 22962) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6430) * $signed(input_fmap_221[7:0]) +
	( 16'sd 23481) * $signed(input_fmap_222[7:0]) +
	( 16'sd 30156) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7669) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20002) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30068) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13298) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2635) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26771) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28735) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10465) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8207) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11952) * $signed(input_fmap_233[7:0]) +
	( 14'sd 6065) * $signed(input_fmap_234[7:0]) +
	( 14'sd 6425) * $signed(input_fmap_235[7:0]) +
	( 15'sd 15718) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2076) * $signed(input_fmap_237[7:0]) +
	( 16'sd 29486) * $signed(input_fmap_238[7:0]) +
	( 12'sd 1248) * $signed(input_fmap_239[7:0]) +
	( 16'sd 28164) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21908) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1994) * $signed(input_fmap_242[7:0]) +
	( 15'sd 16058) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30356) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5565) * $signed(input_fmap_245[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15852) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26744) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9855) * $signed(input_fmap_249[7:0]) +
	( 16'sd 18440) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22173) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5436) * $signed(input_fmap_252[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_253[7:0]) +
	( 15'sd 11905) * $signed(input_fmap_254[7:0]) +
	( 14'sd 4555) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_27;
assign conv_mac_27 = 
	( 16'sd 18590) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9901) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9960) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17380) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17897) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4966) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7441) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19090) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28422) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12049) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8330) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24745) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25681) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17571) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25791) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23129) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21222) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30338) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10824) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29010) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29010) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5671) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8501) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7442) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28143) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26761) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30892) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22064) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20483) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30928) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8371) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2923) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14523) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8583) * $signed(input_fmap_35[7:0]) +
	( 11'sd 552) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27049) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7635) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31220) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25372) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26598) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18246) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30392) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8475) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29010) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3153) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24345) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15579) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24793) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19598) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15535) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12659) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18056) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23158) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4151) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29036) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20169) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13979) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27022) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2188) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13722) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13839) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9422) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14342) * $signed(input_fmap_65[7:0]) +
	( 9'sd 196) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29675) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31928) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20885) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25658) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25089) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21106) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8624) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24222) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26360) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30696) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29079) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25720) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7702) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17209) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32437) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2983) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19882) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31666) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25187) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16613) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13992) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7967) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16599) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31954) * $signed(input_fmap_94[7:0]) +
	( 13'sd 4092) * $signed(input_fmap_95[7:0]) +
	( 10'sd 328) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30703) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2370) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2847) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5148) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20246) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13182) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17780) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29419) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3751) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2361) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22257) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27388) * $signed(input_fmap_109[7:0]) +
	( 13'sd 4064) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15147) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25394) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3990) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2605) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27740) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27847) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30797) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27780) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1848) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2690) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3420) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12541) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9273) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15691) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4124) * $signed(input_fmap_127[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24019) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31814) * $signed(input_fmap_130[7:0]) +
	( 16'sd 18426) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14609) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12229) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11978) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21839) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26512) * $signed(input_fmap_137[7:0]) +
	( 15'sd 13912) * $signed(input_fmap_138[7:0]) +
	( 16'sd 17519) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29768) * $signed(input_fmap_140[7:0]) +
	( 16'sd 32722) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25697) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5975) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19320) * $signed(input_fmap_144[7:0]) +
	( 16'sd 19235) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24072) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30604) * $signed(input_fmap_147[7:0]) +
	( 16'sd 18658) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2652) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18127) * $signed(input_fmap_150[7:0]) +
	( 15'sd 10458) * $signed(input_fmap_151[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_152[7:0]) +
	( 11'sd 560) * $signed(input_fmap_153[7:0]) +
	( 15'sd 12240) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19558) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13122) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27775) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20145) * $signed(input_fmap_158[7:0]) +
	( 16'sd 22129) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17977) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22409) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2996) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20935) * $signed(input_fmap_163[7:0]) +
	( 16'sd 26575) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28821) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17066) * $signed(input_fmap_167[7:0]) +
	( 15'sd 10218) * $signed(input_fmap_168[7:0]) +
	( 16'sd 31842) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_170[7:0]) +
	( 16'sd 29095) * $signed(input_fmap_171[7:0]) +
	( 16'sd 26668) * $signed(input_fmap_172[7:0]) +
	( 16'sd 22387) * $signed(input_fmap_173[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7606) * $signed(input_fmap_175[7:0]) +
	( 16'sd 30955) * $signed(input_fmap_176[7:0]) +
	( 15'sd 14720) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2601) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3688) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28155) * $signed(input_fmap_181[7:0]) +
	( 16'sd 20444) * $signed(input_fmap_182[7:0]) +
	( 12'sd 1739) * $signed(input_fmap_183[7:0]) +
	( 14'sd 4331) * $signed(input_fmap_184[7:0]) +
	( 16'sd 32069) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2102) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18289) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31866) * $signed(input_fmap_188[7:0]) +
	( 15'sd 15666) * $signed(input_fmap_189[7:0]) +
	( 16'sd 25135) * $signed(input_fmap_190[7:0]) +
	( 15'sd 12121) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28293) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11627) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30667) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5666) * $signed(input_fmap_195[7:0]) +
	( 16'sd 28839) * $signed(input_fmap_196[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10398) * $signed(input_fmap_198[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20253) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1430) * $signed(input_fmap_201[7:0]) +
	( 13'sd 3431) * $signed(input_fmap_202[7:0]) +
	( 16'sd 27317) * $signed(input_fmap_203[7:0]) +
	( 16'sd 21220) * $signed(input_fmap_204[7:0]) +
	( 16'sd 26567) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9735) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_207[7:0]) +
	( 14'sd 7121) * $signed(input_fmap_208[7:0]) +
	( 16'sd 27360) * $signed(input_fmap_209[7:0]) +
	( 16'sd 27396) * $signed(input_fmap_210[7:0]) +
	( 15'sd 11529) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29436) * $signed(input_fmap_213[7:0]) +
	( 16'sd 25293) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17885) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32225) * $signed(input_fmap_217[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_218[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22846) * $signed(input_fmap_220[7:0]) +
	( 16'sd 18761) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18926) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9069) * $signed(input_fmap_223[7:0]) +
	( 16'sd 24926) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1969) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27895) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14108) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4928) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29106) * $signed(input_fmap_229[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_230[7:0]) +
	( 14'sd 4632) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12823) * $signed(input_fmap_232[7:0]) +
	( 16'sd 29281) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15523) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29988) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5708) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14561) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23451) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9951) * $signed(input_fmap_239[7:0]) +
	( 16'sd 32352) * $signed(input_fmap_240[7:0]) +
	( 16'sd 17959) * $signed(input_fmap_241[7:0]) +
	( 9'sd 230) * $signed(input_fmap_242[7:0]) +
	( 15'sd 15544) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30977) * $signed(input_fmap_244[7:0]) +
	( 16'sd 16686) * $signed(input_fmap_245[7:0]) +
	( 16'sd 24909) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26591) * $signed(input_fmap_248[7:0]) +
	( 16'sd 22609) * $signed(input_fmap_249[7:0]) +
	( 16'sd 18035) * $signed(input_fmap_250[7:0]) +
	( 12'sd 1934) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13536) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13559) * $signed(input_fmap_253[7:0]) +
	( 16'sd 16661) * $signed(input_fmap_254[7:0]) +
	( 14'sd 6019) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_28;
assign conv_mac_28 = 
	( 16'sd 16559) * $signed(input_fmap_0[7:0]) +
	( 14'sd 8055) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14760) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11513) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6559) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2113) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4535) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27044) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10134) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5453) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26217) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9684) * $signed(input_fmap_12[7:0]) +
	( 15'sd 16286) * $signed(input_fmap_13[7:0]) +
	( 10'sd 382) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5139) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25946) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22005) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2670) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32284) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6095) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18805) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31633) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25254) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24408) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4876) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14411) * $signed(input_fmap_28[7:0]) +
	( 13'sd 4044) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4378) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26909) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19986) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2254) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23029) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25109) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6748) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22700) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1583) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25822) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6353) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29083) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18286) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26918) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6008) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20412) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23752) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5171) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29332) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6958) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26317) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10524) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6949) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26655) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9930) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32605) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22122) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18040) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10804) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8183) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18831) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7290) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24342) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20421) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17363) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13505) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1788) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25588) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1752) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3327) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27126) * $signed(input_fmap_72[7:0]) +
	( 6'sd 16) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9031) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23177) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28262) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1936) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6929) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10011) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2905) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27756) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3512) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5781) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1957) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15185) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3351) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8970) * $signed(input_fmap_88[7:0]) +
	( 9'sd 160) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6416) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20557) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30176) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16964) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16043) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13883) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13479) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21814) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9759) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29877) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26310) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11707) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12803) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31040) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30189) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7699) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1812) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12315) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26897) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25318) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1848) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23156) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13264) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10037) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18288) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4376) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27740) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32132) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29352) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18284) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24484) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23952) * $signed(input_fmap_122[7:0]) +
	( 13'sd 4021) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5305) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28981) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23559) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19120) * $signed(input_fmap_129[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_130[7:0]) +
	( 16'sd 25769) * $signed(input_fmap_131[7:0]) +
	( 16'sd 28265) * $signed(input_fmap_132[7:0]) +
	( 16'sd 23846) * $signed(input_fmap_133[7:0]) +
	( 15'sd 8641) * $signed(input_fmap_134[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4818) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4868) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17763) * $signed(input_fmap_138[7:0]) +
	( 15'sd 16083) * $signed(input_fmap_139[7:0]) +
	( 14'sd 4443) * $signed(input_fmap_140[7:0]) +
	( 16'sd 26654) * $signed(input_fmap_141[7:0]) +
	( 16'sd 20716) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10755) * $signed(input_fmap_143[7:0]) +
	( 16'sd 32063) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2944) * $signed(input_fmap_145[7:0]) +
	( 15'sd 8531) * $signed(input_fmap_146[7:0]) +
	( 12'sd 1160) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_148[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9730) * $signed(input_fmap_150[7:0]) +
	( 16'sd 25031) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6686) * $signed(input_fmap_152[7:0]) +
	( 16'sd 18433) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24554) * $signed(input_fmap_154[7:0]) +
	( 12'sd 1445) * $signed(input_fmap_155[7:0]) +
	( 9'sd 187) * $signed(input_fmap_156[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_157[7:0]) +
	( 15'sd 16345) * $signed(input_fmap_158[7:0]) +
	( 10'sd 306) * $signed(input_fmap_159[7:0]) +
	( 15'sd 15469) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19072) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_162[7:0]) +
	( 10'sd 379) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_164[7:0]) +
	( 11'sd 722) * $signed(input_fmap_165[7:0]) +
	( 16'sd 25353) * $signed(input_fmap_166[7:0]) +
	( 16'sd 22225) * $signed(input_fmap_167[7:0]) +
	( 16'sd 23245) * $signed(input_fmap_168[7:0]) +
	( 16'sd 19236) * $signed(input_fmap_169[7:0]) +
	( 15'sd 8282) * $signed(input_fmap_170[7:0]) +
	( 14'sd 6324) * $signed(input_fmap_171[7:0]) +
	( 16'sd 27019) * $signed(input_fmap_172[7:0]) +
	( 15'sd 15366) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17970) * $signed(input_fmap_175[7:0]) +
	( 16'sd 32104) * $signed(input_fmap_176[7:0]) +
	( 16'sd 28977) * $signed(input_fmap_177[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_178[7:0]) +
	( 14'sd 7316) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32176) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28190) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10112) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25079) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22510) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5240) * $signed(input_fmap_185[7:0]) +
	( 16'sd 22951) * $signed(input_fmap_186[7:0]) +
	( 16'sd 32591) * $signed(input_fmap_187[7:0]) +
	( 14'sd 5551) * $signed(input_fmap_188[7:0]) +
	( 15'sd 16225) * $signed(input_fmap_189[7:0]) +
	( 14'sd 7587) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14699) * $signed(input_fmap_191[7:0]) +
	( 16'sd 21744) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30983) * $signed(input_fmap_193[7:0]) +
	( 16'sd 22970) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22911) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11311) * $signed(input_fmap_196[7:0]) +
	( 16'sd 30654) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24780) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_199[7:0]) +
	( 15'sd 11906) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21904) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18340) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_203[7:0]) +
	( 15'sd 10133) * $signed(input_fmap_204[7:0]) +
	( 11'sd 933) * $signed(input_fmap_205[7:0]) +
	( 14'sd 5135) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17208) * $signed(input_fmap_207[7:0]) +
	( 14'sd 5747) * $signed(input_fmap_208[7:0]) +
	( 16'sd 31875) * $signed(input_fmap_209[7:0]) +
	( 16'sd 21641) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15442) * $signed(input_fmap_211[7:0]) +
	( 14'sd 8049) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6890) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29345) * $signed(input_fmap_215[7:0]) +
	( 16'sd 16747) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24355) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5393) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20439) * $signed(input_fmap_219[7:0]) +
	( 16'sd 16804) * $signed(input_fmap_220[7:0]) +
	( 16'sd 32335) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15123) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12870) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14157) * $signed(input_fmap_224[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30852) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24405) * $signed(input_fmap_227[7:0]) +
	( 13'sd 3028) * $signed(input_fmap_228[7:0]) +
	( 15'sd 11509) * $signed(input_fmap_229[7:0]) +
	( 16'sd 20815) * $signed(input_fmap_230[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_231[7:0]) +
	( 15'sd 11728) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27378) * $signed(input_fmap_233[7:0]) +
	( 13'sd 2181) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5332) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31572) * $signed(input_fmap_236[7:0]) +
	( 16'sd 25303) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12265) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20534) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22675) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26860) * $signed(input_fmap_241[7:0]) +
	( 13'sd 3297) * $signed(input_fmap_242[7:0]) +
	( 11'sd 835) * $signed(input_fmap_243[7:0]) +
	( 15'sd 14268) * $signed(input_fmap_244[7:0]) +
	( 16'sd 31166) * $signed(input_fmap_245[7:0]) +
	( 14'sd 5073) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27051) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1388) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21284) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12276) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28040) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31387) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_29;
assign conv_mac_29 = 
	( 14'sd 6961) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14617) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27570) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14955) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27869) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14068) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13527) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6269) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_8[7:0]) +
	( 9'sd 210) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15805) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8493) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6848) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25782) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4439) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8737) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11515) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29329) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29807) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5281) * $signed(input_fmap_26[7:0]) +
	( 11'sd 569) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21693) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2960) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8921) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8487) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2205) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16260) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8772) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13628) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5061) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25575) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32264) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26730) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14440) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20040) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14668) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16301) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19065) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12919) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9075) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17526) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15257) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13012) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5387) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10595) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18641) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14910) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28588) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16672) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17188) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24124) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12027) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26159) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12690) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12771) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20334) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12655) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16110) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12065) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8308) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8557) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25315) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4466) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3975) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32199) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19356) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24854) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15484) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24600) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25854) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11267) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27231) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4268) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9281) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2668) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9308) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11931) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7563) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6553) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8118) * $signed(input_fmap_93[7:0]) +
	( 11'sd 644) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7371) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20985) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17419) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28439) * $signed(input_fmap_98[7:0]) +
	( 11'sd 1002) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19253) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12212) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10713) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4870) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26583) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13154) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22495) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7128) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19713) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24042) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1969) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14046) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17427) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26539) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21076) * $signed(input_fmap_114[7:0]) +
	( 10'sd 292) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_116[7:0]) +
	( 13'sd 4002) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4308) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30866) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17341) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32183) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26281) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18374) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23036) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20440) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24748) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6130) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9943) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24131) * $signed(input_fmap_129[7:0]) +
	( 10'sd 340) * $signed(input_fmap_130[7:0]) +
	( 15'sd 11872) * $signed(input_fmap_131[7:0]) +
	( 16'sd 24481) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12160) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24312) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_135[7:0]) +
	( 16'sd 22705) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11590) * $signed(input_fmap_137[7:0]) +
	( 13'sd 2853) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24278) * $signed(input_fmap_139[7:0]) +
	( 15'sd 8304) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18830) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_142[7:0]) +
	( 16'sd 19538) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22704) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8741) * $signed(input_fmap_145[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24222) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22768) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4290) * $signed(input_fmap_149[7:0]) +
	( 12'sd 1709) * $signed(input_fmap_150[7:0]) +
	( 15'sd 9070) * $signed(input_fmap_151[7:0]) +
	( 16'sd 27459) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23322) * $signed(input_fmap_153[7:0]) +
	( 15'sd 14414) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30947) * $signed(input_fmap_155[7:0]) +
	( 14'sd 5383) * $signed(input_fmap_156[7:0]) +
	( 15'sd 9781) * $signed(input_fmap_157[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12571) * $signed(input_fmap_159[7:0]) +
	( 16'sd 25281) * $signed(input_fmap_160[7:0]) +
	( 15'sd 14167) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21211) * $signed(input_fmap_162[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_163[7:0]) +
	( 16'sd 22648) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9495) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8861) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17575) * $signed(input_fmap_167[7:0]) +
	( 16'sd 31433) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10692) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2293) * $signed(input_fmap_170[7:0]) +
	( 15'sd 13233) * $signed(input_fmap_171[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1432) * $signed(input_fmap_173[7:0]) +
	( 13'sd 2891) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7424) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20099) * $signed(input_fmap_176[7:0]) +
	( 15'sd 14024) * $signed(input_fmap_177[7:0]) +
	( 14'sd 6239) * $signed(input_fmap_178[7:0]) +
	( 13'sd 4085) * $signed(input_fmap_179[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6579) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_182[7:0]) +
	( 16'sd 20005) * $signed(input_fmap_183[7:0]) +
	( 16'sd 19703) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6908) * $signed(input_fmap_185[7:0]) +
	( 15'sd 15960) * $signed(input_fmap_186[7:0]) +
	( 15'sd 13748) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29642) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30797) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_190[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_191[7:0]) +
	( 15'sd 9412) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26797) * $signed(input_fmap_193[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_194[7:0]) +
	( 13'sd 3762) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_196[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19108) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23790) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31259) * $signed(input_fmap_200[7:0]) +
	( 14'sd 5712) * $signed(input_fmap_201[7:0]) +
	( 10'sd 371) * $signed(input_fmap_202[7:0]) +
	( 14'sd 4379) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12648) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28721) * $signed(input_fmap_205[7:0]) +
	( 15'sd 16018) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13523) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8951) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26017) * $signed(input_fmap_209[7:0]) +
	( 16'sd 20088) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5487) * $signed(input_fmap_211[7:0]) +
	( 16'sd 30748) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5789) * $signed(input_fmap_213[7:0]) +
	( 13'sd 3626) * $signed(input_fmap_214[7:0]) +
	( 16'sd 30167) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20965) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32590) * $signed(input_fmap_217[7:0]) +
	( 10'sd 411) * $signed(input_fmap_218[7:0]) +
	( 14'sd 7006) * $signed(input_fmap_219[7:0]) +
	( 15'sd 11767) * $signed(input_fmap_220[7:0]) +
	( 15'sd 14310) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_222[7:0]) +
	( 15'sd 13174) * $signed(input_fmap_223[7:0]) +
	( 16'sd 16909) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18796) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14579) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2262) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1921) * $signed(input_fmap_228[7:0]) +
	( 15'sd 15732) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7186) * $signed(input_fmap_230[7:0]) +
	( 16'sd 32017) * $signed(input_fmap_231[7:0]) +
	( 15'sd 10717) * $signed(input_fmap_232[7:0]) +
	( 10'sd 403) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5431) * $signed(input_fmap_234[7:0]) +
	( 16'sd 18741) * $signed(input_fmap_235[7:0]) +
	( 15'sd 9833) * $signed(input_fmap_236[7:0]) +
	( 15'sd 8960) * $signed(input_fmap_237[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_238[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_239[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29852) * $signed(input_fmap_241[7:0]) +
	( 15'sd 13580) * $signed(input_fmap_242[7:0]) +
	( 12'sd 1060) * $signed(input_fmap_243[7:0]) +
	( 16'sd 17724) * $signed(input_fmap_244[7:0]) +
	( 16'sd 27205) * $signed(input_fmap_245[7:0]) +
	( 15'sd 13241) * $signed(input_fmap_246[7:0]) +
	( 16'sd 31505) * $signed(input_fmap_247[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14406) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30496) * $signed(input_fmap_250[7:0]) +
	( 16'sd 24294) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13202) * $signed(input_fmap_252[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_253[7:0]) +
	( 16'sd 27098) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_30;
assign conv_mac_30 = 
	( 11'sd 964) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24614) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28248) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26384) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7774) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18815) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13070) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30604) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30160) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2982) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7097) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3696) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28305) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10628) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30790) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17151) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4150) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12155) * $signed(input_fmap_18[7:0]) +
	( 11'sd 939) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13268) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19819) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1033) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21335) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19758) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10191) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28845) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28917) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28189) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14174) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27686) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19846) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4640) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25832) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30250) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15359) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6329) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22441) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31766) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9850) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31409) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18813) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24343) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32140) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6490) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26363) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1095) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31468) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26284) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11914) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16742) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9049) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31123) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24304) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18065) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22981) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25246) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21598) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25006) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1024) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19606) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28306) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12484) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29242) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9078) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29514) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2423) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29440) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23857) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26965) * $signed(input_fmap_70[7:0]) +
	( 11'sd 1003) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29969) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28492) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28521) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24691) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16908) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20833) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23675) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12515) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2695) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13172) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10098) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11835) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20431) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14455) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21496) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17580) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16237) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15034) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20549) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28069) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21394) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_97[7:0]) +
	( 13'sd 4019) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11197) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11470) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1944) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11639) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21499) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1718) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6844) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4103) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1948) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24638) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4129) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3827) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8845) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8541) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26504) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23813) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16192) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30539) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18265) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13697) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5985) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12876) * $signed(input_fmap_124[7:0]) +
	( 11'sd 688) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20993) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22188) * $signed(input_fmap_127[7:0]) +
	( 16'sd 28508) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14690) * $signed(input_fmap_129[7:0]) +
	( 16'sd 20459) * $signed(input_fmap_130[7:0]) +
	( 14'sd 7926) * $signed(input_fmap_131[7:0]) +
	( 16'sd 19482) * $signed(input_fmap_132[7:0]) +
	( 14'sd 6465) * $signed(input_fmap_133[7:0]) +
	( 16'sd 29882) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28699) * $signed(input_fmap_135[7:0]) +
	( 15'sd 10199) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13981) * $signed(input_fmap_137[7:0]) +
	( 16'sd 20235) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24580) * $signed(input_fmap_139[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_140[7:0]) +
	( 15'sd 8302) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30119) * $signed(input_fmap_142[7:0]) +
	( 16'sd 16453) * $signed(input_fmap_143[7:0]) +
	( 16'sd 20939) * $signed(input_fmap_144[7:0]) +
	( 15'sd 10308) * $signed(input_fmap_145[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17947) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26007) * $signed(input_fmap_148[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_149[7:0]) +
	( 16'sd 20011) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_151[7:0]) +
	( 15'sd 9814) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25226) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23176) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28712) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18867) * $signed(input_fmap_157[7:0]) +
	( 16'sd 21207) * $signed(input_fmap_158[7:0]) +
	( 16'sd 17517) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27486) * $signed(input_fmap_160[7:0]) +
	( 15'sd 13132) * $signed(input_fmap_161[7:0]) +
	( 16'sd 32123) * $signed(input_fmap_162[7:0]) +
	( 14'sd 7835) * $signed(input_fmap_163[7:0]) +
	( 16'sd 17117) * $signed(input_fmap_164[7:0]) +
	( 16'sd 29538) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4966) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26430) * $signed(input_fmap_167[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11760) * $signed(input_fmap_169[7:0]) +
	( 16'sd 26698) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15572) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4940) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1030) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11134) * $signed(input_fmap_174[7:0]) +
	( 16'sd 29065) * $signed(input_fmap_175[7:0]) +
	( 15'sd 11060) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5779) * $signed(input_fmap_177[7:0]) +
	( 16'sd 19658) * $signed(input_fmap_178[7:0]) +
	( 16'sd 26821) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26436) * $signed(input_fmap_180[7:0]) +
	( 16'sd 20647) * $signed(input_fmap_181[7:0]) +
	( 13'sd 2674) * $signed(input_fmap_182[7:0]) +
	( 16'sd 16522) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8669) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6387) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17317) * $signed(input_fmap_186[7:0]) +
	( 15'sd 10662) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17721) * $signed(input_fmap_188[7:0]) +
	( 15'sd 9470) * $signed(input_fmap_189[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_190[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_191[7:0]) +
	( 14'sd 5524) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15043) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30823) * $signed(input_fmap_194[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_195[7:0]) +
	( 14'sd 4808) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32005) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27769) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14161) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18354) * $signed(input_fmap_200[7:0]) +
	( 15'sd 8710) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_202[7:0]) +
	( 15'sd 8957) * $signed(input_fmap_203[7:0]) +
	( 16'sd 20568) * $signed(input_fmap_204[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6885) * $signed(input_fmap_206[7:0]) +
	( 15'sd 14195) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28954) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18237) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17085) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29706) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30629) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5279) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18821) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25204) * $signed(input_fmap_217[7:0]) +
	( 16'sd 27186) * $signed(input_fmap_218[7:0]) +
	( 16'sd 26139) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1482) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15355) * $signed(input_fmap_221[7:0]) +
	( 16'sd 20774) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9303) * $signed(input_fmap_223[7:0]) +
	( 16'sd 23659) * $signed(input_fmap_224[7:0]) +
	( 16'sd 22197) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22966) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24909) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4449) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20356) * $signed(input_fmap_229[7:0]) +
	( 16'sd 31223) * $signed(input_fmap_230[7:0]) +
	( 15'sd 15075) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9142) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3564) * $signed(input_fmap_233[7:0]) +
	( 16'sd 30219) * $signed(input_fmap_234[7:0]) +
	( 16'sd 20907) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_236[7:0]) +
	( 15'sd 13122) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3111) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5970) * $signed(input_fmap_239[7:0]) +
	( 16'sd 16777) * $signed(input_fmap_240[7:0]) +
	( 16'sd 19258) * $signed(input_fmap_241[7:0]) +
	( 14'sd 6651) * $signed(input_fmap_242[7:0]) +
	( 16'sd 19469) * $signed(input_fmap_243[7:0]) +
	( 16'sd 29064) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19031) * $signed(input_fmap_245[7:0]) +
	( 14'sd 6124) * $signed(input_fmap_246[7:0]) +
	( 13'sd 2518) * $signed(input_fmap_247[7:0]) +
	( 16'sd 27296) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9581) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26704) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13826) * $signed(input_fmap_251[7:0]) +
	( 15'sd 8583) * $signed(input_fmap_252[7:0]) +
	( 16'sd 20776) * $signed(input_fmap_253[7:0]) +
	( 16'sd 22720) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23471) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_31;
assign conv_mac_31 = 
	( 16'sd 17472) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20404) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25157) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23259) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23141) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17100) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12347) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27831) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28409) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2347) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17659) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17548) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22927) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23351) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18550) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25237) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25989) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28015) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1743) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16100) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29746) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7863) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3745) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29795) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25556) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6895) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13530) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18860) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22278) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25405) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13671) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31503) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10446) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27148) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7209) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3357) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31673) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2646) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26702) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3939) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27125) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9605) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21193) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12135) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14111) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25835) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11531) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29358) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22517) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1460) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18389) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32250) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26459) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26926) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2853) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21729) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8240) * $signed(input_fmap_66[7:0]) +
	( 11'sd 966) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8325) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18575) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3756) * $signed(input_fmap_70[7:0]) +
	( 14'sd 8073) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31856) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13199) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9084) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4148) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3055) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10112) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16179) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29351) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18639) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25091) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9787) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16030) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30493) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7453) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12602) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20074) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20301) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21660) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17425) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3873) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26946) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10955) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29256) * $signed(input_fmap_102[7:0]) +
	( 11'sd 582) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27452) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20068) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19252) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20874) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17186) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30591) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14560) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6999) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6864) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7129) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14079) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27502) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30417) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23340) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8436) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8484) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12022) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30309) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29920) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32385) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5275) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29904) * $signed(input_fmap_128[7:0]) +
	( 13'sd 3526) * $signed(input_fmap_129[7:0]) +
	( 16'sd 24496) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19572) * $signed(input_fmap_131[7:0]) +
	( 14'sd 4360) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11534) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19325) * $signed(input_fmap_134[7:0]) +
	( 16'sd 29335) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13620) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9384) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10330) * $signed(input_fmap_138[7:0]) +
	( 16'sd 17383) * $signed(input_fmap_139[7:0]) +
	( 11'sd 904) * $signed(input_fmap_140[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_141[7:0]) +
	( 15'sd 15244) * $signed(input_fmap_142[7:0]) +
	( 16'sd 22204) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_144[7:0]) +
	( 16'sd 30954) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_146[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_147[7:0]) +
	( 16'sd 25333) * $signed(input_fmap_148[7:0]) +
	( 16'sd 32764) * $signed(input_fmap_149[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4249) * $signed(input_fmap_151[7:0]) +
	( 15'sd 11287) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_153[7:0]) +
	( 16'sd 19258) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27096) * $signed(input_fmap_155[7:0]) +
	( 13'sd 3214) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31704) * $signed(input_fmap_157[7:0]) +
	( 16'sd 30818) * $signed(input_fmap_158[7:0]) +
	( 16'sd 17919) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24636) * $signed(input_fmap_160[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_161[7:0]) +
	( 16'sd 16740) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20854) * $signed(input_fmap_163[7:0]) +
	( 14'sd 8140) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30321) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12192) * $signed(input_fmap_166[7:0]) +
	( 14'sd 5995) * $signed(input_fmap_167[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_168[7:0]) +
	( 16'sd 29679) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_170[7:0]) +
	( 15'sd 14431) * $signed(input_fmap_171[7:0]) +
	( 16'sd 26269) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_174[7:0]) +
	( 15'sd 12795) * $signed(input_fmap_175[7:0]) +
	( 16'sd 31205) * $signed(input_fmap_176[7:0]) +
	( 16'sd 21303) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10753) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21970) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11683) * $signed(input_fmap_181[7:0]) +
	( 16'sd 24051) * $signed(input_fmap_182[7:0]) +
	( 15'sd 13563) * $signed(input_fmap_183[7:0]) +
	( 15'sd 12181) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1512) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4410) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9047) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21153) * $signed(input_fmap_188[7:0]) +
	( 15'sd 15554) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32452) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28642) * $signed(input_fmap_192[7:0]) +
	( 12'sd 1863) * $signed(input_fmap_193[7:0]) +
	( 16'sd 16890) * $signed(input_fmap_194[7:0]) +
	( 15'sd 8595) * $signed(input_fmap_195[7:0]) +
	( 15'sd 8224) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14277) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29188) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_199[7:0]) +
	( 16'sd 32403) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15721) * $signed(input_fmap_201[7:0]) +
	( 16'sd 29519) * $signed(input_fmap_202[7:0]) +
	( 16'sd 18514) * $signed(input_fmap_203[7:0]) +
	( 16'sd 20901) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31825) * $signed(input_fmap_205[7:0]) +
	( 16'sd 23099) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_207[7:0]) +
	( 14'sd 5467) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7784) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23937) * $signed(input_fmap_210[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24010) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28265) * $signed(input_fmap_214[7:0]) +
	( 14'sd 4184) * $signed(input_fmap_215[7:0]) +
	( 15'sd 12815) * $signed(input_fmap_216[7:0]) +
	( 16'sd 23283) * $signed(input_fmap_217[7:0]) +
	( 16'sd 29647) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17399) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22729) * $signed(input_fmap_220[7:0]) +
	( 16'sd 20740) * $signed(input_fmap_221[7:0]) +
	( 11'sd 696) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25716) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13206) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18992) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30834) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22953) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26064) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8678) * $signed(input_fmap_229[7:0]) +
	( 15'sd 8629) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24844) * $signed(input_fmap_231[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_232[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_233[7:0]) +
	( 14'sd 6777) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7111) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25081) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28613) * $signed(input_fmap_237[7:0]) +
	( 15'sd 11755) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26683) * $signed(input_fmap_239[7:0]) +
	( 13'sd 4075) * $signed(input_fmap_240[7:0]) +
	( 14'sd 4739) * $signed(input_fmap_241[7:0]) +
	( 16'sd 22127) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25899) * $signed(input_fmap_243[7:0]) +
	( 16'sd 17406) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24409) * $signed(input_fmap_245[7:0]) +
	( 11'sd 543) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15013) * $signed(input_fmap_247[7:0]) +
	( 15'sd 16124) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21475) * $signed(input_fmap_249[7:0]) +
	( 15'sd 15622) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4754) * $signed(input_fmap_251[7:0]) +
	( 16'sd 19173) * $signed(input_fmap_252[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_253[7:0]) +
	( 15'sd 15537) * $signed(input_fmap_254[7:0]) +
	( 12'sd 1967) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_32;
assign conv_mac_32 = 
	( 16'sd 19034) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13706) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3944) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10149) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31432) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9991) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10972) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26988) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22092) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11517) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9184) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13436) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26979) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26825) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1452) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8363) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18038) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9900) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15076) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23546) * $signed(input_fmap_20[7:0]) +
	( 5'sd 13) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1335) * $signed(input_fmap_23[7:0]) +
	( 9'sd 169) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6493) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30814) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1379) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8803) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17526) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13679) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2660) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13535) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21365) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1379) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21801) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4121) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24385) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20003) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10886) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20831) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7659) * $signed(input_fmap_43[7:0]) +
	( 9'sd 161) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18191) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9388) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20504) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29387) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26094) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21002) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7849) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11532) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23419) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11309) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29114) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4551) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8472) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6895) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12536) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20311) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25047) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31373) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12908) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9051) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10451) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25937) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12365) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19108) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8409) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28224) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21249) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17870) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32170) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21861) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2414) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1648) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29607) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21537) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32241) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2324) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9459) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28693) * $signed(input_fmap_85[7:0]) +
	( 11'sd 913) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23642) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32583) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27871) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16424) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17205) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19620) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22240) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19251) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25929) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14567) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20813) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18301) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14180) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31514) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17181) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22211) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13147) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8659) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19859) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30543) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26623) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7534) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3789) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7688) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12117) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7295) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4535) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17158) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16437) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9767) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15253) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32216) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26212) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29393) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8121) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24857) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27111) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11692) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3435) * $signed(input_fmap_127[7:0]) +
	( 13'sd 3773) * $signed(input_fmap_128[7:0]) +
	( 15'sd 11716) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1628) * $signed(input_fmap_130[7:0]) +
	( 14'sd 6762) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10132) * $signed(input_fmap_132[7:0]) +
	( 16'sd 26368) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25115) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32192) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1459) * $signed(input_fmap_136[7:0]) +
	( 13'sd 3083) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29578) * $signed(input_fmap_138[7:0]) +
	( 15'sd 9213) * $signed(input_fmap_139[7:0]) +
	( 16'sd 18521) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3016) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22738) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5718) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8211) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29290) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29621) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20139) * $signed(input_fmap_148[7:0]) +
	( 16'sd 20588) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25161) * $signed(input_fmap_150[7:0]) +
	( 12'sd 1556) * $signed(input_fmap_151[7:0]) +
	( 14'sd 5695) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3095) * $signed(input_fmap_153[7:0]) +
	( 10'sd 438) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27608) * $signed(input_fmap_155[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_156[7:0]) +
	( 14'sd 7595) * $signed(input_fmap_157[7:0]) +
	( 15'sd 16316) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4805) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_160[7:0]) +
	( 16'sd 17146) * $signed(input_fmap_161[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_162[7:0]) +
	( 16'sd 21449) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13507) * $signed(input_fmap_164[7:0]) +
	( 16'sd 21013) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4770) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23497) * $signed(input_fmap_167[7:0]) +
	( 16'sd 25484) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27841) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24391) * $signed(input_fmap_170[7:0]) +
	( 15'sd 9489) * $signed(input_fmap_171[7:0]) +
	( 16'sd 32572) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27528) * $signed(input_fmap_173[7:0]) +
	( 16'sd 17085) * $signed(input_fmap_174[7:0]) +
	( 16'sd 30005) * $signed(input_fmap_175[7:0]) +
	( 15'sd 16176) * $signed(input_fmap_176[7:0]) +
	( 15'sd 11433) * $signed(input_fmap_177[7:0]) +
	( 14'sd 7216) * $signed(input_fmap_178[7:0]) +
	( 16'sd 31395) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28872) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25233) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19566) * $signed(input_fmap_182[7:0]) +
	( 14'sd 4298) * $signed(input_fmap_183[7:0]) +
	( 14'sd 7723) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1420) * $signed(input_fmap_185[7:0]) +
	( 16'sd 25130) * $signed(input_fmap_186[7:0]) +
	( 16'sd 17618) * $signed(input_fmap_187[7:0]) +
	( 16'sd 28279) * $signed(input_fmap_188[7:0]) +
	( 16'sd 28147) * $signed(input_fmap_189[7:0]) +
	( 16'sd 29089) * $signed(input_fmap_190[7:0]) +
	( 9'sd 161) * $signed(input_fmap_191[7:0]) +
	( 13'sd 2092) * $signed(input_fmap_192[7:0]) +
	( 16'sd 31960) * $signed(input_fmap_193[7:0]) +
	( 16'sd 25382) * $signed(input_fmap_194[7:0]) +
	( 14'sd 6172) * $signed(input_fmap_195[7:0]) +
	( 16'sd 30927) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14094) * $signed(input_fmap_197[7:0]) +
	( 16'sd 20554) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5016) * $signed(input_fmap_199[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16391) * $signed(input_fmap_201[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_202[7:0]) +
	( 16'sd 31235) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14739) * $signed(input_fmap_204[7:0]) +
	( 12'sd 2027) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3710) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30977) * $signed(input_fmap_207[7:0]) +
	( 16'sd 20916) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7399) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_210[7:0]) +
	( 16'sd 19228) * $signed(input_fmap_211[7:0]) +
	( 11'sd 919) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6140) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30727) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2073) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11145) * $signed(input_fmap_216[7:0]) +
	( 16'sd 18181) * $signed(input_fmap_217[7:0]) +
	( 16'sd 25872) * $signed(input_fmap_218[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_219[7:0]) +
	( 16'sd 27448) * $signed(input_fmap_220[7:0]) +
	( 16'sd 22296) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2683) * $signed(input_fmap_222[7:0]) +
	( 11'sd 547) * $signed(input_fmap_223[7:0]) +
	( 15'sd 16235) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2721) * $signed(input_fmap_225[7:0]) +
	( 16'sd 26194) * $signed(input_fmap_226[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10769) * $signed(input_fmap_228[7:0]) +
	( 16'sd 32088) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27070) * $signed(input_fmap_230[7:0]) +
	( 15'sd 8993) * $signed(input_fmap_231[7:0]) +
	( 13'sd 3611) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15296) * $signed(input_fmap_233[7:0]) +
	( 16'sd 20294) * $signed(input_fmap_234[7:0]) +
	( 15'sd 16232) * $signed(input_fmap_235[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29952) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22384) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22700) * $signed(input_fmap_239[7:0]) +
	( 8'sd 96) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20237) * $signed(input_fmap_241[7:0]) +
	( 14'sd 7300) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25325) * $signed(input_fmap_243[7:0]) +
	( 14'sd 4432) * $signed(input_fmap_244[7:0]) +
	( 16'sd 27417) * $signed(input_fmap_245[7:0]) +
	( 16'sd 24598) * $signed(input_fmap_246[7:0]) +
	( 16'sd 23153) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32078) * $signed(input_fmap_248[7:0]) +
	( 16'sd 29145) * $signed(input_fmap_249[7:0]) +
	( 16'sd 21889) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15649) * $signed(input_fmap_251[7:0]) +
	( 15'sd 11751) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11724) * $signed(input_fmap_253[7:0]) +
	( 15'sd 8914) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24288) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_33;
assign conv_mac_33 = 
	( 14'sd 7967) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3011) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15762) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19082) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26857) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19508) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3278) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11112) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11605) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21876) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19726) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28877) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24248) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17057) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15940) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22341) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7881) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3649) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8504) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29600) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22256) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11412) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23418) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31781) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25278) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5124) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3516) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1919) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17036) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24165) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15537) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8339) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15561) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1702) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24434) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7231) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23206) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23845) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18387) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15722) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11944) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28167) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1080) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4327) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15497) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23520) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31958) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21480) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24271) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5492) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16715) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32754) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27840) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31508) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31135) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24308) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24370) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13440) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6814) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23594) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31372) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14651) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3966) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6338) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30640) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16243) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22777) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11835) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3651) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30420) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26082) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26034) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23741) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10432) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17399) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5888) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18902) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24271) * $signed(input_fmap_88[7:0]) +
	( 9'sd 152) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15426) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26631) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27075) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13726) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7051) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14557) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14767) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19624) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14029) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21239) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16572) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17779) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9080) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7724) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23158) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14907) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28515) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26510) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31961) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19552) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27269) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20528) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15075) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12773) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4525) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10779) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25640) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5242) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4102) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28264) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14065) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20337) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30384) * $signed(input_fmap_128[7:0]) +
	( 16'sd 25098) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1647) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24678) * $signed(input_fmap_131[7:0]) +
	( 14'sd 7293) * $signed(input_fmap_132[7:0]) +
	( 15'sd 13684) * $signed(input_fmap_133[7:0]) +
	( 16'sd 26972) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10681) * $signed(input_fmap_135[7:0]) +
	( 15'sd 14199) * $signed(input_fmap_136[7:0]) +
	( 15'sd 14058) * $signed(input_fmap_137[7:0]) +
	( 15'sd 12119) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14562) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26487) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19835) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11033) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7515) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31218) * $signed(input_fmap_144[7:0]) +
	( 16'sd 18996) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17698) * $signed(input_fmap_147[7:0]) +
	( 12'sd 1232) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_149[7:0]) +
	( 16'sd 17557) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30023) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24252) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_153[7:0]) +
	( 15'sd 13564) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23007) * $signed(input_fmap_155[7:0]) +
	( 16'sd 23339) * $signed(input_fmap_156[7:0]) +
	( 16'sd 21517) * $signed(input_fmap_157[7:0]) +
	( 11'sd 811) * $signed(input_fmap_158[7:0]) +
	( 16'sd 23525) * $signed(input_fmap_159[7:0]) +
	( 14'sd 7418) * $signed(input_fmap_160[7:0]) +
	( 16'sd 30931) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2206) * $signed(input_fmap_162[7:0]) +
	( 15'sd 13580) * $signed(input_fmap_163[7:0]) +
	( 14'sd 7968) * $signed(input_fmap_164[7:0]) +
	( 16'sd 31094) * $signed(input_fmap_165[7:0]) +
	( 12'sd 1767) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23765) * $signed(input_fmap_167[7:0]) +
	( 15'sd 13150) * $signed(input_fmap_168[7:0]) +
	( 16'sd 29380) * $signed(input_fmap_169[7:0]) +
	( 16'sd 21296) * $signed(input_fmap_170[7:0]) +
	( 16'sd 25342) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14509) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23506) * $signed(input_fmap_173[7:0]) +
	( 16'sd 29954) * $signed(input_fmap_174[7:0]) +
	( 15'sd 16075) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10711) * $signed(input_fmap_176[7:0]) +
	( 15'sd 13194) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2741) * $signed(input_fmap_178[7:0]) +
	( 15'sd 11521) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29233) * $signed(input_fmap_180[7:0]) +
	( 16'sd 31117) * $signed(input_fmap_181[7:0]) +
	( 11'sd 723) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2321) * $signed(input_fmap_183[7:0]) +
	( 15'sd 12825) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17955) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4857) * $signed(input_fmap_187[7:0]) +
	( 14'sd 6387) * $signed(input_fmap_188[7:0]) +
	( 16'sd 23697) * $signed(input_fmap_189[7:0]) +
	( 11'sd 981) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26415) * $signed(input_fmap_191[7:0]) +
	( 15'sd 9454) * $signed(input_fmap_192[7:0]) +
	( 16'sd 21858) * $signed(input_fmap_193[7:0]) +
	( 16'sd 28814) * $signed(input_fmap_194[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22315) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22786) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19788) * $signed(input_fmap_198[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8566) * $signed(input_fmap_200[7:0]) +
	( 16'sd 24239) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_202[7:0]) +
	( 15'sd 10551) * $signed(input_fmap_203[7:0]) +
	( 13'sd 3481) * $signed(input_fmap_204[7:0]) +
	( 15'sd 9985) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21123) * $signed(input_fmap_206[7:0]) +
	( 15'sd 15328) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6800) * $signed(input_fmap_208[7:0]) +
	( 16'sd 28560) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15907) * $signed(input_fmap_211[7:0]) +
	( 16'sd 25533) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23567) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23271) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7369) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18509) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13900) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12848) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4114) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5540) * $signed(input_fmap_221[7:0]) +
	( 12'sd 1599) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9377) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25754) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26902) * $signed(input_fmap_225[7:0]) +
	( 16'sd 19301) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9369) * $signed(input_fmap_227[7:0]) +
	( 15'sd 12198) * $signed(input_fmap_228[7:0]) +
	( 16'sd 16598) * $signed(input_fmap_229[7:0]) +
	( 15'sd 11215) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13727) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9118) * $signed(input_fmap_232[7:0]) +
	( 16'sd 17822) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18068) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14015) * $signed(input_fmap_235[7:0]) +
	( 14'sd 7129) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14333) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23517) * $signed(input_fmap_238[7:0]) +
	( 14'sd 6941) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25469) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26226) * $signed(input_fmap_241[7:0]) +
	( 14'sd 7627) * $signed(input_fmap_242[7:0]) +
	( 16'sd 19693) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18143) * $signed(input_fmap_244[7:0]) +
	( 16'sd 21217) * $signed(input_fmap_245[7:0]) +
	( 14'sd 5735) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12340) * $signed(input_fmap_247[7:0]) +
	( 15'sd 11905) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4201) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_250[7:0]) +
	( 16'sd 16632) * $signed(input_fmap_251[7:0]) +
	( 9'sd 202) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_253[7:0]) +
	( 16'sd 27839) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_34;
assign conv_mac_34 = 
	( 16'sd 19453) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19975) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31667) * $signed(input_fmap_2[7:0]) +
	( 11'sd 711) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17585) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23706) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24317) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2829) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26710) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30543) * $signed(input_fmap_10[7:0]) +
	( 9'sd 144) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28114) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23041) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1052) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4271) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6898) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15053) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1102) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25814) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21123) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19861) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24342) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27475) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14950) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16546) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26151) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23520) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11750) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13296) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27134) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8902) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24364) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9047) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13921) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28017) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4407) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11985) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9259) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10188) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24985) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31432) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28763) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16460) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17448) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18316) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23048) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22039) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26080) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14913) * $signed(input_fmap_56[7:0]) +
	( 11'sd 1015) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12408) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25534) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17294) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23522) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2051) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13887) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31534) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21302) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24637) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_69[7:0]) +
	( 11'sd 672) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16663) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12948) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25828) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32470) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31858) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21795) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29382) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12526) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5533) * $signed(input_fmap_80[7:0]) +
	( 7'sd 54) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12001) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6578) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20604) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21636) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8434) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24645) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9321) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14537) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24533) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17647) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13997) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29892) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3495) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25833) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28863) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30174) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2835) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28001) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2794) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3121) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2780) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13681) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25001) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21405) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6999) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28643) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3306) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6474) * $signed(input_fmap_111[7:0]) +
	( 10'sd 301) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20021) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1551) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26439) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17510) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25585) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_121[7:0]) +
	( 12'sd 2028) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32262) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15694) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1983) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10317) * $signed(input_fmap_127[7:0]) +
	( 16'sd 22472) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13226) * $signed(input_fmap_129[7:0]) +
	( 16'sd 29132) * $signed(input_fmap_130[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_131[7:0]) +
	( 8'sd 85) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29124) * $signed(input_fmap_133[7:0]) +
	( 16'sd 26093) * $signed(input_fmap_134[7:0]) +
	( 13'sd 2683) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_136[7:0]) +
	( 15'sd 14385) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29737) * $signed(input_fmap_138[7:0]) +
	( 16'sd 29656) * $signed(input_fmap_139[7:0]) +
	( 10'sd 358) * $signed(input_fmap_140[7:0]) +
	( 15'sd 9391) * $signed(input_fmap_141[7:0]) +
	( 13'sd 2590) * $signed(input_fmap_142[7:0]) +
	( 16'sd 25603) * $signed(input_fmap_143[7:0]) +
	( 16'sd 25762) * $signed(input_fmap_144[7:0]) +
	( 15'sd 14743) * $signed(input_fmap_145[7:0]) +
	( 16'sd 30872) * $signed(input_fmap_146[7:0]) +
	( 16'sd 31163) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26053) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17775) * $signed(input_fmap_149[7:0]) +
	( 10'sd 502) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19908) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21498) * $signed(input_fmap_152[7:0]) +
	( 16'sd 29159) * $signed(input_fmap_153[7:0]) +
	( 16'sd 32228) * $signed(input_fmap_154[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_155[7:0]) +
	( 16'sd 21351) * $signed(input_fmap_156[7:0]) +
	( 13'sd 2477) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20249) * $signed(input_fmap_158[7:0]) +
	( 16'sd 31885) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31074) * $signed(input_fmap_160[7:0]) +
	( 16'sd 21184) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24164) * $signed(input_fmap_162[7:0]) +
	( 16'sd 23278) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8516) * $signed(input_fmap_164[7:0]) +
	( 16'sd 26474) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_166[7:0]) +
	( 16'sd 19891) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5433) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25922) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24338) * $signed(input_fmap_170[7:0]) +
	( 14'sd 6503) * $signed(input_fmap_171[7:0]) +
	( 16'sd 27865) * $signed(input_fmap_172[7:0]) +
	( 15'sd 15252) * $signed(input_fmap_173[7:0]) +
	( 16'sd 17653) * $signed(input_fmap_174[7:0]) +
	( 16'sd 27128) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29164) * $signed(input_fmap_176[7:0]) +
	( 15'sd 8383) * $signed(input_fmap_177[7:0]) +
	( 14'sd 5823) * $signed(input_fmap_178[7:0]) +
	( 9'sd 242) * $signed(input_fmap_179[7:0]) +
	( 16'sd 31711) * $signed(input_fmap_180[7:0]) +
	( 15'sd 14250) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4718) * $signed(input_fmap_182[7:0]) +
	( 16'sd 23808) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14426) * $signed(input_fmap_184[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_185[7:0]) +
	( 16'sd 22673) * $signed(input_fmap_186[7:0]) +
	( 16'sd 24742) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32029) * $signed(input_fmap_188[7:0]) +
	( 15'sd 8789) * $signed(input_fmap_189[7:0]) +
	( 16'sd 26705) * $signed(input_fmap_190[7:0]) +
	( 15'sd 10478) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27594) * $signed(input_fmap_192[7:0]) +
	( 16'sd 24848) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9284) * $signed(input_fmap_194[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_195[7:0]) +
	( 16'sd 16985) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26191) * $signed(input_fmap_197[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28552) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8463) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22020) * $signed(input_fmap_201[7:0]) +
	( 16'sd 24891) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5357) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5608) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21819) * $signed(input_fmap_206[7:0]) +
	( 13'sd 2332) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15577) * $signed(input_fmap_208[7:0]) +
	( 14'sd 5472) * $signed(input_fmap_209[7:0]) +
	( 16'sd 25871) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28363) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18591) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6842) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31754) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25713) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28100) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19754) * $signed(input_fmap_217[7:0]) +
	( 15'sd 16262) * $signed(input_fmap_218[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_219[7:0]) +
	( 16'sd 20910) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28750) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3108) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1678) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14121) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11082) * $signed(input_fmap_226[7:0]) +
	( 14'sd 7704) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2587) * $signed(input_fmap_228[7:0]) +
	( 15'sd 14258) * $signed(input_fmap_229[7:0]) +
	( 15'sd 9915) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18944) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15223) * $signed(input_fmap_232[7:0]) +
	( 16'sd 32357) * $signed(input_fmap_233[7:0]) +
	( 16'sd 28968) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12642) * $signed(input_fmap_235[7:0]) +
	( 11'sd 744) * $signed(input_fmap_236[7:0]) +
	( 15'sd 15658) * $signed(input_fmap_237[7:0]) +
	( 15'sd 11374) * $signed(input_fmap_238[7:0]) +
	( 13'sd 3005) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25596) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32121) * $signed(input_fmap_241[7:0]) +
	( 16'sd 30448) * $signed(input_fmap_242[7:0]) +
	( 14'sd 5741) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22199) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10880) * $signed(input_fmap_246[7:0]) +
	( 16'sd 22630) * $signed(input_fmap_247[7:0]) +
	( 15'sd 15841) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15637) * $signed(input_fmap_249[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13295) * $signed(input_fmap_251[7:0]) +
	( 16'sd 22170) * $signed(input_fmap_252[7:0]) +
	( 14'sd 7908) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1990) * $signed(input_fmap_254[7:0]) +
	( 15'sd 12028) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_35;
assign conv_mac_35 = 
	( 16'sd 19307) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8649) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30931) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27947) * $signed(input_fmap_3[7:0]) +
	( 11'sd 565) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15123) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16201) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29295) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26689) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24352) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30199) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29600) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12539) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5214) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18444) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29220) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15961) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7471) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22922) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24766) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20582) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14141) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6452) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26628) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14481) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22869) * $signed(input_fmap_26[7:0]) +
	( 14'sd 8107) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26670) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10572) * $signed(input_fmap_29[7:0]) +
	( 10'sd 292) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11739) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30981) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11028) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9724) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1134) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8596) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20906) * $signed(input_fmap_38[7:0]) +
	( 13'sd 4065) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6168) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29394) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13550) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1083) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27456) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23759) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17713) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23909) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16342) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19868) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5937) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3899) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20795) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17737) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8320) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12659) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20719) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18845) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27812) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25097) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18808) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2499) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21602) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22787) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13577) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29770) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21151) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1140) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23017) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25149) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1784) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12561) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20068) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19290) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30340) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7237) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14947) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8526) * $signed(input_fmap_80[7:0]) +
	( 9'sd 155) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22314) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21127) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29454) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9758) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13255) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20935) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14804) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5326) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29158) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2734) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30785) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7382) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5368) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11591) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17256) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18469) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21537) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7761) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27927) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5163) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14833) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3901) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32625) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17489) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30385) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15699) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13341) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1103) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5694) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1608) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4551) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21639) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19955) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22213) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12476) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9062) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16464) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20769) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23283) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10581) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31817) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31264) * $signed(input_fmap_126[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_127[7:0]) +
	( 14'sd 7114) * $signed(input_fmap_128[7:0]) +
	( 16'sd 21340) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6271) * $signed(input_fmap_130[7:0]) +
	( 16'sd 25547) * $signed(input_fmap_131[7:0]) +
	( 16'sd 21714) * $signed(input_fmap_132[7:0]) +
	( 13'sd 3043) * $signed(input_fmap_133[7:0]) +
	( 15'sd 9647) * $signed(input_fmap_134[7:0]) +
	( 16'sd 29743) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25127) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15195) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27598) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24899) * $signed(input_fmap_139[7:0]) +
	( 12'sd 2012) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3587) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6517) * $signed(input_fmap_142[7:0]) +
	( 16'sd 22125) * $signed(input_fmap_143[7:0]) +
	( 16'sd 30351) * $signed(input_fmap_144[7:0]) +
	( 11'sd 737) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1516) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11423) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20164) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18108) * $signed(input_fmap_149[7:0]) +
	( 16'sd 28252) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6217) * $signed(input_fmap_151[7:0]) +
	( 16'sd 25237) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27099) * $signed(input_fmap_153[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20198) * $signed(input_fmap_156[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_157[7:0]) +
	( 16'sd 24304) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27476) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26085) * $signed(input_fmap_160[7:0]) +
	( 15'sd 11274) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24707) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26074) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25081) * $signed(input_fmap_164[7:0]) +
	( 16'sd 26100) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_166[7:0]) +
	( 16'sd 29906) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5876) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20210) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20358) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16650) * $signed(input_fmap_171[7:0]) +
	( 16'sd 29485) * $signed(input_fmap_172[7:0]) +
	( 15'sd 15868) * $signed(input_fmap_173[7:0]) +
	( 15'sd 16135) * $signed(input_fmap_174[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_175[7:0]) +
	( 14'sd 4454) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24728) * $signed(input_fmap_177[7:0]) +
	( 15'sd 13286) * $signed(input_fmap_178[7:0]) +
	( 16'sd 24946) * $signed(input_fmap_179[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_180[7:0]) +
	( 13'sd 2122) * $signed(input_fmap_181[7:0]) +
	( 15'sd 14078) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_183[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_184[7:0]) +
	( 16'sd 18916) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4779) * $signed(input_fmap_186[7:0]) +
	( 13'sd 3056) * $signed(input_fmap_187[7:0]) +
	( 7'sd 63) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11689) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20579) * $signed(input_fmap_190[7:0]) +
	( 11'sd 888) * $signed(input_fmap_191[7:0]) +
	( 14'sd 6335) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10275) * $signed(input_fmap_193[7:0]) +
	( 15'sd 15534) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22674) * $signed(input_fmap_195[7:0]) +
	( 16'sd 27099) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11809) * $signed(input_fmap_197[7:0]) +
	( 16'sd 20502) * $signed(input_fmap_198[7:0]) +
	( 15'sd 11166) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15751) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27683) * $signed(input_fmap_201[7:0]) +
	( 16'sd 30274) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6350) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11900) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24407) * $signed(input_fmap_205[7:0]) +
	( 16'sd 32245) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30974) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11066) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_209[7:0]) +
	( 16'sd 20825) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30388) * $signed(input_fmap_211[7:0]) +
	( 15'sd 10535) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23110) * $signed(input_fmap_213[7:0]) +
	( 15'sd 11836) * $signed(input_fmap_214[7:0]) +
	( 16'sd 26857) * $signed(input_fmap_215[7:0]) +
	( 16'sd 26838) * $signed(input_fmap_216[7:0]) +
	( 16'sd 27766) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8444) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_219[7:0]) +
	( 13'sd 4055) * $signed(input_fmap_220[7:0]) +
	( 13'sd 3152) * $signed(input_fmap_221[7:0]) +
	( 16'sd 32739) * $signed(input_fmap_222[7:0]) +
	( 14'sd 7670) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7946) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15837) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6115) * $signed(input_fmap_226[7:0]) +
	( 16'sd 32728) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25010) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24004) * $signed(input_fmap_229[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_230[7:0]) +
	( 14'sd 4922) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29149) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28831) * $signed(input_fmap_233[7:0]) +
	( 16'sd 29849) * $signed(input_fmap_234[7:0]) +
	( 16'sd 17429) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10858) * $signed(input_fmap_236[7:0]) +
	( 16'sd 31220) * $signed(input_fmap_237[7:0]) +
	( 16'sd 20540) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5012) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22987) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26899) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23313) * $signed(input_fmap_242[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30978) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6714) * $signed(input_fmap_245[7:0]) +
	( 15'sd 13860) * $signed(input_fmap_246[7:0]) +
	( 16'sd 29143) * $signed(input_fmap_247[7:0]) +
	( 15'sd 8216) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_249[7:0]) +
	( 16'sd 28565) * $signed(input_fmap_250[7:0]) +
	( 16'sd 25108) * $signed(input_fmap_251[7:0]) +
	( 15'sd 16133) * $signed(input_fmap_252[7:0]) +
	( 16'sd 31976) * $signed(input_fmap_253[7:0]) +
	( 16'sd 24271) * $signed(input_fmap_254[7:0]) +
	( 16'sd 30394) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_36;
assign conv_mac_36 = 
	( 14'sd 6416) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11567) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10153) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26974) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9643) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28603) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29971) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5484) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29690) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5321) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24153) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25315) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31557) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25980) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20626) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2145) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29376) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9390) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27856) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3329) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14240) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24956) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27123) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7808) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29506) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15879) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30523) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9463) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3906) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10594) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28538) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11142) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21290) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28523) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32482) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9089) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27273) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25266) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14457) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19425) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3568) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8407) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14924) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14175) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9208) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2408) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23847) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23654) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17542) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19293) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18886) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20545) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24268) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9953) * $signed(input_fmap_63[7:0]) +
	( 9'sd 217) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17403) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28340) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21606) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14292) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23449) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8563) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22326) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14377) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2932) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22313) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31271) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26364) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27059) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26953) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1744) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24864) * $signed(input_fmap_80[7:0]) +
	( 11'sd 582) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23433) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25552) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2203) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7759) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11614) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25840) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9320) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12721) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14634) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12684) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16906) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21622) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23069) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12357) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12340) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25824) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11822) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13033) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20967) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2409) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21249) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3063) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5224) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27154) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20606) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28088) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1191) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21579) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5470) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14893) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28853) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24108) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25967) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24676) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16868) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19355) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11663) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7627) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16861) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27930) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24058) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17084) * $signed(input_fmap_127[7:0]) +
	( 14'sd 6093) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7866) * $signed(input_fmap_129[7:0]) +
	( 16'sd 21363) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3331) * $signed(input_fmap_131[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16426) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3517) * $signed(input_fmap_134[7:0]) +
	( 15'sd 8196) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1368) * $signed(input_fmap_136[7:0]) +
	( 16'sd 17906) * $signed(input_fmap_137[7:0]) +
	( 15'sd 15327) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14639) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29076) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12480) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11380) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10527) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9218) * $signed(input_fmap_144[7:0]) +
	( 15'sd 12935) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19339) * $signed(input_fmap_146[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20963) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23769) * $signed(input_fmap_149[7:0]) +
	( 14'sd 6742) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12171) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23592) * $signed(input_fmap_152[7:0]) +
	( 16'sd 28050) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24731) * $signed(input_fmap_154[7:0]) +
	( 13'sd 2931) * $signed(input_fmap_155[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27506) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14137) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17926) * $signed(input_fmap_160[7:0]) +
	( 15'sd 8298) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29581) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26959) * $signed(input_fmap_163[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30202) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9023) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_168[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24459) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3820) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12289) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_173[7:0]) +
	( 13'sd 3794) * $signed(input_fmap_174[7:0]) +
	( 16'sd 20197) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21796) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24462) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9456) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_179[7:0]) +
	( 16'sd 17261) * $signed(input_fmap_180[7:0]) +
	( 10'sd 380) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5412) * $signed(input_fmap_182[7:0]) +
	( 16'sd 20961) * $signed(input_fmap_183[7:0]) +
	( 14'sd 7607) * $signed(input_fmap_184[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_185[7:0]) +
	( 16'sd 31006) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2876) * $signed(input_fmap_187[7:0]) +
	( 16'sd 20891) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25053) * $signed(input_fmap_189[7:0]) +
	( 16'sd 22319) * $signed(input_fmap_190[7:0]) +
	( 15'sd 13507) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24915) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27844) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14663) * $signed(input_fmap_194[7:0]) +
	( 13'sd 3961) * $signed(input_fmap_195[7:0]) +
	( 14'sd 4583) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24646) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_198[7:0]) +
	( 16'sd 31849) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18904) * $signed(input_fmap_200[7:0]) +
	( 16'sd 19815) * $signed(input_fmap_201[7:0]) +
	( 16'sd 29784) * $signed(input_fmap_202[7:0]) +
	( 14'sd 7964) * $signed(input_fmap_203[7:0]) +
	( 16'sd 30245) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12595) * $signed(input_fmap_205[7:0]) +
	( 16'sd 19678) * $signed(input_fmap_206[7:0]) +
	( 14'sd 4780) * $signed(input_fmap_207[7:0]) +
	( 15'sd 9493) * $signed(input_fmap_208[7:0]) +
	( 16'sd 32728) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_210[7:0]) +
	( 15'sd 14207) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26386) * $signed(input_fmap_212[7:0]) +
	( 16'sd 17414) * $signed(input_fmap_213[7:0]) +
	( 15'sd 12124) * $signed(input_fmap_214[7:0]) +
	( 16'sd 20202) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28720) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30609) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_218[7:0]) +
	( 16'sd 28664) * $signed(input_fmap_219[7:0]) +
	( 15'sd 8843) * $signed(input_fmap_220[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15394) * $signed(input_fmap_222[7:0]) +
	( 14'sd 6985) * $signed(input_fmap_223[7:0]) +
	( 10'sd 267) * $signed(input_fmap_224[7:0]) +
	( 16'sd 23460) * $signed(input_fmap_225[7:0]) +
	( 13'sd 2866) * $signed(input_fmap_226[7:0]) +
	( 16'sd 30815) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25883) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6275) * $signed(input_fmap_229[7:0]) +
	( 16'sd 22359) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7070) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9638) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_233[7:0]) +
	( 15'sd 12330) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29446) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30597) * $signed(input_fmap_236[7:0]) +
	( 15'sd 8777) * $signed(input_fmap_237[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_238[7:0]) +
	( 9'sd 235) * $signed(input_fmap_239[7:0]) +
	( 15'sd 12321) * $signed(input_fmap_240[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_241[7:0]) +
	( 15'sd 14349) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10277) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28301) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2919) * $signed(input_fmap_245[7:0]) +
	( 16'sd 24079) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21853) * $signed(input_fmap_247[7:0]) +
	( 16'sd 17045) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9208) * $signed(input_fmap_249[7:0]) +
	( 15'sd 15917) * $signed(input_fmap_250[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6665) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25101) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2085) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23254) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_37;
assign conv_mac_37 = 
	( 16'sd 32031) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24834) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9118) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18573) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14946) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5387) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4220) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18682) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5195) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23611) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17393) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12898) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5447) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8551) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24123) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14160) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4898) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16936) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26937) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8924) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13248) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8583) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16775) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16732) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15588) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10982) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22348) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15760) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32571) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17666) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29932) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19663) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8436) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14891) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12451) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32041) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18676) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20085) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22522) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13853) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27251) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16522) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29309) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26108) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17438) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27088) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9319) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6731) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10045) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5180) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18227) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4761) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5308) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20107) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20651) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13994) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10152) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31261) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10263) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18415) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25926) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1171) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30224) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26131) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14533) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31118) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25742) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28759) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30455) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3928) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4435) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10632) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19776) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15246) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25214) * $signed(input_fmap_87[7:0]) +
	( 9'sd 225) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19673) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13399) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19883) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32370) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29739) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22874) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31464) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1313) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29157) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2450) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19379) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10457) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31492) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8792) * $signed(input_fmap_102[7:0]) +
	( 10'sd 370) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16158) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27534) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2787) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4397) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1150) * $signed(input_fmap_108[7:0]) +
	( 11'sd 797) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8893) * $signed(input_fmap_110[7:0]) +
	( 11'sd 786) * $signed(input_fmap_111[7:0]) +
	( 10'sd 431) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31992) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2392) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16595) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12266) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15159) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4652) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32416) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9674) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19590) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12326) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31067) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18896) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28769) * $signed(input_fmap_127[7:0]) +
	( 15'sd 14101) * $signed(input_fmap_128[7:0]) +
	( 16'sd 25693) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_130[7:0]) +
	( 15'sd 8767) * $signed(input_fmap_131[7:0]) +
	( 16'sd 32392) * $signed(input_fmap_132[7:0]) +
	( 16'sd 17553) * $signed(input_fmap_133[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_134[7:0]) +
	( 14'sd 7858) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8455) * $signed(input_fmap_136[7:0]) +
	( 16'sd 30930) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19507) * $signed(input_fmap_138[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_139[7:0]) +
	( 15'sd 12212) * $signed(input_fmap_140[7:0]) +
	( 14'sd 4904) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4901) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9817) * $signed(input_fmap_144[7:0]) +
	( 15'sd 12231) * $signed(input_fmap_145[7:0]) +
	( 10'sd 311) * $signed(input_fmap_146[7:0]) +
	( 16'sd 28080) * $signed(input_fmap_147[7:0]) +
	( 15'sd 15534) * $signed(input_fmap_148[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_149[7:0]) +
	( 15'sd 16005) * $signed(input_fmap_150[7:0]) +
	( 16'sd 20662) * $signed(input_fmap_151[7:0]) +
	( 15'sd 13976) * $signed(input_fmap_152[7:0]) +
	( 15'sd 13444) * $signed(input_fmap_153[7:0]) +
	( 16'sd 28283) * $signed(input_fmap_154[7:0]) +
	( 16'sd 16767) * $signed(input_fmap_155[7:0]) +
	( 16'sd 32621) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20402) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11754) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32617) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18699) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22892) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30485) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30259) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6780) * $signed(input_fmap_164[7:0]) +
	( 7'sd 33) * $signed(input_fmap_165[7:0]) +
	( 14'sd 6826) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_167[7:0]) +
	( 16'sd 30827) * $signed(input_fmap_168[7:0]) +
	( 15'sd 9556) * $signed(input_fmap_169[7:0]) +
	( 16'sd 29590) * $signed(input_fmap_170[7:0]) +
	( 16'sd 22855) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6490) * $signed(input_fmap_172[7:0]) +
	( 16'sd 21600) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11276) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28348) * $signed(input_fmap_175[7:0]) +
	( 10'sd 443) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6312) * $signed(input_fmap_177[7:0]) +
	( 16'sd 20465) * $signed(input_fmap_178[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4111) * $signed(input_fmap_180[7:0]) +
	( 10'sd 444) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29818) * $signed(input_fmap_182[7:0]) +
	( 15'sd 10935) * $signed(input_fmap_183[7:0]) +
	( 16'sd 16860) * $signed(input_fmap_184[7:0]) +
	( 15'sd 12975) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2217) * $signed(input_fmap_186[7:0]) +
	( 15'sd 8198) * $signed(input_fmap_187[7:0]) +
	( 16'sd 25759) * $signed(input_fmap_188[7:0]) +
	( 16'sd 22748) * $signed(input_fmap_189[7:0]) +
	( 16'sd 19593) * $signed(input_fmap_190[7:0]) +
	( 16'sd 25013) * $signed(input_fmap_191[7:0]) +
	( 16'sd 18847) * $signed(input_fmap_192[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_193[7:0]) +
	( 16'sd 31978) * $signed(input_fmap_194[7:0]) +
	( 14'sd 4260) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24220) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_198[7:0]) +
	( 16'sd 31059) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26567) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6700) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5934) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21180) * $signed(input_fmap_203[7:0]) +
	( 14'sd 7091) * $signed(input_fmap_204[7:0]) +
	( 14'sd 4861) * $signed(input_fmap_205[7:0]) +
	( 13'sd 4042) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28661) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11695) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26720) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3794) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6178) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18051) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29474) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30658) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29708) * $signed(input_fmap_215[7:0]) +
	( 16'sd 25037) * $signed(input_fmap_216[7:0]) +
	( 16'sd 29867) * $signed(input_fmap_217[7:0]) +
	( 16'sd 24690) * $signed(input_fmap_218[7:0]) +
	( 16'sd 28209) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19531) * $signed(input_fmap_220[7:0]) +
	( 16'sd 20396) * $signed(input_fmap_221[7:0]) +
	( 16'sd 17399) * $signed(input_fmap_222[7:0]) +
	( 14'sd 8134) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27155) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27755) * $signed(input_fmap_225[7:0]) +
	( 15'sd 9570) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6382) * $signed(input_fmap_227[7:0]) +
	( 16'sd 30701) * $signed(input_fmap_228[7:0]) +
	( 16'sd 32003) * $signed(input_fmap_229[7:0]) +
	( 10'sd 423) * $signed(input_fmap_230[7:0]) +
	( 16'sd 23789) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20019) * $signed(input_fmap_232[7:0]) +
	( 15'sd 9197) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19266) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14369) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_236[7:0]) +
	( 15'sd 9425) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3956) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20758) * $signed(input_fmap_239[7:0]) +
	( 15'sd 11780) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25275) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5806) * $signed(input_fmap_242[7:0]) +
	( 14'sd 4965) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30680) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6074) * $signed(input_fmap_245[7:0]) +
	( 15'sd 13165) * $signed(input_fmap_246[7:0]) +
	( 15'sd 10729) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_249[7:0]) +
	( 15'sd 14737) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7277) * $signed(input_fmap_251[7:0]) +
	( 13'sd 3635) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_253[7:0]) +
	( 9'sd 228) * $signed(input_fmap_254[7:0]) +
	( 12'sd 1194) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_38;
assign conv_mac_38 = 
	( 14'sd 4715) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12365) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21263) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23375) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3225) * $signed(input_fmap_5[7:0]) +
	( 14'sd 8144) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22587) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29706) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20921) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25382) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12511) * $signed(input_fmap_12[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14222) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5689) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17786) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5621) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18789) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20919) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4463) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30367) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21838) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3425) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30630) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25021) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14394) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32650) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31920) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11288) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29448) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4579) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2374) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8737) * $signed(input_fmap_34[7:0]) +
	( 8'sd 66) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2128) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16645) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6001) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5541) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30034) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13782) * $signed(input_fmap_44[7:0]) +
	( 10'sd 506) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8518) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21287) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14076) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11919) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4312) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4533) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10300) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6912) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9111) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8461) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20054) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10823) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27386) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10660) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13745) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19007) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32518) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6759) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6669) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29634) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10185) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15750) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15149) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1470) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28537) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22587) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15276) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19786) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1438) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16356) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19235) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5933) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5442) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25507) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18824) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31447) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8380) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26214) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14336) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22991) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30099) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13143) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23534) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29037) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7511) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20514) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30851) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21590) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31440) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25887) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31157) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23789) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26661) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8691) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4405) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27406) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1776) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16083) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12276) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19952) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30302) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29580) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24697) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11654) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22672) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4693) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28319) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20388) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11127) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22048) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27090) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7216) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21771) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13480) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19084) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6247) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19974) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18624) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31321) * $signed(input_fmap_133[7:0]) +
	( 15'sd 15910) * $signed(input_fmap_134[7:0]) +
	( 14'sd 4432) * $signed(input_fmap_135[7:0]) +
	( 16'sd 24944) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11764) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27991) * $signed(input_fmap_138[7:0]) +
	( 15'sd 13638) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1600) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22462) * $signed(input_fmap_141[7:0]) +
	( 14'sd 4690) * $signed(input_fmap_142[7:0]) +
	( 16'sd 32616) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2346) * $signed(input_fmap_144[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_145[7:0]) +
	( 16'sd 23975) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29124) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6895) * $signed(input_fmap_148[7:0]) +
	( 14'sd 6336) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5191) * $signed(input_fmap_150[7:0]) +
	( 16'sd 27380) * $signed(input_fmap_151[7:0]) +
	( 16'sd 19853) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23147) * $signed(input_fmap_153[7:0]) +
	( 16'sd 29485) * $signed(input_fmap_154[7:0]) +
	( 13'sd 2306) * $signed(input_fmap_155[7:0]) +
	( 16'sd 23917) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25920) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11660) * $signed(input_fmap_158[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_159[7:0]) +
	( 9'sd 254) * $signed(input_fmap_160[7:0]) +
	( 10'sd 331) * $signed(input_fmap_161[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22224) * $signed(input_fmap_163[7:0]) +
	( 16'sd 17736) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11140) * $signed(input_fmap_165[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_166[7:0]) +
	( 11'sd 649) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_168[7:0]) +
	( 15'sd 16352) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17038) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20866) * $signed(input_fmap_171[7:0]) +
	( 11'sd 955) * $signed(input_fmap_172[7:0]) +
	( 16'sd 22615) * $signed(input_fmap_173[7:0]) +
	( 12'sd 1672) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7035) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10321) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15610) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14362) * $signed(input_fmap_178[7:0]) +
	( 16'sd 21425) * $signed(input_fmap_179[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3582) * $signed(input_fmap_181[7:0]) +
	( 14'sd 7088) * $signed(input_fmap_182[7:0]) +
	( 15'sd 15772) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31328) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17256) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3884) * $signed(input_fmap_186[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29946) * $signed(input_fmap_188[7:0]) +
	( 16'sd 31746) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3833) * $signed(input_fmap_191[7:0]) +
	( 12'sd 1773) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10451) * $signed(input_fmap_193[7:0]) +
	( 15'sd 10026) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29074) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7942) * $signed(input_fmap_196[7:0]) +
	( 14'sd 7729) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19434) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12837) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2322) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12048) * $signed(input_fmap_203[7:0]) +
	( 14'sd 7676) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12310) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20053) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13139) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25361) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6187) * $signed(input_fmap_211[7:0]) +
	( 13'sd 2233) * $signed(input_fmap_212[7:0]) +
	( 16'sd 16851) * $signed(input_fmap_213[7:0]) +
	( 15'sd 12170) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1436) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19256) * $signed(input_fmap_216[7:0]) +
	( 14'sd 5861) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5992) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5761) * $signed(input_fmap_219[7:0]) +
	( 14'sd 5514) * $signed(input_fmap_220[7:0]) +
	( 16'sd 16448) * $signed(input_fmap_221[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17090) * $signed(input_fmap_223[7:0]) +
	( 14'sd 5558) * $signed(input_fmap_224[7:0]) +
	( 16'sd 25281) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27441) * $signed(input_fmap_226[7:0]) +
	( 16'sd 19530) * $signed(input_fmap_227[7:0]) +
	( 16'sd 30636) * $signed(input_fmap_228[7:0]) +
	( 15'sd 15584) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6500) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3903) * $signed(input_fmap_231[7:0]) +
	( 16'sd 27520) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18803) * $signed(input_fmap_233[7:0]) +
	( 13'sd 2740) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26752) * $signed(input_fmap_235[7:0]) +
	( 15'sd 9328) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19315) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13881) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20506) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31652) * $signed(input_fmap_240[7:0]) +
	( 8'sd 67) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23590) * $signed(input_fmap_242[7:0]) +
	( 16'sd 32555) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12884) * $signed(input_fmap_244[7:0]) +
	( 16'sd 26031) * $signed(input_fmap_245[7:0]) +
	( 16'sd 32331) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9368) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10566) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30078) * $signed(input_fmap_249[7:0]) +
	( 16'sd 21572) * $signed(input_fmap_250[7:0]) +
	( 13'sd 3304) * $signed(input_fmap_251[7:0]) +
	( 8'sd 89) * $signed(input_fmap_252[7:0]) +
	( 14'sd 7189) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31054) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24257) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_39;
assign conv_mac_39 = 
	( 15'sd 9362) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22675) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12400) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21472) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27822) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20375) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23645) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18399) * $signed(input_fmap_8[7:0]) +
	( 10'sd 357) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3567) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5701) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2999) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16396) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26259) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14395) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11597) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32054) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23267) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23932) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7517) * $signed(input_fmap_22[7:0]) +
	( 12'sd 2013) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5647) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25088) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21859) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25123) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5000) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22182) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9508) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27175) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27517) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15021) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6502) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27795) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15644) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5777) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10766) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8586) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18357) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3156) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29244) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17987) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8993) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26839) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32149) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18847) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29087) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32244) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7036) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29475) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15468) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24502) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23709) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25269) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18897) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24012) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13897) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27592) * $signed(input_fmap_65[7:0]) +
	( 11'sd 615) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23770) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21491) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24986) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10816) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28041) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14395) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25910) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1699) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32295) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27103) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24941) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9089) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25231) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28359) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26119) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14458) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23633) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10603) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15763) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2884) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22364) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30576) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19746) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10637) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19819) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9993) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21432) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22816) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19232) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28284) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1299) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17409) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7723) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1249) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3103) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20983) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26127) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20747) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5221) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6093) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28403) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29261) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10725) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21785) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2969) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22924) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8624) * $signed(input_fmap_118[7:0]) +
	( 11'sd 939) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3861) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3844) * $signed(input_fmap_121[7:0]) +
	( 11'sd 627) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22194) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25666) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31355) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24648) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1643) * $signed(input_fmap_127[7:0]) +
	( 16'sd 19123) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24442) * $signed(input_fmap_129[7:0]) +
	( 15'sd 11090) * $signed(input_fmap_130[7:0]) +
	( 14'sd 7852) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11606) * $signed(input_fmap_132[7:0]) +
	( 15'sd 13498) * $signed(input_fmap_133[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_134[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_135[7:0]) +
	( 13'sd 3310) * $signed(input_fmap_136[7:0]) +
	( 16'sd 16389) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17551) * $signed(input_fmap_138[7:0]) +
	( 15'sd 9388) * $signed(input_fmap_139[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_140[7:0]) +
	( 16'sd 16454) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31845) * $signed(input_fmap_142[7:0]) +
	( 16'sd 30689) * $signed(input_fmap_143[7:0]) +
	( 16'sd 16933) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27616) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14783) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29930) * $signed(input_fmap_147[7:0]) +
	( 16'sd 32531) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_149[7:0]) +
	( 15'sd 10830) * $signed(input_fmap_150[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27008) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24667) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28833) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7858) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11424) * $signed(input_fmap_157[7:0]) +
	( 16'sd 32728) * $signed(input_fmap_158[7:0]) +
	( 15'sd 11146) * $signed(input_fmap_159[7:0]) +
	( 15'sd 9709) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28606) * $signed(input_fmap_161[7:0]) +
	( 15'sd 16096) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3703) * $signed(input_fmap_163[7:0]) +
	( 15'sd 14149) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28799) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3739) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7561) * $signed(input_fmap_167[7:0]) +
	( 15'sd 10392) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21964) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2550) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14968) * $signed(input_fmap_172[7:0]) +
	( 15'sd 13610) * $signed(input_fmap_173[7:0]) +
	( 16'sd 18603) * $signed(input_fmap_174[7:0]) +
	( 16'sd 24645) * $signed(input_fmap_175[7:0]) +
	( 14'sd 6346) * $signed(input_fmap_176[7:0]) +
	( 15'sd 16294) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27048) * $signed(input_fmap_178[7:0]) +
	( 16'sd 19690) * $signed(input_fmap_179[7:0]) +
	( 16'sd 17226) * $signed(input_fmap_180[7:0]) +
	( 10'sd 348) * $signed(input_fmap_181[7:0]) +
	( 15'sd 15431) * $signed(input_fmap_182[7:0]) +
	( 15'sd 10359) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26999) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22849) * $signed(input_fmap_185[7:0]) +
	( 15'sd 11861) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_187[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_188[7:0]) +
	( 16'sd 22926) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20038) * $signed(input_fmap_190[7:0]) +
	( 12'sd 1987) * $signed(input_fmap_191[7:0]) +
	( 15'sd 10301) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_193[7:0]) +
	( 15'sd 10586) * $signed(input_fmap_194[7:0]) +
	( 16'sd 20342) * $signed(input_fmap_195[7:0]) +
	( 13'sd 4010) * $signed(input_fmap_196[7:0]) +
	( 15'sd 12953) * $signed(input_fmap_197[7:0]) +
	( 16'sd 31801) * $signed(input_fmap_198[7:0]) +
	( 13'sd 2918) * $signed(input_fmap_199[7:0]) +
	( 16'sd 32233) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1460) * $signed(input_fmap_201[7:0]) +
	( 16'sd 28271) * $signed(input_fmap_202[7:0]) +
	( 15'sd 10011) * $signed(input_fmap_203[7:0]) +
	( 16'sd 22471) * $signed(input_fmap_204[7:0]) +
	( 16'sd 20710) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12827) * $signed(input_fmap_206[7:0]) +
	( 15'sd 16118) * $signed(input_fmap_207[7:0]) +
	( 16'sd 27982) * $signed(input_fmap_208[7:0]) +
	( 16'sd 29752) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11165) * $signed(input_fmap_210[7:0]) +
	( 15'sd 14095) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24425) * $signed(input_fmap_212[7:0]) +
	( 15'sd 13352) * $signed(input_fmap_213[7:0]) +
	( 14'sd 4653) * $signed(input_fmap_214[7:0]) +
	( 16'sd 26782) * $signed(input_fmap_215[7:0]) +
	( 16'sd 31626) * $signed(input_fmap_216[7:0]) +
	( 14'sd 4305) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28093) * $signed(input_fmap_218[7:0]) +
	( 11'sd 891) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25137) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12214) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3900) * $signed(input_fmap_222[7:0]) +
	( 15'sd 16131) * $signed(input_fmap_223[7:0]) +
	( 14'sd 4694) * $signed(input_fmap_224[7:0]) +
	( 16'sd 30436) * $signed(input_fmap_225[7:0]) +
	( 16'sd 28400) * $signed(input_fmap_226[7:0]) +
	( 16'sd 17560) * $signed(input_fmap_227[7:0]) +
	( 14'sd 5496) * $signed(input_fmap_228[7:0]) +
	( 16'sd 25556) * $signed(input_fmap_229[7:0]) +
	( 16'sd 23391) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25892) * $signed(input_fmap_231[7:0]) +
	( 14'sd 6823) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21915) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18386) * $signed(input_fmap_234[7:0]) +
	( 15'sd 8567) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10979) * $signed(input_fmap_236[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_237[7:0]) +
	( 14'sd 4239) * $signed(input_fmap_238[7:0]) +
	( 14'sd 6083) * $signed(input_fmap_239[7:0]) +
	( 13'sd 2350) * $signed(input_fmap_240[7:0]) +
	( 14'sd 6183) * $signed(input_fmap_241[7:0]) +
	( 16'sd 30916) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2402) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12758) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_245[7:0]) +
	( 14'sd 6092) * $signed(input_fmap_246[7:0]) +
	( 12'sd 1226) * $signed(input_fmap_247[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28745) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32447) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18425) * $signed(input_fmap_251[7:0]) +
	( 16'sd 19039) * $signed(input_fmap_252[7:0]) +
	( 16'sd 31429) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26569) * $signed(input_fmap_254[7:0]) +
	( 15'sd 15183) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_40;
assign conv_mac_40 = 
	( 15'sd 13633) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28377) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26572) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25899) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11864) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22923) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4448) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28946) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13267) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13613) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25933) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20210) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13946) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18134) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12696) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15724) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32445) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16499) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22895) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22664) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8467) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22417) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15116) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8633) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21311) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21363) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26777) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30118) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17286) * $signed(input_fmap_35[7:0]) +
	( 11'sd 819) * $signed(input_fmap_36[7:0]) +
	( 11'sd 783) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26942) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4902) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32213) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25240) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31101) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4717) * $signed(input_fmap_43[7:0]) +
	( 11'sd 973) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25944) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12082) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26057) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21801) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1501) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30780) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29455) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2939) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30299) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12187) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25484) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9487) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9569) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8630) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28596) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19046) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29738) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21931) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18632) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31847) * $signed(input_fmap_65[7:0]) +
	( 9'sd 209) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21123) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3250) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17639) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30366) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13902) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21063) * $signed(input_fmap_73[7:0]) +
	( 9'sd 252) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3333) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27060) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18134) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22920) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7374) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24999) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13005) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17152) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30081) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19568) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9894) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2253) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8953) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10278) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18595) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_92[7:0]) +
	( 11'sd 793) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12468) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3138) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30191) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9624) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3603) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20571) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14142) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19261) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6016) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31965) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28210) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1670) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3586) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21873) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16078) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20515) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29083) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25837) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23259) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1339) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6256) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8673) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24946) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23982) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30461) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8192) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20497) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18027) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32511) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14487) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15225) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29668) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8916) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27231) * $signed(input_fmap_129[7:0]) +
	( 15'sd 8662) * $signed(input_fmap_130[7:0]) +
	( 13'sd 2945) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18191) * $signed(input_fmap_132[7:0]) +
	( 16'sd 32447) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19819) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21447) * $signed(input_fmap_136[7:0]) +
	( 16'sd 29922) * $signed(input_fmap_137[7:0]) +
	( 15'sd 14239) * $signed(input_fmap_138[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_139[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_140[7:0]) +
	( 12'sd 1118) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31626) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4315) * $signed(input_fmap_143[7:0]) +
	( 16'sd 17994) * $signed(input_fmap_144[7:0]) +
	( 16'sd 29060) * $signed(input_fmap_145[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_146[7:0]) +
	( 10'sd 473) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21053) * $signed(input_fmap_148[7:0]) +
	( 15'sd 9625) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21677) * $signed(input_fmap_150[7:0]) +
	( 15'sd 9063) * $signed(input_fmap_151[7:0]) +
	( 16'sd 19178) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12687) * $signed(input_fmap_153[7:0]) +
	( 15'sd 9914) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23813) * $signed(input_fmap_155[7:0]) +
	( 15'sd 8379) * $signed(input_fmap_156[7:0]) +
	( 16'sd 26330) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4714) * $signed(input_fmap_158[7:0]) +
	( 15'sd 9932) * $signed(input_fmap_159[7:0]) +
	( 15'sd 15038) * $signed(input_fmap_160[7:0]) +
	( 15'sd 14624) * $signed(input_fmap_161[7:0]) +
	( 14'sd 5461) * $signed(input_fmap_162[7:0]) +
	( 15'sd 14039) * $signed(input_fmap_163[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_164[7:0]) +
	( 15'sd 16052) * $signed(input_fmap_165[7:0]) +
	( 16'sd 27210) * $signed(input_fmap_166[7:0]) +
	( 15'sd 15071) * $signed(input_fmap_167[7:0]) +
	( 13'sd 2374) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3877) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28092) * $signed(input_fmap_170[7:0]) +
	( 16'sd 29706) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_172[7:0]) +
	( 16'sd 24639) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10046) * $signed(input_fmap_174[7:0]) +
	( 16'sd 27469) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27400) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22028) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17861) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5861) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27674) * $signed(input_fmap_180[7:0]) +
	( 16'sd 29183) * $signed(input_fmap_181[7:0]) +
	( 16'sd 23070) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_183[7:0]) +
	( 14'sd 6015) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26805) * $signed(input_fmap_186[7:0]) +
	( 16'sd 32462) * $signed(input_fmap_187[7:0]) +
	( 14'sd 7792) * $signed(input_fmap_188[7:0]) +
	( 15'sd 13454) * $signed(input_fmap_189[7:0]) +
	( 16'sd 16629) * $signed(input_fmap_190[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28014) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19201) * $signed(input_fmap_193[7:0]) +
	( 12'sd 1258) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29451) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5101) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19427) * $signed(input_fmap_197[7:0]) +
	( 16'sd 25172) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10972) * $signed(input_fmap_199[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_200[7:0]) +
	( 16'sd 17499) * $signed(input_fmap_201[7:0]) +
	( 15'sd 12201) * $signed(input_fmap_202[7:0]) +
	( 16'sd 22983) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5457) * $signed(input_fmap_204[7:0]) +
	( 13'sd 3377) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3236) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4315) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11482) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11989) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26854) * $signed(input_fmap_211[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_213[7:0]) +
	( 16'sd 21745) * $signed(input_fmap_214[7:0]) +
	( 13'sd 3972) * $signed(input_fmap_215[7:0]) +
	( 16'sd 29882) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_217[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21969) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31400) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13706) * $signed(input_fmap_221[7:0]) +
	( 16'sd 26771) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14170) * $signed(input_fmap_223[7:0]) +
	( 16'sd 31033) * $signed(input_fmap_224[7:0]) +
	( 16'sd 31455) * $signed(input_fmap_225[7:0]) +
	( 15'sd 12417) * $signed(input_fmap_226[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_227[7:0]) +
	( 14'sd 5340) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10006) * $signed(input_fmap_229[7:0]) +
	( 11'sd 532) * $signed(input_fmap_230[7:0]) +
	( 15'sd 15780) * $signed(input_fmap_231[7:0]) +
	( 16'sd 27123) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27441) * $signed(input_fmap_233[7:0]) +
	( 16'sd 24934) * $signed(input_fmap_234[7:0]) +
	( 14'sd 4913) * $signed(input_fmap_235[7:0]) +
	( 15'sd 13647) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20474) * $signed(input_fmap_237[7:0]) +
	( 16'sd 18481) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19296) * $signed(input_fmap_239[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18451) * $signed(input_fmap_241[7:0]) +
	( 16'sd 16744) * $signed(input_fmap_242[7:0]) +
	( 16'sd 24417) * $signed(input_fmap_243[7:0]) +
	( 15'sd 15247) * $signed(input_fmap_244[7:0]) +
	( 15'sd 9059) * $signed(input_fmap_245[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17209) * $signed(input_fmap_247[7:0]) +
	( 16'sd 17399) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25406) * $signed(input_fmap_249[7:0]) +
	( 15'sd 13842) * $signed(input_fmap_250[7:0]) +
	( 16'sd 31475) * $signed(input_fmap_251[7:0]) +
	( 16'sd 24685) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9379) * $signed(input_fmap_254[7:0]) +
	( 15'sd 9365) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_41;
assign conv_mac_41 = 
	( 16'sd 30891) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6619) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22097) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16874) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25731) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29012) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5951) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20924) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13515) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30972) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22697) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1070) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30292) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15902) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32516) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3290) * $signed(input_fmap_16[7:0]) +
	( 9'sd 139) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21417) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18630) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26489) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18243) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30928) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6755) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11602) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2174) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2830) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2487) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5006) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24410) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22368) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14996) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8274) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27496) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13400) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21449) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19041) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12315) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3835) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22857) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27295) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13416) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16096) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2138) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7046) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31851) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11661) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1916) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15960) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9196) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12152) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10295) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3681) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9066) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30275) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17077) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3794) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13980) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17312) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14525) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6734) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12368) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1038) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13948) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32716) * $signed(input_fmap_69[7:0]) +
	( 9'sd 205) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15967) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13711) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29582) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20744) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16036) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28436) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2597) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23126) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30091) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3691) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1242) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6337) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17862) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1211) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16020) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4689) * $signed(input_fmap_86[7:0]) +
	( 13'sd 4059) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30781) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15741) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7592) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8973) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7010) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2088) * $signed(input_fmap_93[7:0]) +
	( 13'sd 4023) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3105) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17984) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20892) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32763) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10027) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11968) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12851) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29933) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24046) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15556) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20588) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5559) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8337) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23367) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17905) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8480) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21926) * $signed(input_fmap_112[7:0]) +
	( 11'sd 1014) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13993) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2067) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8052) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15209) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24096) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29650) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20293) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19572) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12184) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1167) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23030) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1256) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15506) * $signed(input_fmap_128[7:0]) +
	( 16'sd 18952) * $signed(input_fmap_129[7:0]) +
	( 16'sd 23322) * $signed(input_fmap_130[7:0]) +
	( 16'sd 27901) * $signed(input_fmap_131[7:0]) +
	( 14'sd 6189) * $signed(input_fmap_132[7:0]) +
	( 16'sd 30038) * $signed(input_fmap_133[7:0]) +
	( 16'sd 28057) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26909) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4962) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6691) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27611) * $signed(input_fmap_138[7:0]) +
	( 16'sd 23326) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30211) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24594) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28438) * $signed(input_fmap_142[7:0]) +
	( 16'sd 21463) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28550) * $signed(input_fmap_144[7:0]) +
	( 15'sd 14720) * $signed(input_fmap_145[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24914) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3296) * $signed(input_fmap_148[7:0]) +
	( 15'sd 14659) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25044) * $signed(input_fmap_150[7:0]) +
	( 16'sd 27677) * $signed(input_fmap_151[7:0]) +
	( 14'sd 4891) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3692) * $signed(input_fmap_153[7:0]) +
	( 16'sd 20936) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10944) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13859) * $signed(input_fmap_156[7:0]) +
	( 16'sd 26597) * $signed(input_fmap_157[7:0]) +
	( 15'sd 16105) * $signed(input_fmap_158[7:0]) +
	( 16'sd 22798) * $signed(input_fmap_159[7:0]) +
	( 16'sd 23912) * $signed(input_fmap_160[7:0]) +
	( 16'sd 25552) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27951) * $signed(input_fmap_162[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_163[7:0]) +
	( 16'sd 27310) * $signed(input_fmap_164[7:0]) +
	( 16'sd 31632) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4845) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9797) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1214) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12914) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23110) * $signed(input_fmap_170[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_171[7:0]) +
	( 15'sd 13739) * $signed(input_fmap_172[7:0]) +
	( 16'sd 30598) * $signed(input_fmap_173[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_174[7:0]) +
	( 15'sd 12504) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10845) * $signed(input_fmap_176[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_177[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28587) * $signed(input_fmap_180[7:0]) +
	( 14'sd 8128) * $signed(input_fmap_181[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25567) * $signed(input_fmap_183[7:0]) +
	( 16'sd 19385) * $signed(input_fmap_184[7:0]) +
	( 15'sd 12023) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9535) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4906) * $signed(input_fmap_187[7:0]) +
	( 16'sd 26361) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30041) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9369) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20043) * $signed(input_fmap_191[7:0]) +
	( 16'sd 17703) * $signed(input_fmap_192[7:0]) +
	( 16'sd 18798) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_194[7:0]) +
	( 15'sd 10333) * $signed(input_fmap_195[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26788) * $signed(input_fmap_197[7:0]) +
	( 15'sd 12097) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28235) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8910) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15648) * $signed(input_fmap_201[7:0]) +
	( 16'sd 30850) * $signed(input_fmap_202[7:0]) +
	( 11'sd 667) * $signed(input_fmap_203[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1191) * $signed(input_fmap_205[7:0]) +
	( 15'sd 11720) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28133) * $signed(input_fmap_207[7:0]) +
	( 12'sd 1343) * $signed(input_fmap_208[7:0]) +
	( 12'sd 1566) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15210) * $signed(input_fmap_210[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_211[7:0]) +
	( 14'sd 4866) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11651) * $signed(input_fmap_213[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2931) * $signed(input_fmap_215[7:0]) +
	( 11'sd 799) * $signed(input_fmap_216[7:0]) +
	( 15'sd 11515) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22569) * $signed(input_fmap_218[7:0]) +
	( 14'sd 4454) * $signed(input_fmap_219[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6487) * $signed(input_fmap_221[7:0]) +
	( 15'sd 9874) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2843) * $signed(input_fmap_223[7:0]) +
	( 16'sd 32127) * $signed(input_fmap_224[7:0]) +
	( 15'sd 9096) * $signed(input_fmap_225[7:0]) +
	( 16'sd 19559) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13990) * $signed(input_fmap_227[7:0]) +
	( 16'sd 23211) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8196) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_230[7:0]) +
	( 16'sd 26843) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12069) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1919) * $signed(input_fmap_233[7:0]) +
	( 16'sd 24310) * $signed(input_fmap_234[7:0]) +
	( 15'sd 9218) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_236[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22117) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1431) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25096) * $signed(input_fmap_241[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23388) * $signed(input_fmap_243[7:0]) +
	( 16'sd 32566) * $signed(input_fmap_244[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1097) * $signed(input_fmap_246[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_247[7:0]) +
	( 14'sd 5256) * $signed(input_fmap_248[7:0]) +
	( 10'sd 306) * $signed(input_fmap_249[7:0]) +
	( 2'sd 1) * $signed(input_fmap_250[7:0]) +
	( 12'sd 1718) * $signed(input_fmap_251[7:0]) +
	( 9'sd 253) * $signed(input_fmap_252[7:0]) +
	( 15'sd 10802) * $signed(input_fmap_253[7:0]) +
	( 16'sd 22968) * $signed(input_fmap_254[7:0]) +
	( 15'sd 12526) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_42;
assign conv_mac_42 = 
	( 16'sd 32378) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5885) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17155) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11339) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26245) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17462) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8441) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21453) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30785) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29889) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4289) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14482) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12682) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14994) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17645) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13278) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13939) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15543) * $signed(input_fmap_19[7:0]) +
	( 10'sd 311) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30067) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24202) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28238) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31998) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1655) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21332) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14228) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18429) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16551) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20948) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29176) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1988) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25165) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12801) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9064) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26040) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20481) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2640) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22202) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13183) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13868) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25686) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28320) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14145) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30012) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1127) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16565) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12304) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30799) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30645) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12359) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32317) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12277) * $signed(input_fmap_55[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28798) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27310) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11201) * $signed(input_fmap_60[7:0]) +
	( 9'sd 141) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25549) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11061) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27624) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3558) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16564) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22267) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8358) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4380) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18658) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25506) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13201) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22435) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13049) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17623) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10080) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21605) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32645) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10453) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13603) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6768) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19851) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19967) * $signed(input_fmap_86[7:0]) +
	( 11'sd 861) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14144) * $signed(input_fmap_88[7:0]) +
	( 11'sd 756) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29843) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29197) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30995) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2993) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24880) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10038) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29431) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14121) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25252) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25630) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19803) * $signed(input_fmap_100[7:0]) +
	( 10'sd 483) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21040) * $signed(input_fmap_102[7:0]) +
	( 9'sd 224) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6020) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4568) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7268) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7288) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16193) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21859) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27514) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28836) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30192) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32703) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8930) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8017) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6265) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22206) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18433) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31547) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26579) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11820) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18732) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9648) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25034) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25413) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26457) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31701) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1047) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30178) * $signed(input_fmap_130[7:0]) +
	( 15'sd 10496) * $signed(input_fmap_131[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_132[7:0]) +
	( 10'sd 410) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21426) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32144) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17460) * $signed(input_fmap_136[7:0]) +
	( 14'sd 8073) * $signed(input_fmap_137[7:0]) +
	( 14'sd 5316) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_139[7:0]) +
	( 13'sd 2278) * $signed(input_fmap_140[7:0]) +
	( 15'sd 11033) * $signed(input_fmap_141[7:0]) +
	( 14'sd 5649) * $signed(input_fmap_142[7:0]) +
	( 15'sd 15082) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22477) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25176) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27764) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8298) * $signed(input_fmap_147[7:0]) +
	( 16'sd 24213) * $signed(input_fmap_148[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_149[7:0]) +
	( 16'sd 32075) * $signed(input_fmap_150[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_151[7:0]) +
	( 14'sd 5709) * $signed(input_fmap_152[7:0]) +
	( 16'sd 22197) * $signed(input_fmap_153[7:0]) +
	( 15'sd 16074) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20478) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29874) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8392) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26439) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31400) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23422) * $signed(input_fmap_161[7:0]) +
	( 11'sd 803) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28640) * $signed(input_fmap_163[7:0]) +
	( 16'sd 22545) * $signed(input_fmap_164[7:0]) +
	( 14'sd 5057) * $signed(input_fmap_165[7:0]) +
	( 14'sd 8022) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20483) * $signed(input_fmap_167[7:0]) +
	( 14'sd 7807) * $signed(input_fmap_168[7:0]) +
	( 12'sd 1125) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14619) * $signed(input_fmap_170[7:0]) +
	( 10'sd 313) * $signed(input_fmap_171[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_172[7:0]) +
	( 8'sd 79) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26450) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7635) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27131) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29032) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10467) * $signed(input_fmap_178[7:0]) +
	( 11'sd 693) * $signed(input_fmap_179[7:0]) +
	( 15'sd 16195) * $signed(input_fmap_180[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_181[7:0]) +
	( 15'sd 14951) * $signed(input_fmap_182[7:0]) +
	( 13'sd 4075) * $signed(input_fmap_183[7:0]) +
	( 16'sd 25477) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6089) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3825) * $signed(input_fmap_186[7:0]) +
	( 15'sd 10908) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21488) * $signed(input_fmap_188[7:0]) +
	( 16'sd 27508) * $signed(input_fmap_189[7:0]) +
	( 15'sd 11853) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17219) * $signed(input_fmap_191[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5214) * $signed(input_fmap_193[7:0]) +
	( 13'sd 2619) * $signed(input_fmap_194[7:0]) +
	( 16'sd 26692) * $signed(input_fmap_195[7:0]) +
	( 13'sd 3899) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19908) * $signed(input_fmap_197[7:0]) +
	( 15'sd 15290) * $signed(input_fmap_198[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21715) * $signed(input_fmap_201[7:0]) +
	( 14'sd 6382) * $signed(input_fmap_202[7:0]) +
	( 16'sd 32383) * $signed(input_fmap_203[7:0]) +
	( 16'sd 20088) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15153) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2290) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1766) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12784) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9550) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_211[7:0]) +
	( 15'sd 16289) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23934) * $signed(input_fmap_213[7:0]) +
	( 15'sd 11013) * $signed(input_fmap_214[7:0]) +
	( 15'sd 14371) * $signed(input_fmap_215[7:0]) +
	( 15'sd 8643) * $signed(input_fmap_216[7:0]) +
	( 15'sd 8850) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_218[7:0]) +
	( 16'sd 24730) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13962) * $signed(input_fmap_220[7:0]) +
	( 16'sd 16787) * $signed(input_fmap_221[7:0]) +
	( 15'sd 8673) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2962) * $signed(input_fmap_223[7:0]) +
	( 16'sd 18459) * $signed(input_fmap_224[7:0]) +
	( 14'sd 6354) * $signed(input_fmap_225[7:0]) +
	( 15'sd 8711) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9908) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26255) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17433) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_230[7:0]) +
	( 16'sd 32239) * $signed(input_fmap_231[7:0]) +
	( 16'sd 27093) * $signed(input_fmap_232[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13351) * $signed(input_fmap_234[7:0]) +
	( 13'sd 2842) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25650) * $signed(input_fmap_236[7:0]) +
	( 16'sd 26553) * $signed(input_fmap_237[7:0]) +
	( 14'sd 8047) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26546) * $signed(input_fmap_239[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_240[7:0]) +
	( 16'sd 17055) * $signed(input_fmap_241[7:0]) +
	( 16'sd 16469) * $signed(input_fmap_242[7:0]) +
	( 16'sd 29384) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2777) * $signed(input_fmap_244[7:0]) +
	( 12'sd 1117) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11484) * $signed(input_fmap_246[7:0]) +
	( 15'sd 10231) * $signed(input_fmap_247[7:0]) +
	( 14'sd 8058) * $signed(input_fmap_248[7:0]) +
	( 14'sd 7258) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17385) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6061) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13749) * $signed(input_fmap_253[7:0]) +
	( 16'sd 30407) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10949) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_43;
assign conv_mac_43 = 
	( 16'sd 19755) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19994) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10222) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17505) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8904) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26405) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23444) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8233) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15945) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15537) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30077) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17007) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11889) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7482) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28216) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17559) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25202) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11138) * $signed(input_fmap_18[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21721) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29185) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12397) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3431) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22169) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17360) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28573) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17204) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15633) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11012) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2194) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19426) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19155) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3258) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22770) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3336) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13244) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20044) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28258) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30028) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24279) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30929) * $signed(input_fmap_46[7:0]) +
	( 10'sd 398) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15640) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14747) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21672) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7981) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16325) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5689) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31615) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30707) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5603) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28173) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11177) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23282) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5044) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20341) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15749) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17998) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14676) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3340) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22532) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26874) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29828) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25147) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20745) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31743) * $signed(input_fmap_74[7:0]) +
	( 11'sd 694) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16635) * $signed(input_fmap_76[7:0]) +
	( 14'sd 8139) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23670) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22556) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6640) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4448) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25679) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13645) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28636) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3156) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4914) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18004) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8606) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31017) * $signed(input_fmap_91[7:0]) +
	( 10'sd 499) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6767) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9199) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12859) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2084) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16907) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1342) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17952) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4918) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19769) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8801) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9713) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32246) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6471) * $signed(input_fmap_105[7:0]) +
	( 8'sd 92) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25252) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20038) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4443) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25602) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19989) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25913) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30843) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9005) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5026) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14116) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27696) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1103) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3096) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2775) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25417) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28240) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30593) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21979) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5335) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4958) * $signed(input_fmap_127[7:0]) +
	( 16'sd 21769) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27330) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12536) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3367) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18221) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16534) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24459) * $signed(input_fmap_134[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_135[7:0]) +
	( 11'sd 967) * $signed(input_fmap_136[7:0]) +
	( 16'sd 19731) * $signed(input_fmap_137[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_138[7:0]) +
	( 16'sd 17368) * $signed(input_fmap_139[7:0]) +
	( 16'sd 25975) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12725) * $signed(input_fmap_141[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_142[7:0]) +
	( 16'sd 29744) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4156) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22477) * $signed(input_fmap_145[7:0]) +
	( 16'sd 32711) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27078) * $signed(input_fmap_147[7:0]) +
	( 15'sd 15282) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25720) * $signed(input_fmap_149[7:0]) +
	( 16'sd 24502) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30645) * $signed(input_fmap_151[7:0]) +
	( 15'sd 15456) * $signed(input_fmap_152[7:0]) +
	( 14'sd 5217) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4548) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7791) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20092) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27035) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25770) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14466) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26792) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1330) * $signed(input_fmap_161[7:0]) +
	( 16'sd 22468) * $signed(input_fmap_162[7:0]) +
	( 12'sd 1300) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24659) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10940) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22316) * $signed(input_fmap_166[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5383) * $signed(input_fmap_168[7:0]) +
	( 11'sd 759) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2270) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16684) * $signed(input_fmap_171[7:0]) +
	( 11'sd 594) * $signed(input_fmap_172[7:0]) +
	( 15'sd 14033) * $signed(input_fmap_173[7:0]) +
	( 16'sd 25561) * $signed(input_fmap_174[7:0]) +
	( 15'sd 9872) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18709) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1819) * $signed(input_fmap_178[7:0]) +
	( 16'sd 17738) * $signed(input_fmap_179[7:0]) +
	( 16'sd 30360) * $signed(input_fmap_180[7:0]) +
	( 15'sd 9901) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5555) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27627) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14030) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1486) * $signed(input_fmap_185[7:0]) +
	( 16'sd 28243) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25069) * $signed(input_fmap_187[7:0]) +
	( 14'sd 7767) * $signed(input_fmap_188[7:0]) +
	( 15'sd 10920) * $signed(input_fmap_189[7:0]) +
	( 16'sd 18417) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5125) * $signed(input_fmap_191[7:0]) +
	( 15'sd 10386) * $signed(input_fmap_192[7:0]) +
	( 16'sd 17592) * $signed(input_fmap_193[7:0]) +
	( 16'sd 22001) * $signed(input_fmap_194[7:0]) +
	( 15'sd 11189) * $signed(input_fmap_195[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_196[7:0]) +
	( 8'sd 89) * $signed(input_fmap_197[7:0]) +
	( 12'sd 1418) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6758) * $signed(input_fmap_199[7:0]) +
	( 16'sd 23501) * $signed(input_fmap_200[7:0]) +
	( 14'sd 5727) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_202[7:0]) +
	( 16'sd 32241) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12908) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31567) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29986) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18789) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22056) * $signed(input_fmap_208[7:0]) +
	( 16'sd 17040) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30477) * $signed(input_fmap_210[7:0]) +
	( 16'sd 29301) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17063) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2479) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_214[7:0]) +
	( 16'sd 27140) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17257) * $signed(input_fmap_216[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_217[7:0]) +
	( 16'sd 16687) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21938) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19880) * $signed(input_fmap_220[7:0]) +
	( 16'sd 29010) * $signed(input_fmap_221[7:0]) +
	( 14'sd 8134) * $signed(input_fmap_222[7:0]) +
	( 13'sd 3168) * $signed(input_fmap_223[7:0]) +
	( 16'sd 32741) * $signed(input_fmap_224[7:0]) +
	( 15'sd 11806) * $signed(input_fmap_225[7:0]) +
	( 15'sd 13476) * $signed(input_fmap_226[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_229[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_230[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_231[7:0]) +
	( 16'sd 16391) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14089) * $signed(input_fmap_233[7:0]) +
	( 16'sd 24576) * $signed(input_fmap_234[7:0]) +
	( 16'sd 25850) * $signed(input_fmap_235[7:0]) +
	( 14'sd 6116) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_237[7:0]) +
	( 16'sd 31006) * $signed(input_fmap_238[7:0]) +
	( 16'sd 30174) * $signed(input_fmap_239[7:0]) +
	( 16'sd 21592) * $signed(input_fmap_240[7:0]) +
	( 15'sd 14216) * $signed(input_fmap_241[7:0]) +
	( 16'sd 24076) * $signed(input_fmap_242[7:0]) +
	( 16'sd 26361) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20801) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24630) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31058) * $signed(input_fmap_246[7:0]) +
	( 13'sd 2912) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32093) * $signed(input_fmap_248[7:0]) +
	( 16'sd 29460) * $signed(input_fmap_249[7:0]) +
	( 14'sd 5729) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15717) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5962) * $signed(input_fmap_252[7:0]) +
	( 15'sd 9012) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19245) * $signed(input_fmap_254[7:0]) +
	( 16'sd 28226) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_44;
assign conv_mac_44 = 
	( 16'sd 16839) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29052) * $signed(input_fmap_2[7:0]) +
	( 11'sd 807) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28827) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19829) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28328) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13968) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11159) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25517) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24294) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15115) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16429) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15822) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10292) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10209) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1522) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16289) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22772) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32471) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17254) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2711) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31837) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8317) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17136) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16153) * $signed(input_fmap_26[7:0]) +
	( 10'sd 401) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13951) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8482) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13724) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30768) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31502) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14719) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21731) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17205) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26873) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31546) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3416) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7329) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16345) * $signed(input_fmap_43[7:0]) +
	( 11'sd 719) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6827) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4366) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7290) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22619) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32277) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11458) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9072) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19896) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29472) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3663) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8214) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4328) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32009) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27371) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28105) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_64[7:0]) +
	( 13'sd 4015) * $signed(input_fmap_65[7:0]) +
	( 8'sd 91) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20701) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17329) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30292) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22903) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11539) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17278) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14693) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11942) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29507) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25853) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16918) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8611) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21827) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9825) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25000) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23984) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1045) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1540) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6735) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15842) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8758) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21460) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27570) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27601) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11575) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21580) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18692) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14548) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29684) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24199) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9232) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18895) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30028) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23547) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1772) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29034) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6446) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5679) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21288) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23170) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14472) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20593) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11915) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24755) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3054) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29903) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3879) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15988) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8910) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23685) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15891) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6075) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13907) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27247) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16415) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16455) * $signed(input_fmap_127[7:0]) +
	( 16'sd 21052) * $signed(input_fmap_128[7:0]) +
	( 15'sd 16346) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18923) * $signed(input_fmap_130[7:0]) +
	( 13'sd 2373) * $signed(input_fmap_131[7:0]) +
	( 16'sd 32022) * $signed(input_fmap_132[7:0]) +
	( 16'sd 19494) * $signed(input_fmap_133[7:0]) +
	( 16'sd 23845) * $signed(input_fmap_134[7:0]) +
	( 16'sd 17157) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12190) * $signed(input_fmap_136[7:0]) +
	( 16'sd 18845) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27955) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3990) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1274) * $signed(input_fmap_140[7:0]) +
	( 15'sd 9492) * $signed(input_fmap_141[7:0]) +
	( 15'sd 12442) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1073) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22417) * $signed(input_fmap_145[7:0]) +
	( 16'sd 32296) * $signed(input_fmap_146[7:0]) +
	( 16'sd 23334) * $signed(input_fmap_147[7:0]) +
	( 15'sd 13943) * $signed(input_fmap_148[7:0]) +
	( 15'sd 13909) * $signed(input_fmap_149[7:0]) +
	( 15'sd 13409) * $signed(input_fmap_150[7:0]) +
	( 16'sd 29390) * $signed(input_fmap_151[7:0]) +
	( 15'sd 15252) * $signed(input_fmap_152[7:0]) +
	( 14'sd 7959) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24472) * $signed(input_fmap_154[7:0]) +
	( 15'sd 11962) * $signed(input_fmap_155[7:0]) +
	( 13'sd 2873) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6483) * $signed(input_fmap_157[7:0]) +
	( 16'sd 19899) * $signed(input_fmap_158[7:0]) +
	( 16'sd 17801) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11399) * $signed(input_fmap_160[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10846) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15213) * $signed(input_fmap_163[7:0]) +
	( 16'sd 29057) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19231) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22103) * $signed(input_fmap_166[7:0]) +
	( 16'sd 25046) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1194) * $signed(input_fmap_168[7:0]) +
	( 16'sd 32582) * $signed(input_fmap_169[7:0]) +
	( 11'sd 615) * $signed(input_fmap_170[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6956) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27915) * $signed(input_fmap_173[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3675) * $signed(input_fmap_175[7:0]) +
	( 16'sd 25102) * $signed(input_fmap_176[7:0]) +
	( 15'sd 9151) * $signed(input_fmap_177[7:0]) +
	( 14'sd 4435) * $signed(input_fmap_178[7:0]) +
	( 15'sd 11613) * $signed(input_fmap_179[7:0]) +
	( 16'sd 31136) * $signed(input_fmap_180[7:0]) +
	( 14'sd 4278) * $signed(input_fmap_181[7:0]) +
	( 16'sd 17173) * $signed(input_fmap_182[7:0]) +
	( 16'sd 26528) * $signed(input_fmap_183[7:0]) +
	( 16'sd 19818) * $signed(input_fmap_184[7:0]) +
	( 15'sd 10237) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18297) * $signed(input_fmap_186[7:0]) +
	( 16'sd 24951) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13327) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30431) * $signed(input_fmap_189[7:0]) +
	( 15'sd 12836) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19682) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20052) * $signed(input_fmap_192[7:0]) +
	( 13'sd 2079) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9069) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29345) * $signed(input_fmap_195[7:0]) +
	( 9'sd 150) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22588) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9926) * $signed(input_fmap_198[7:0]) +
	( 15'sd 15130) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_200[7:0]) +
	( 15'sd 16115) * $signed(input_fmap_201[7:0]) +
	( 16'sd 29675) * $signed(input_fmap_202[7:0]) +
	( 16'sd 27914) * $signed(input_fmap_203[7:0]) +
	( 16'sd 25364) * $signed(input_fmap_204[7:0]) +
	( 16'sd 32644) * $signed(input_fmap_205[7:0]) +
	( 16'sd 22122) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30847) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4560) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3369) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9749) * $signed(input_fmap_210[7:0]) +
	( 15'sd 8592) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14538) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2701) * $signed(input_fmap_213[7:0]) +
	( 14'sd 4268) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22293) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17742) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_217[7:0]) +
	( 15'sd 15383) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21839) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25987) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27964) * $signed(input_fmap_221[7:0]) +
	( 16'sd 17967) * $signed(input_fmap_222[7:0]) +
	( 14'sd 5245) * $signed(input_fmap_223[7:0]) +
	( 15'sd 15593) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26273) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31998) * $signed(input_fmap_226[7:0]) +
	( 16'sd 29260) * $signed(input_fmap_227[7:0]) +
	( 16'sd 23815) * $signed(input_fmap_228[7:0]) +
	( 16'sd 21010) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_230[7:0]) +
	( 16'sd 23762) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9170) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27652) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15641) * $signed(input_fmap_234[7:0]) +
	( 14'sd 6106) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27898) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19129) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28792) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20982) * $signed(input_fmap_239[7:0]) +
	( 15'sd 11811) * $signed(input_fmap_240[7:0]) +
	( 16'sd 31347) * $signed(input_fmap_241[7:0]) +
	( 15'sd 13969) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22154) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18380) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24041) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1703) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21887) * $signed(input_fmap_247[7:0]) +
	( 15'sd 8240) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2763) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17968) * $signed(input_fmap_250[7:0]) +
	( 16'sd 28283) * $signed(input_fmap_251[7:0]) +
	( 14'sd 8034) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29892) * $signed(input_fmap_253[7:0]) +
	( 16'sd 25195) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14678) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_45;
assign conv_mac_45 = 
	( 13'sd 3619) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5271) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27215) * $signed(input_fmap_2[7:0]) +
	( 11'sd 799) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22521) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27189) * $signed(input_fmap_5[7:0]) +
	( 11'sd 827) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13192) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11744) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22012) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7559) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29653) * $signed(input_fmap_11[7:0]) +
	( 9'sd 137) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14273) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30715) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7385) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21764) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27262) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31338) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25200) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1296) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21873) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13240) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2755) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21963) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7661) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6081) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25830) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9537) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26593) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8866) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5610) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3151) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23413) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18339) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2478) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4294) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18920) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11889) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19026) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29366) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21623) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28992) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7621) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6272) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25441) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25078) * $signed(input_fmap_50[7:0]) +
	( 10'sd 475) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19599) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22952) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1931) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17144) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9127) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4800) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13215) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6020) * $signed(input_fmap_60[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28070) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29864) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28014) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16318) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2581) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28307) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18642) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12929) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16617) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3559) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1693) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8475) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20413) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3133) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11344) * $signed(input_fmap_80[7:0]) +
	( 10'sd 494) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12294) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10916) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28853) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16983) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22238) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25297) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28544) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2095) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11056) * $signed(input_fmap_91[7:0]) +
	( 11'sd 804) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27368) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9655) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25036) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31715) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4322) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27703) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5384) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31895) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9126) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21271) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5505) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10249) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8257) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4224) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13256) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17471) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4934) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2505) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10397) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13064) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18268) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9030) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20254) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16612) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10180) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19031) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12240) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14766) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4179) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3987) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15610) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13802) * $signed(input_fmap_129[7:0]) +
	( 16'sd 28863) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31806) * $signed(input_fmap_131[7:0]) +
	( 16'sd 20196) * $signed(input_fmap_132[7:0]) +
	( 16'sd 23245) * $signed(input_fmap_133[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21447) * $signed(input_fmap_135[7:0]) +
	( 14'sd 5402) * $signed(input_fmap_136[7:0]) +
	( 11'sd 749) * $signed(input_fmap_137[7:0]) +
	( 16'sd 25366) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8945) * $signed(input_fmap_139[7:0]) +
	( 14'sd 4306) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_142[7:0]) +
	( 16'sd 30662) * $signed(input_fmap_143[7:0]) +
	( 16'sd 26243) * $signed(input_fmap_144[7:0]) +
	( 14'sd 4455) * $signed(input_fmap_145[7:0]) +
	( 16'sd 31229) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27793) * $signed(input_fmap_147[7:0]) +
	( 16'sd 29293) * $signed(input_fmap_148[7:0]) +
	( 14'sd 8118) * $signed(input_fmap_149[7:0]) +
	( 15'sd 14967) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24919) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20372) * $signed(input_fmap_152[7:0]) +
	( 16'sd 19281) * $signed(input_fmap_153[7:0]) +
	( 16'sd 32739) * $signed(input_fmap_154[7:0]) +
	( 16'sd 26176) * $signed(input_fmap_155[7:0]) +
	( 14'sd 6105) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17017) * $signed(input_fmap_158[7:0]) +
	( 15'sd 15400) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22253) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30030) * $signed(input_fmap_162[7:0]) +
	( 16'sd 23709) * $signed(input_fmap_163[7:0]) +
	( 16'sd 30340) * $signed(input_fmap_164[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2741) * $signed(input_fmap_166[7:0]) +
	( 16'sd 29504) * $signed(input_fmap_167[7:0]) +
	( 16'sd 18577) * $signed(input_fmap_168[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7716) * $signed(input_fmap_170[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14368) * $signed(input_fmap_172[7:0]) +
	( 14'sd 7313) * $signed(input_fmap_173[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_174[7:0]) +
	( 16'sd 23436) * $signed(input_fmap_175[7:0]) +
	( 9'sd 217) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29408) * $signed(input_fmap_177[7:0]) +
	( 16'sd 28822) * $signed(input_fmap_178[7:0]) +
	( 11'sd 608) * $signed(input_fmap_179[7:0]) +
	( 15'sd 12795) * $signed(input_fmap_180[7:0]) +
	( 15'sd 12878) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29190) * $signed(input_fmap_183[7:0]) +
	( 15'sd 15837) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_185[7:0]) +
	( 15'sd 11239) * $signed(input_fmap_186[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_187[7:0]) +
	( 15'sd 10065) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2082) * $signed(input_fmap_189[7:0]) +
	( 12'sd 1934) * $signed(input_fmap_190[7:0]) +
	( 16'sd 27013) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15750) * $signed(input_fmap_192[7:0]) +
	( 12'sd 2029) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21020) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22247) * $signed(input_fmap_195[7:0]) +
	( 13'sd 3327) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1048) * $signed(input_fmap_197[7:0]) +
	( 15'sd 15142) * $signed(input_fmap_198[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_199[7:0]) +
	( 11'sd 591) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6572) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31546) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24936) * $signed(input_fmap_203[7:0]) +
	( 16'sd 26425) * $signed(input_fmap_204[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12068) * $signed(input_fmap_206[7:0]) +
	( 16'sd 25929) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15504) * $signed(input_fmap_208[7:0]) +
	( 16'sd 29297) * $signed(input_fmap_209[7:0]) +
	( 15'sd 14732) * $signed(input_fmap_210[7:0]) +
	( 14'sd 7918) * $signed(input_fmap_211[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_212[7:0]) +
	( 16'sd 26268) * $signed(input_fmap_213[7:0]) +
	( 16'sd 26472) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9426) * $signed(input_fmap_215[7:0]) +
	( 16'sd 29388) * $signed(input_fmap_216[7:0]) +
	( 15'sd 16241) * $signed(input_fmap_217[7:0]) +
	( 15'sd 9774) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10679) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13684) * $signed(input_fmap_220[7:0]) +
	( 14'sd 7019) * $signed(input_fmap_221[7:0]) +
	( 16'sd 22267) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2616) * $signed(input_fmap_223[7:0]) +
	( 16'sd 28807) * $signed(input_fmap_224[7:0]) +
	( 16'sd 30943) * $signed(input_fmap_225[7:0]) +
	( 15'sd 12974) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9064) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29010) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29955) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3392) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7307) * $signed(input_fmap_232[7:0]) +
	( 16'sd 26902) * $signed(input_fmap_233[7:0]) +
	( 16'sd 17202) * $signed(input_fmap_234[7:0]) +
	( 15'sd 10052) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10014) * $signed(input_fmap_236[7:0]) +
	( 16'sd 24201) * $signed(input_fmap_237[7:0]) +
	( 16'sd 29169) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20215) * $signed(input_fmap_239[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_240[7:0]) +
	( 11'sd 754) * $signed(input_fmap_241[7:0]) +
	( 15'sd 13441) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7214) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22699) * $signed(input_fmap_244[7:0]) +
	( 14'sd 4707) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14979) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17228) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32439) * $signed(input_fmap_248[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9832) * $signed(input_fmap_250[7:0]) +
	( 16'sd 31882) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12202) * $signed(input_fmap_252[7:0]) +
	( 15'sd 9467) * $signed(input_fmap_253[7:0]) +
	( 16'sd 17654) * $signed(input_fmap_254[7:0]) +
	( 10'sd 483) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_46;
assign conv_mac_46 = 
	( 14'sd 6552) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4570) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3663) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11413) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4591) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11748) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5673) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8533) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21172) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10559) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19395) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31539) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23548) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12376) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2992) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7244) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24439) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2927) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24876) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23757) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27329) * $signed(input_fmap_24[7:0]) +
	( 7'sd 49) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8227) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30489) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31322) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18024) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16614) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5708) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30074) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14291) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3085) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24912) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26992) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11286) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22762) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25228) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17780) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29033) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11164) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27428) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_46[7:0]) +
	( 10'sd 369) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5992) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1905) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8445) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5220) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22804) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1741) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5176) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23496) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23367) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20676) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10530) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10454) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5175) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29643) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16118) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10689) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8415) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2249) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4858) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3586) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28573) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1164) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31686) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4919) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2954) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31376) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6404) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15664) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5131) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24383) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7352) * $signed(input_fmap_79[7:0]) +
	( 9'sd 196) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8247) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8871) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9165) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20029) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30047) * $signed(input_fmap_86[7:0]) +
	( 11'sd 864) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25907) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23433) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25882) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20915) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2516) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7044) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26102) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17481) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15160) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28249) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13357) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21558) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23656) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1855) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20937) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23703) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30563) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13496) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31080) * $signed(input_fmap_106[7:0]) +
	( 11'sd 544) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5106) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2228) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7717) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25049) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23440) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29176) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3159) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11892) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2706) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7468) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32172) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29565) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19416) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4329) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28813) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6422) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24289) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23386) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2748) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7259) * $signed(input_fmap_127[7:0]) +
	( 16'sd 26169) * $signed(input_fmap_128[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_129[7:0]) +
	( 15'sd 13114) * $signed(input_fmap_130[7:0]) +
	( 11'sd 1018) * $signed(input_fmap_131[7:0]) +
	( 16'sd 31063) * $signed(input_fmap_132[7:0]) +
	( 15'sd 15376) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19842) * $signed(input_fmap_134[7:0]) +
	( 14'sd 7221) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17059) * $signed(input_fmap_136[7:0]) +
	( 16'sd 29674) * $signed(input_fmap_137[7:0]) +
	( 16'sd 30565) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30604) * $signed(input_fmap_140[7:0]) +
	( 16'sd 23259) * $signed(input_fmap_141[7:0]) +
	( 13'sd 3136) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26496) * $signed(input_fmap_143[7:0]) +
	( 11'sd 899) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26995) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18020) * $signed(input_fmap_146[7:0]) +
	( 16'sd 22188) * $signed(input_fmap_147[7:0]) +
	( 12'sd 2032) * $signed(input_fmap_148[7:0]) +
	( 15'sd 11383) * $signed(input_fmap_149[7:0]) +
	( 14'sd 7503) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19303) * $signed(input_fmap_151[7:0]) +
	( 13'sd 3393) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1949) * $signed(input_fmap_153[7:0]) +
	( 13'sd 2659) * $signed(input_fmap_154[7:0]) +
	( 16'sd 25697) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29757) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13796) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4967) * $signed(input_fmap_158[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_159[7:0]) +
	( 13'sd 2440) * $signed(input_fmap_160[7:0]) +
	( 14'sd 6907) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29332) * $signed(input_fmap_162[7:0]) +
	( 15'sd 13579) * $signed(input_fmap_163[7:0]) +
	( 14'sd 7470) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_165[7:0]) +
	( 16'sd 21074) * $signed(input_fmap_166[7:0]) +
	( 13'sd 2225) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_169[7:0]) +
	( 16'sd 19748) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4730) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29707) * $signed(input_fmap_173[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_174[7:0]) +
	( 10'sd 430) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7503) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15706) * $signed(input_fmap_177[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18881) * $signed(input_fmap_179[7:0]) +
	( 16'sd 20547) * $signed(input_fmap_180[7:0]) +
	( 15'sd 8389) * $signed(input_fmap_181[7:0]) +
	( 14'sd 7517) * $signed(input_fmap_182[7:0]) +
	( 15'sd 14343) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24715) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17256) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4367) * $signed(input_fmap_187[7:0]) +
	( 16'sd 26434) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25990) * $signed(input_fmap_189[7:0]) +
	( 16'sd 25046) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23157) * $signed(input_fmap_191[7:0]) +
	( 14'sd 4883) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30196) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27305) * $signed(input_fmap_194[7:0]) +
	( 15'sd 15212) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17875) * $signed(input_fmap_196[7:0]) +
	( 9'sd 219) * $signed(input_fmap_197[7:0]) +
	( 9'sd 183) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1048) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5454) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9373) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31272) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21263) * $signed(input_fmap_203[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_204[7:0]) +
	( 14'sd 4777) * $signed(input_fmap_205[7:0]) +
	( 16'sd 26916) * $signed(input_fmap_206[7:0]) +
	( 15'sd 9197) * $signed(input_fmap_207[7:0]) +
	( 6'sd 31) * $signed(input_fmap_208[7:0]) +
	( 14'sd 5778) * $signed(input_fmap_209[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_210[7:0]) +
	( 16'sd 27693) * $signed(input_fmap_211[7:0]) +
	( 16'sd 32458) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28831) * $signed(input_fmap_213[7:0]) +
	( 13'sd 3528) * $signed(input_fmap_214[7:0]) +
	( 16'sd 18439) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1922) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19450) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13293) * $signed(input_fmap_218[7:0]) +
	( 14'sd 7553) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19605) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19538) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10711) * $signed(input_fmap_222[7:0]) +
	( 16'sd 31966) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_224[7:0]) +
	( 16'sd 21420) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32489) * $signed(input_fmap_226[7:0]) +
	( 16'sd 26866) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22170) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_229[7:0]) +
	( 14'sd 5981) * $signed(input_fmap_230[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_231[7:0]) +
	( 16'sd 24894) * $signed(input_fmap_232[7:0]) +
	( 16'sd 20756) * $signed(input_fmap_233[7:0]) +
	( 15'sd 9175) * $signed(input_fmap_234[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10892) * $signed(input_fmap_236[7:0]) +
	( 15'sd 8318) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16836) * $signed(input_fmap_238[7:0]) +
	( 15'sd 15607) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19361) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20730) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23053) * $signed(input_fmap_242[7:0]) +
	( 16'sd 26500) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24096) * $signed(input_fmap_244[7:0]) +
	( 15'sd 11967) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1474) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15277) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3989) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21780) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24376) * $signed(input_fmap_250[7:0]) +
	( 16'sd 32211) * $signed(input_fmap_251[7:0]) +
	( 13'sd 3724) * $signed(input_fmap_252[7:0]) +
	( 14'sd 8102) * $signed(input_fmap_253[7:0]) +
	( 16'sd 28082) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10858) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_47;
assign conv_mac_47 = 
	( 10'sd 311) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_1[7:0]) +
	( 13'sd 4085) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31232) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14695) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27084) * $signed(input_fmap_5[7:0]) +
	( 11'sd 529) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12205) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19478) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24784) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16789) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13023) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3907) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28721) * $signed(input_fmap_13[7:0]) +
	( 12'sd 2039) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3587) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5918) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4645) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21410) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6833) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18231) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3666) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30228) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23861) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17274) * $signed(input_fmap_25[7:0]) +
	( 11'sd 1001) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14011) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5339) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8506) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10376) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1105) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27701) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21807) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30232) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19646) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32632) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10434) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29531) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13942) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7303) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10292) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9085) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16157) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17649) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11162) * $signed(input_fmap_47[7:0]) +
	( 11'sd 643) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32678) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27363) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30532) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13853) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5851) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2146) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22090) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5487) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10054) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16585) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10937) * $signed(input_fmap_61[7:0]) +
	( 11'sd 901) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22942) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16612) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20370) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8571) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15685) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4876) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31527) * $signed(input_fmap_69[7:0]) +
	( 13'sd 4021) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12316) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13835) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6777) * $signed(input_fmap_73[7:0]) +
	( 9'sd 203) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14721) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15743) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5616) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3513) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18558) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8534) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17863) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11733) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9109) * $signed(input_fmap_88[7:0]) +
	( 13'sd 4021) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29393) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12291) * $signed(input_fmap_91[7:0]) +
	( 9'sd 196) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20768) * $signed(input_fmap_93[7:0]) +
	( 9'sd 132) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4196) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3746) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29388) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6863) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8800) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15997) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16556) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16516) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18926) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31747) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9940) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6571) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_108[7:0]) +
	( 14'sd 8137) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12630) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19547) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3939) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17135) * $signed(input_fmap_113[7:0]) +
	( 11'sd 863) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15881) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11605) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24522) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7931) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15571) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28039) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16789) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5837) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25969) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5444) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23310) * $signed(input_fmap_128[7:0]) +
	( 16'sd 22689) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_130[7:0]) +
	( 16'sd 27258) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25109) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22784) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11901) * $signed(input_fmap_134[7:0]) +
	( 15'sd 9114) * $signed(input_fmap_135[7:0]) +
	( 15'sd 11842) * $signed(input_fmap_136[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_138[7:0]) +
	( 12'sd 1314) * $signed(input_fmap_139[7:0]) +
	( 15'sd 8727) * $signed(input_fmap_140[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_141[7:0]) +
	( 15'sd 9492) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7504) * $signed(input_fmap_143[7:0]) +
	( 16'sd 21126) * $signed(input_fmap_144[7:0]) +
	( 14'sd 4971) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19630) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17422) * $signed(input_fmap_147[7:0]) +
	( 15'sd 13525) * $signed(input_fmap_148[7:0]) +
	( 16'sd 20608) * $signed(input_fmap_149[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17036) * $signed(input_fmap_151[7:0]) +
	( 16'sd 25272) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23726) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4595) * $signed(input_fmap_154[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28723) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25141) * $signed(input_fmap_157[7:0]) +
	( 15'sd 15277) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5843) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_160[7:0]) +
	( 16'sd 17402) * $signed(input_fmap_161[7:0]) +
	( 16'sd 16646) * $signed(input_fmap_162[7:0]) +
	( 14'sd 6666) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_164[7:0]) +
	( 16'sd 29110) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30237) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20402) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14750) * $signed(input_fmap_168[7:0]) +
	( 16'sd 31937) * $signed(input_fmap_169[7:0]) +
	( 15'sd 15990) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11469) * $signed(input_fmap_171[7:0]) +
	( 9'sd 149) * $signed(input_fmap_172[7:0]) +
	( 13'sd 3571) * $signed(input_fmap_173[7:0]) +
	( 16'sd 23726) * $signed(input_fmap_174[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13555) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29386) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32621) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28694) * $signed(input_fmap_179[7:0]) +
	( 15'sd 10348) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18692) * $signed(input_fmap_181[7:0]) +
	( 13'sd 3807) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27246) * $signed(input_fmap_183[7:0]) +
	( 16'sd 27615) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26513) * $signed(input_fmap_185[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_186[7:0]) +
	( 9'sd 157) * $signed(input_fmap_187[7:0]) +
	( 16'sd 16732) * $signed(input_fmap_188[7:0]) +
	( 15'sd 10967) * $signed(input_fmap_189[7:0]) +
	( 15'sd 10387) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20647) * $signed(input_fmap_191[7:0]) +
	( 16'sd 32697) * $signed(input_fmap_192[7:0]) +
	( 13'sd 2075) * $signed(input_fmap_193[7:0]) +
	( 16'sd 20539) * $signed(input_fmap_194[7:0]) +
	( 16'sd 28239) * $signed(input_fmap_195[7:0]) +
	( 16'sd 31602) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26044) * $signed(input_fmap_197[7:0]) +
	( 15'sd 12955) * $signed(input_fmap_198[7:0]) +
	( 16'sd 22503) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3311) * $signed(input_fmap_200[7:0]) +
	( 16'sd 20316) * $signed(input_fmap_201[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_202[7:0]) +
	( 16'sd 29327) * $signed(input_fmap_203[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_204[7:0]) +
	( 13'sd 4022) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2432) * $signed(input_fmap_206[7:0]) +
	( 16'sd 24999) * $signed(input_fmap_207[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20190) * $signed(input_fmap_209[7:0]) +
	( 11'sd 633) * $signed(input_fmap_210[7:0]) +
	( 15'sd 16258) * $signed(input_fmap_211[7:0]) +
	( 16'sd 21961) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12712) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31287) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2781) * $signed(input_fmap_215[7:0]) +
	( 16'sd 16863) * $signed(input_fmap_216[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28028) * $signed(input_fmap_218[7:0]) +
	( 13'sd 2729) * $signed(input_fmap_219[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15107) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_222[7:0]) +
	( 16'sd 30175) * $signed(input_fmap_223[7:0]) +
	( 15'sd 16118) * $signed(input_fmap_224[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29541) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22920) * $signed(input_fmap_227[7:0]) +
	( 15'sd 12592) * $signed(input_fmap_228[7:0]) +
	( 16'sd 31570) * $signed(input_fmap_229[7:0]) +
	( 16'sd 25517) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7614) * $signed(input_fmap_231[7:0]) +
	( 14'sd 4356) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5095) * $signed(input_fmap_233[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7804) * $signed(input_fmap_235[7:0]) +
	( 16'sd 26525) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2507) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13534) * $signed(input_fmap_238[7:0]) +
	( 14'sd 7585) * $signed(input_fmap_239[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30378) * $signed(input_fmap_241[7:0]) +
	( 16'sd 21286) * $signed(input_fmap_242[7:0]) +
	( 13'sd 3187) * $signed(input_fmap_243[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_244[7:0]) +
	( 15'sd 9399) * $signed(input_fmap_245[7:0]) +
	( 14'sd 7944) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15992) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18944) * $signed(input_fmap_248[7:0]) +
	( 15'sd 11946) * $signed(input_fmap_249[7:0]) +
	( 14'sd 5255) * $signed(input_fmap_250[7:0]) +
	( 16'sd 29951) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_252[7:0]) +
	( 16'sd 20510) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19373) * $signed(input_fmap_254[7:0]) +
	( 13'sd 3016) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_48;
assign conv_mac_48 = 
	( 15'sd 14784) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30259) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5621) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4791) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17917) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1820) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2911) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31130) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8536) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5365) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23284) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24441) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11250) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32676) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12755) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18295) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28947) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18367) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9195) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7050) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17682) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11349) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1727) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7138) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21113) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29355) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17730) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26919) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31016) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5901) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26030) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30923) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22774) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9383) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17827) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27195) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24204) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7436) * $signed(input_fmap_40[7:0]) +
	( 10'sd 291) * $signed(input_fmap_41[7:0]) +
	( 11'sd 636) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2779) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3010) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9185) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18428) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28997) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20410) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5339) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8637) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9688) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22777) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20905) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22700) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17730) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22264) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5203) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32547) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5204) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16194) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9437) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16192) * $signed(input_fmap_63[7:0]) +
	( 7'sd 36) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19495) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14248) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26263) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24622) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11244) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27878) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32607) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23299) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26559) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14785) * $signed(input_fmap_75[7:0]) +
	( 9'sd 233) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_77[7:0]) +
	( 11'sd 815) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23947) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25545) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_81[7:0]) +
	( 13'sd 4046) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4741) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6018) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7191) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21169) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29489) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15435) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1186) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16808) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2110) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2243) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2202) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17246) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26552) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10620) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10259) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15216) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23678) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22461) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32232) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25194) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26141) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31127) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27928) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10562) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14123) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12213) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12612) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1695) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26695) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4735) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24295) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19041) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15477) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11659) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11327) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29397) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8169) * $signed(input_fmap_127[7:0]) +
	( 16'sd 22692) * $signed(input_fmap_128[7:0]) +
	( 15'sd 11910) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6075) * $signed(input_fmap_130[7:0]) +
	( 10'sd 505) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_132[7:0]) +
	( 15'sd 14894) * $signed(input_fmap_133[7:0]) +
	( 16'sd 27619) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26167) * $signed(input_fmap_135[7:0]) +
	( 15'sd 11158) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15449) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9398) * $signed(input_fmap_138[7:0]) +
	( 16'sd 19576) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_140[7:0]) +
	( 15'sd 16060) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30699) * $signed(input_fmap_142[7:0]) +
	( 16'sd 18624) * $signed(input_fmap_143[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_144[7:0]) +
	( 12'sd 1880) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7347) * $signed(input_fmap_146[7:0]) +
	( 15'sd 10569) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22863) * $signed(input_fmap_148[7:0]) +
	( 16'sd 31268) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15615) * $signed(input_fmap_150[7:0]) +
	( 16'sd 16458) * $signed(input_fmap_151[7:0]) +
	( 15'sd 15752) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24140) * $signed(input_fmap_153[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_154[7:0]) +
	( 15'sd 15962) * $signed(input_fmap_155[7:0]) +
	( 16'sd 27545) * $signed(input_fmap_156[7:0]) +
	( 16'sd 26241) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17250) * $signed(input_fmap_158[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_159[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_160[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_161[7:0]) +
	( 16'sd 17938) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3525) * $signed(input_fmap_163[7:0]) +
	( 16'sd 21848) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4280) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3131) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23746) * $signed(input_fmap_167[7:0]) +
	( 13'sd 2484) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12818) * $signed(input_fmap_169[7:0]) +
	( 15'sd 8607) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_171[7:0]) +
	( 16'sd 23886) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6941) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21835) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_176[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_177[7:0]) +
	( 14'sd 5524) * $signed(input_fmap_178[7:0]) +
	( 15'sd 12640) * $signed(input_fmap_179[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18227) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6708) * $signed(input_fmap_182[7:0]) +
	( 16'sd 19319) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31408) * $signed(input_fmap_184[7:0]) +
	( 15'sd 14192) * $signed(input_fmap_185[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_186[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_187[7:0]) +
	( 16'sd 20602) * $signed(input_fmap_188[7:0]) +
	( 15'sd 9553) * $signed(input_fmap_189[7:0]) +
	( 14'sd 7366) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20273) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31935) * $signed(input_fmap_192[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_193[7:0]) +
	( 16'sd 20095) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1934) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19128) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1565) * $signed(input_fmap_197[7:0]) +
	( 15'sd 16035) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20228) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8939) * $signed(input_fmap_200[7:0]) +
	( 16'sd 23785) * $signed(input_fmap_201[7:0]) +
	( 12'sd 1842) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19472) * $signed(input_fmap_203[7:0]) +
	( 16'sd 16788) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6530) * $signed(input_fmap_205[7:0]) +
	( 15'sd 16115) * $signed(input_fmap_206[7:0]) +
	( 15'sd 15323) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8229) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19349) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11634) * $signed(input_fmap_210[7:0]) +
	( 12'sd 1559) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_212[7:0]) +
	( 14'sd 7048) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20791) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6831) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30081) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8713) * $signed(input_fmap_218[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_219[7:0]) +
	( 15'sd 8754) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23104) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28398) * $signed(input_fmap_222[7:0]) +
	( 13'sd 3389) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25953) * $signed(input_fmap_224[7:0]) +
	( 15'sd 16226) * $signed(input_fmap_225[7:0]) +
	( 14'sd 8175) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13365) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8539) * $signed(input_fmap_228[7:0]) +
	( 16'sd 21435) * $signed(input_fmap_229[7:0]) +
	( 13'sd 3427) * $signed(input_fmap_230[7:0]) +
	( 16'sd 22746) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15297) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27661) * $signed(input_fmap_233[7:0]) +
	( 16'sd 27059) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7051) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28701) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20037) * $signed(input_fmap_237[7:0]) +
	( 16'sd 24998) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31956) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19121) * $signed(input_fmap_240[7:0]) +
	( 13'sd 2541) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27995) * $signed(input_fmap_242[7:0]) +
	( 16'sd 16954) * $signed(input_fmap_243[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7522) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9104) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3230) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21071) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24540) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28860) * $signed(input_fmap_253[7:0]) +
	( 16'sd 27778) * $signed(input_fmap_254[7:0]) +
	( 14'sd 4501) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_49;
assign conv_mac_49 = 
	( 16'sd 19848) * $signed(input_fmap_0[7:0]) +
	( 15'sd 12712) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5830) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24294) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28149) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31167) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20112) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2175) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17417) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15786) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32745) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21998) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1746) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18048) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6307) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29599) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13246) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16949) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31002) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20675) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22177) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7407) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28919) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32703) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1179) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13375) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20633) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27734) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6397) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19313) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25997) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25639) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22295) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11780) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9939) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30459) * $signed(input_fmap_40[7:0]) +
	( 12'sd 2006) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12642) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26077) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9187) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28060) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8430) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29928) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29053) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22032) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20408) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14257) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31033) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17834) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25041) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16161) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7590) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20529) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19688) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9375) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28519) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23906) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12085) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11062) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27328) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15527) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7591) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28618) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18722) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6592) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19515) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24041) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5470) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5326) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21871) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21979) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7349) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26104) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21585) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1438) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19217) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23815) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8479) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13118) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22995) * $signed(input_fmap_88[7:0]) +
	( 11'sd 527) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23373) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17136) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14475) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24273) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10315) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12131) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8491) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12350) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15916) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1535) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24107) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12057) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14494) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2730) * $signed(input_fmap_104[7:0]) +
	( 10'sd 325) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29889) * $signed(input_fmap_108[7:0]) +
	( 16'sd 27661) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22426) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31639) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30990) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18654) * $signed(input_fmap_113[7:0]) +
	( 10'sd 506) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23956) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1501) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4251) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26650) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25026) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6078) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16758) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13555) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23004) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25599) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13444) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22964) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8170) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4521) * $signed(input_fmap_128[7:0]) +
	( 15'sd 8295) * $signed(input_fmap_129[7:0]) +
	( 16'sd 23914) * $signed(input_fmap_130[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_131[7:0]) +
	( 13'sd 2209) * $signed(input_fmap_132[7:0]) +
	( 16'sd 27627) * $signed(input_fmap_133[7:0]) +
	( 15'sd 15332) * $signed(input_fmap_134[7:0]) +
	( 11'sd 883) * $signed(input_fmap_135[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26810) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29148) * $signed(input_fmap_138[7:0]) +
	( 16'sd 30613) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28396) * $signed(input_fmap_140[7:0]) +
	( 10'sd 402) * $signed(input_fmap_141[7:0]) +
	( 16'sd 16572) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31270) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3689) * $signed(input_fmap_144[7:0]) +
	( 12'sd 2041) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27501) * $signed(input_fmap_146[7:0]) +
	( 16'sd 25147) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28431) * $signed(input_fmap_148[7:0]) +
	( 16'sd 32373) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15138) * $signed(input_fmap_150[7:0]) +
	( 16'sd 21803) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29838) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24473) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6560) * $signed(input_fmap_154[7:0]) +
	( 16'sd 31714) * $signed(input_fmap_155[7:0]) +
	( 15'sd 11042) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22369) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14487) * $signed(input_fmap_159[7:0]) +
	( 16'sd 19200) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4693) * $signed(input_fmap_161[7:0]) +
	( 16'sd 23995) * $signed(input_fmap_162[7:0]) +
	( 16'sd 17054) * $signed(input_fmap_163[7:0]) +
	( 16'sd 29869) * $signed(input_fmap_164[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_165[7:0]) +
	( 16'sd 24755) * $signed(input_fmap_166[7:0]) +
	( 15'sd 12231) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5481) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6518) * $signed(input_fmap_169[7:0]) +
	( 10'sd 351) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20245) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7074) * $signed(input_fmap_172[7:0]) +
	( 13'sd 3789) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_174[7:0]) +
	( 15'sd 11593) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29673) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31080) * $signed(input_fmap_177[7:0]) +
	( 14'sd 4347) * $signed(input_fmap_178[7:0]) +
	( 10'sd 477) * $signed(input_fmap_179[7:0]) +
	( 10'sd 450) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3213) * $signed(input_fmap_181[7:0]) +
	( 14'sd 7961) * $signed(input_fmap_182[7:0]) +
	( 13'sd 3122) * $signed(input_fmap_183[7:0]) +
	( 14'sd 6650) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_185[7:0]) +
	( 16'sd 20830) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1037) * $signed(input_fmap_187[7:0]) +
	( 16'sd 26904) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2073) * $signed(input_fmap_189[7:0]) +
	( 12'sd 1512) * $signed(input_fmap_190[7:0]) +
	( 15'sd 15274) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27870) * $signed(input_fmap_192[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_193[7:0]) +
	( 16'sd 32325) * $signed(input_fmap_194[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_195[7:0]) +
	( 16'sd 28626) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22111) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5572) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13336) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12895) * $signed(input_fmap_201[7:0]) +
	( 11'sd 769) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30173) * $signed(input_fmap_203[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5986) * $signed(input_fmap_205[7:0]) +
	( 14'sd 7374) * $signed(input_fmap_206[7:0]) +
	( 14'sd 6099) * $signed(input_fmap_207[7:0]) +
	( 15'sd 10953) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19346) * $signed(input_fmap_209[7:0]) +
	( 16'sd 21352) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26914) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23466) * $signed(input_fmap_213[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_214[7:0]) +
	( 16'sd 31257) * $signed(input_fmap_215[7:0]) +
	( 16'sd 22575) * $signed(input_fmap_216[7:0]) +
	( 15'sd 12145) * $signed(input_fmap_217[7:0]) +
	( 13'sd 4001) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10030) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24368) * $signed(input_fmap_220[7:0]) +
	( 16'sd 21728) * $signed(input_fmap_221[7:0]) +
	( 16'sd 27468) * $signed(input_fmap_222[7:0]) +
	( 11'sd 515) * $signed(input_fmap_223[7:0]) +
	( 16'sd 21438) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26815) * $signed(input_fmap_225[7:0]) +
	( 16'sd 25174) * $signed(input_fmap_226[7:0]) +
	( 14'sd 7794) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19096) * $signed(input_fmap_228[7:0]) +
	( 16'sd 16574) * $signed(input_fmap_229[7:0]) +
	( 12'sd 1208) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3628) * $signed(input_fmap_231[7:0]) +
	( 13'sd 2836) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_233[7:0]) +
	( 15'sd 8356) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19517) * $signed(input_fmap_235[7:0]) +
	( 16'sd 24252) * $signed(input_fmap_236[7:0]) +
	( 14'sd 7186) * $signed(input_fmap_237[7:0]) +
	( 16'sd 21127) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5718) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6461) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29731) * $signed(input_fmap_241[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_242[7:0]) +
	( 16'sd 16799) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18814) * $signed(input_fmap_244[7:0]) +
	( 16'sd 18757) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20964) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13372) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_248[7:0]) +
	( 16'sd 18230) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_250[7:0]) +
	( 16'sd 30908) * $signed(input_fmap_251[7:0]) +
	( 16'sd 16828) * $signed(input_fmap_252[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20407) * $signed(input_fmap_254[7:0]) +
	( 14'sd 4245) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_50;
assign conv_mac_50 = 
	( 16'sd 27417) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16095) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19140) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3076) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5520) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10232) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8874) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4882) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27318) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20838) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12091) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31789) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32402) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23589) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27808) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5912) * $signed(input_fmap_16[7:0]) +
	( 11'sd 893) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23702) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18865) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30951) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21367) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17948) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21835) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1367) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26745) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23495) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27886) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28964) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31671) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4329) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29244) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12955) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10845) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30398) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19667) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6377) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31379) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15807) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11311) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21656) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16038) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14759) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23163) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31713) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20641) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14247) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14595) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8659) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4939) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2759) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11100) * $signed(input_fmap_59[7:0]) +
	( 10'sd 262) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11492) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2371) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5853) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1568) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20531) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21195) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10096) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1872) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20666) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10326) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30139) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8275) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5558) * $signed(input_fmap_75[7:0]) +
	( 11'sd 520) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2983) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10131) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1146) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11469) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22638) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1635) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13903) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20822) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21011) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17685) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31673) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27461) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12020) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30488) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12705) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31705) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6473) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16782) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9006) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31415) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12321) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21863) * $signed(input_fmap_103[7:0]) +
	( 10'sd 504) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15718) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14437) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17072) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19433) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6947) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25867) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30837) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24449) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11225) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26999) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3847) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22892) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5796) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11976) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30672) * $signed(input_fmap_120[7:0]) +
	( 9'sd 171) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9642) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24652) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11635) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8814) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15602) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29967) * $signed(input_fmap_128[7:0]) +
	( 15'sd 8753) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14481) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19755) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11882) * $signed(input_fmap_132[7:0]) +
	( 16'sd 24212) * $signed(input_fmap_133[7:0]) +
	( 15'sd 13982) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26007) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25503) * $signed(input_fmap_136[7:0]) +
	( 14'sd 7488) * $signed(input_fmap_137[7:0]) +
	( 16'sd 26615) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27472) * $signed(input_fmap_139[7:0]) +
	( 16'sd 25973) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31831) * $signed(input_fmap_141[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_142[7:0]) +
	( 16'sd 27275) * $signed(input_fmap_143[7:0]) +
	( 16'sd 29329) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25588) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15432) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29253) * $signed(input_fmap_147[7:0]) +
	( 15'sd 14785) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17404) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21456) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19699) * $signed(input_fmap_151[7:0]) +
	( 16'sd 32429) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3686) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31463) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29596) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11859) * $signed(input_fmap_157[7:0]) +
	( 10'sd 437) * $signed(input_fmap_158[7:0]) +
	( 16'sd 28821) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5570) * $signed(input_fmap_160[7:0]) +
	( 15'sd 13348) * $signed(input_fmap_161[7:0]) +
	( 16'sd 16689) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32057) * $signed(input_fmap_163[7:0]) +
	( 14'sd 4201) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_165[7:0]) +
	( 16'sd 20065) * $signed(input_fmap_166[7:0]) +
	( 16'sd 28350) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4551) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18537) * $signed(input_fmap_169[7:0]) +
	( 16'sd 19131) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11049) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14146) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19111) * $signed(input_fmap_173[7:0]) +
	( 16'sd 28161) * $signed(input_fmap_174[7:0]) +
	( 13'sd 2337) * $signed(input_fmap_175[7:0]) +
	( 14'sd 6047) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6531) * $signed(input_fmap_177[7:0]) +
	( 16'sd 24992) * $signed(input_fmap_178[7:0]) +
	( 15'sd 13967) * $signed(input_fmap_179[7:0]) +
	( 12'sd 1764) * $signed(input_fmap_180[7:0]) +
	( 16'sd 19038) * $signed(input_fmap_181[7:0]) +
	( 15'sd 16120) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25526) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_184[7:0]) +
	( 13'sd 2102) * $signed(input_fmap_185[7:0]) +
	( 14'sd 5324) * $signed(input_fmap_186[7:0]) +
	( 15'sd 15140) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2187) * $signed(input_fmap_188[7:0]) +
	( 8'sd 76) * $signed(input_fmap_189[7:0]) +
	( 15'sd 15667) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32254) * $signed(input_fmap_191[7:0]) +
	( 16'sd 26571) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20424) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18445) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24733) * $signed(input_fmap_197[7:0]) +
	( 15'sd 13744) * $signed(input_fmap_198[7:0]) +
	( 16'sd 21164) * $signed(input_fmap_199[7:0]) +
	( 16'sd 27575) * $signed(input_fmap_200[7:0]) +
	( 16'sd 19773) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19816) * $signed(input_fmap_202[7:0]) +
	( 16'sd 26853) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6473) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18690) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6757) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18801) * $signed(input_fmap_207[7:0]) +
	( 11'sd 720) * $signed(input_fmap_208[7:0]) +
	( 16'sd 32561) * $signed(input_fmap_209[7:0]) +
	( 16'sd 20104) * $signed(input_fmap_210[7:0]) +
	( 15'sd 16332) * $signed(input_fmap_211[7:0]) +
	( 15'sd 10292) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24217) * $signed(input_fmap_213[7:0]) +
	( 14'sd 5030) * $signed(input_fmap_214[7:0]) +
	( 14'sd 8158) * $signed(input_fmap_215[7:0]) +
	( 14'sd 8082) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17605) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_218[7:0]) +
	( 16'sd 25076) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13339) * $signed(input_fmap_220[7:0]) +
	( 16'sd 31003) * $signed(input_fmap_221[7:0]) +
	( 14'sd 7287) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14987) * $signed(input_fmap_223[7:0]) +
	( 16'sd 20466) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13873) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30886) * $signed(input_fmap_226[7:0]) +
	( 12'sd 1166) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19169) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20755) * $signed(input_fmap_229[7:0]) +
	( 16'sd 24169) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17817) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29432) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19748) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21944) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5020) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20801) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17391) * $signed(input_fmap_238[7:0]) +
	( 14'sd 7718) * $signed(input_fmap_239[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_240[7:0]) +
	( 15'sd 8676) * $signed(input_fmap_241[7:0]) +
	( 15'sd 13127) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22877) * $signed(input_fmap_243[7:0]) +
	( 16'sd 23999) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6760) * $signed(input_fmap_245[7:0]) +
	( 14'sd 4192) * $signed(input_fmap_246[7:0]) +
	( 16'sd 16415) * $signed(input_fmap_247[7:0]) +
	( 15'sd 14598) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17636) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12478) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7763) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20067) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_253[7:0]) +
	( 15'sd 12595) * $signed(input_fmap_254[7:0]) +
	( 16'sd 31011) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_51;
assign conv_mac_51 = 
	( 12'sd 1555) * $signed(input_fmap_0[7:0]) +
	( 11'sd 641) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9858) * $signed(input_fmap_2[7:0]) +
	( 10'sd 487) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29009) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14127) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6328) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10491) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2103) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18762) * $signed(input_fmap_9[7:0]) +
	( 11'sd 830) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18041) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25866) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32100) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26914) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26328) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27863) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17566) * $signed(input_fmap_17[7:0]) +
	( 8'sd 109) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12862) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10685) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25357) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21549) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30492) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20545) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30533) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3569) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14763) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2785) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17750) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21017) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31295) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19764) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19351) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5460) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5365) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8430) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5856) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7289) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20656) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19523) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19466) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2070) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24017) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19834) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22598) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32765) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18798) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9588) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14002) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2178) * $signed(input_fmap_54[7:0]) +
	( 13'sd 4052) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20853) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10372) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8708) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1591) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12448) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26518) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10414) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19529) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6795) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15907) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11861) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20156) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22514) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13467) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24742) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11177) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6963) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4704) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11270) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12898) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27043) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16906) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10497) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21960) * $signed(input_fmap_90[7:0]) +
	( 15'sd 16176) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2863) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5546) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24212) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16546) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11641) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9567) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25723) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22992) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8483) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24491) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19586) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31884) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5611) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3639) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25304) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30681) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2847) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10918) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18741) * $signed(input_fmap_111[7:0]) +
	( 14'sd 8161) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29265) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4343) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10533) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19522) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25708) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23760) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16948) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30393) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29984) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25058) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28095) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5922) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29159) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10457) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21565) * $signed(input_fmap_127[7:0]) +
	( 16'sd 22656) * $signed(input_fmap_128[7:0]) +
	( 16'sd 25044) * $signed(input_fmap_129[7:0]) +
	( 15'sd 13184) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13127) * $signed(input_fmap_131[7:0]) +
	( 16'sd 21675) * $signed(input_fmap_132[7:0]) +
	( 16'sd 25557) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21092) * $signed(input_fmap_134[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7286) * $signed(input_fmap_136[7:0]) +
	( 13'sd 2886) * $signed(input_fmap_137[7:0]) +
	( 16'sd 21474) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18162) * $signed(input_fmap_139[7:0]) +
	( 16'sd 23959) * $signed(input_fmap_140[7:0]) +
	( 15'sd 11300) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19268) * $signed(input_fmap_142[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31315) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23314) * $signed(input_fmap_145[7:0]) +
	( 14'sd 5976) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8941) * $signed(input_fmap_147[7:0]) +
	( 16'sd 16591) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18452) * $signed(input_fmap_149[7:0]) +
	( 13'sd 3697) * $signed(input_fmap_150[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2441) * $signed(input_fmap_152[7:0]) +
	( 16'sd 16895) * $signed(input_fmap_153[7:0]) +
	( 15'sd 9642) * $signed(input_fmap_154[7:0]) +
	( 16'sd 25467) * $signed(input_fmap_155[7:0]) +
	( 15'sd 8883) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23652) * $signed(input_fmap_157[7:0]) +
	( 14'sd 5272) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6139) * $signed(input_fmap_159[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28429) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13412) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27202) * $signed(input_fmap_163[7:0]) +
	( 16'sd 32414) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12111) * $signed(input_fmap_165[7:0]) +
	( 14'sd 6551) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20617) * $signed(input_fmap_167[7:0]) +
	( 15'sd 13668) * $signed(input_fmap_168[7:0]) +
	( 15'sd 13472) * $signed(input_fmap_169[7:0]) +
	( 16'sd 19977) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4686) * $signed(input_fmap_172[7:0]) +
	( 15'sd 10338) * $signed(input_fmap_173[7:0]) +
	( 15'sd 9549) * $signed(input_fmap_174[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_175[7:0]) +
	( 14'sd 6058) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7828) * $signed(input_fmap_177[7:0]) +
	( 16'sd 21682) * $signed(input_fmap_178[7:0]) +
	( 10'sd 387) * $signed(input_fmap_179[7:0]) +
	( 16'sd 19889) * $signed(input_fmap_180[7:0]) +
	( 15'sd 14687) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17970) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31810) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3576) * $signed(input_fmap_185[7:0]) +
	( 14'sd 7052) * $signed(input_fmap_186[7:0]) +
	( 15'sd 10680) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12153) * $signed(input_fmap_188[7:0]) +
	( 15'sd 13805) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27046) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5600) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15138) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15732) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27728) * $signed(input_fmap_194[7:0]) +
	( 13'sd 2488) * $signed(input_fmap_195[7:0]) +
	( 12'sd 1230) * $signed(input_fmap_196[7:0]) +
	( 14'sd 7592) * $signed(input_fmap_197[7:0]) +
	( 16'sd 31765) * $signed(input_fmap_198[7:0]) +
	( 16'sd 32259) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5048) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12101) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17900) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25242) * $signed(input_fmap_203[7:0]) +
	( 16'sd 31062) * $signed(input_fmap_204[7:0]) +
	( 14'sd 7806) * $signed(input_fmap_205[7:0]) +
	( 16'sd 19880) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3005) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17296) * $signed(input_fmap_208[7:0]) +
	( 16'sd 32680) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3610) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5236) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17199) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5946) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31032) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22375) * $signed(input_fmap_215[7:0]) +
	( 15'sd 13773) * $signed(input_fmap_216[7:0]) +
	( 16'sd 31267) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21257) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_219[7:0]) +
	( 14'sd 7546) * $signed(input_fmap_220[7:0]) +
	( 16'sd 31544) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28423) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14250) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1046) * $signed(input_fmap_224[7:0]) +
	( 16'sd 16622) * $signed(input_fmap_225[7:0]) +
	( 14'sd 4488) * $signed(input_fmap_226[7:0]) +
	( 16'sd 29084) * $signed(input_fmap_227[7:0]) +
	( 14'sd 7736) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6828) * $signed(input_fmap_229[7:0]) +
	( 13'sd 4009) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10132) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15360) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11134) * $signed(input_fmap_233[7:0]) +
	( 15'sd 11657) * $signed(input_fmap_234[7:0]) +
	( 15'sd 13455) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5550) * $signed(input_fmap_236[7:0]) +
	( 15'sd 15811) * $signed(input_fmap_237[7:0]) +
	( 15'sd 11345) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23020) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26911) * $signed(input_fmap_240[7:0]) +
	( 16'sd 28790) * $signed(input_fmap_241[7:0]) +
	( 16'sd 32592) * $signed(input_fmap_242[7:0]) +
	( 15'sd 15814) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6651) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3218) * $signed(input_fmap_245[7:0]) +
	( 15'sd 13585) * $signed(input_fmap_246[7:0]) +
	( 16'sd 31583) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32264) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14579) * $signed(input_fmap_249[7:0]) +
	( 16'sd 28978) * $signed(input_fmap_250[7:0]) +
	( 12'sd 1630) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4472) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2856) * $signed(input_fmap_253[7:0]) +
	( 15'sd 12337) * $signed(input_fmap_254[7:0]) +
	( 16'sd 18336) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_52;
assign conv_mac_52 = 
	( 16'sd 19867) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2786) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19580) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9508) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14204) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22697) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24136) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1129) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14669) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28492) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12111) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5082) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28114) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28818) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16036) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14284) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13719) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16916) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23375) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25256) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19265) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24089) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28157) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29621) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21987) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6534) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5115) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4322) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12683) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4477) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7484) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6984) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23573) * $signed(input_fmap_36[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24184) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13910) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28048) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8353) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21915) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3766) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4826) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22921) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16387) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2521) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11944) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30158) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10717) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11518) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20538) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13596) * $signed(input_fmap_54[7:0]) +
	( 6'sd 31) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10580) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29671) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22848) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1595) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14201) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9874) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29483) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17059) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25322) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9012) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16095) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26351) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25139) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8963) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19199) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6999) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29844) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2693) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3422) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32701) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32031) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12543) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15374) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21238) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21241) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6768) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7013) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27431) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7828) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7256) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19735) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24010) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22277) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9666) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19229) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9276) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25352) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_94[7:0]) +
	( 11'sd 568) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16959) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7099) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32447) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19529) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18311) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16529) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15589) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4615) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9329) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22430) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9333) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29475) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31737) * $signed(input_fmap_109[7:0]) +
	( 11'sd 614) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19107) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8831) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29747) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20566) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30317) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10808) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23602) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31612) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23001) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9449) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15186) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20957) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31019) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21994) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22765) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31100) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17842) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24082) * $signed(input_fmap_129[7:0]) +
	( 16'sd 29640) * $signed(input_fmap_130[7:0]) +
	( 14'sd 8082) * $signed(input_fmap_131[7:0]) +
	( 16'sd 17759) * $signed(input_fmap_132[7:0]) +
	( 13'sd 3167) * $signed(input_fmap_133[7:0]) +
	( 16'sd 28656) * $signed(input_fmap_134[7:0]) +
	( 15'sd 12545) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21602) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15077) * $signed(input_fmap_137[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_138[7:0]) +
	( 16'sd 19964) * $signed(input_fmap_139[7:0]) +
	( 13'sd 2198) * $signed(input_fmap_140[7:0]) +
	( 16'sd 27667) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31876) * $signed(input_fmap_142[7:0]) +
	( 11'sd 886) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28103) * $signed(input_fmap_144[7:0]) +
	( 16'sd 24176) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7543) * $signed(input_fmap_146[7:0]) +
	( 12'sd 2024) * $signed(input_fmap_147[7:0]) +
	( 16'sd 32010) * $signed(input_fmap_148[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9249) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18389) * $signed(input_fmap_151[7:0]) +
	( 16'sd 19443) * $signed(input_fmap_152[7:0]) +
	( 14'sd 7063) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30159) * $signed(input_fmap_154[7:0]) +
	( 16'sd 32714) * $signed(input_fmap_155[7:0]) +
	( 12'sd 1041) * $signed(input_fmap_156[7:0]) +
	( 16'sd 19104) * $signed(input_fmap_157[7:0]) +
	( 16'sd 31788) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4875) * $signed(input_fmap_159[7:0]) +
	( 15'sd 14504) * $signed(input_fmap_160[7:0]) +
	( 15'sd 10401) * $signed(input_fmap_161[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_162[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11900) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11039) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19469) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31963) * $signed(input_fmap_167[7:0]) +
	( 16'sd 24595) * $signed(input_fmap_168[7:0]) +
	( 15'sd 15113) * $signed(input_fmap_169[7:0]) +
	( 11'sd 815) * $signed(input_fmap_170[7:0]) +
	( 15'sd 10613) * $signed(input_fmap_171[7:0]) +
	( 16'sd 29343) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23224) * $signed(input_fmap_173[7:0]) +
	( 15'sd 12622) * $signed(input_fmap_174[7:0]) +
	( 16'sd 18537) * $signed(input_fmap_175[7:0]) +
	( 15'sd 8194) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19785) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32348) * $signed(input_fmap_178[7:0]) +
	( 14'sd 7417) * $signed(input_fmap_179[7:0]) +
	( 14'sd 5283) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11058) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26396) * $signed(input_fmap_182[7:0]) +
	( 16'sd 31740) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26811) * $signed(input_fmap_184[7:0]) +
	( 13'sd 2939) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2337) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_188[7:0]) +
	( 10'sd 319) * $signed(input_fmap_189[7:0]) +
	( 16'sd 29523) * $signed(input_fmap_190[7:0]) +
	( 15'sd 16021) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31121) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29499) * $signed(input_fmap_193[7:0]) +
	( 15'sd 13128) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19592) * $signed(input_fmap_195[7:0]) +
	( 14'sd 4572) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32013) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1045) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3936) * $signed(input_fmap_200[7:0]) +
	( 16'sd 24792) * $signed(input_fmap_201[7:0]) +
	( 16'sd 22060) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30743) * $signed(input_fmap_203[7:0]) +
	( 12'sd 1414) * $signed(input_fmap_204[7:0]) +
	( 15'sd 10030) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9716) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18790) * $signed(input_fmap_207[7:0]) +
	( 14'sd 5052) * $signed(input_fmap_208[7:0]) +
	( 14'sd 6501) * $signed(input_fmap_209[7:0]) +
	( 15'sd 14829) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6294) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1471) * $signed(input_fmap_212[7:0]) +
	( 14'sd 7955) * $signed(input_fmap_213[7:0]) +
	( 15'sd 8483) * $signed(input_fmap_214[7:0]) +
	( 16'sd 19974) * $signed(input_fmap_215[7:0]) +
	( 14'sd 6592) * $signed(input_fmap_216[7:0]) +
	( 13'sd 3515) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_218[7:0]) +
	( 12'sd 1788) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26588) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6187) * $signed(input_fmap_221[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_222[7:0]) +
	( 14'sd 4279) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6592) * $signed(input_fmap_224[7:0]) +
	( 15'sd 8546) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10782) * $signed(input_fmap_226[7:0]) +
	( 16'sd 29636) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22197) * $signed(input_fmap_228[7:0]) +
	( 13'sd 2693) * $signed(input_fmap_229[7:0]) +
	( 14'sd 4218) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7270) * $signed(input_fmap_231[7:0]) +
	( 15'sd 16294) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24961) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14458) * $signed(input_fmap_234[7:0]) +
	( 16'sd 16469) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28431) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28798) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3257) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9754) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1309) * $signed(input_fmap_240[7:0]) +
	( 16'sd 28176) * $signed(input_fmap_241[7:0]) +
	( 15'sd 12246) * $signed(input_fmap_242[7:0]) +
	( 14'sd 4705) * $signed(input_fmap_243[7:0]) +
	( 14'sd 7777) * $signed(input_fmap_244[7:0]) +
	( 12'sd 1360) * $signed(input_fmap_245[7:0]) +
	( 14'sd 4471) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8982) * $signed(input_fmap_247[7:0]) +
	( 16'sd 23413) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25166) * $signed(input_fmap_249[7:0]) +
	( 12'sd 1747) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18675) * $signed(input_fmap_251[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5675) * $signed(input_fmap_253[7:0]) +
	( 14'sd 4501) * $signed(input_fmap_254[7:0]) +
	( 16'sd 28566) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_53;
assign conv_mac_53 = 
	( 16'sd 29090) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7814) * $signed(input_fmap_1[7:0]) +
	( 13'sd 4023) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27168) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1656) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10213) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9195) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11400) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3823) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24655) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2923) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1880) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3597) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23115) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26703) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14036) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26858) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10137) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25383) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20510) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14435) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6753) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30579) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6316) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9784) * $signed(input_fmap_25[7:0]) +
	( 13'sd 2445) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20243) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3421) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10509) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25610) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1132) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30416) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19451) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28334) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13551) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3051) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9503) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31182) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30621) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23193) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29580) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26891) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24194) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13229) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31844) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10170) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25262) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17787) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8219) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5639) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28106) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10576) * $signed(input_fmap_58[7:0]) +
	( 4'sd 6) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28282) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25698) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28280) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10401) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24346) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17367) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20872) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5010) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10858) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_69[7:0]) +
	( 11'sd 825) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8854) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26370) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15986) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21864) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31886) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31179) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4817) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4472) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32549) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27846) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7045) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15914) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3336) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9423) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9861) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1802) * $signed(input_fmap_88[7:0]) +
	( 11'sd 607) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9604) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19468) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32751) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5778) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9523) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23231) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27850) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28659) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29084) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13445) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3005) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2811) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2490) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30755) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12914) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32652) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5989) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6914) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22089) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7257) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26809) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3614) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31478) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21494) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18592) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20377) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9513) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1113) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8339) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9680) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19938) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21832) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32715) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26158) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29886) * $signed(input_fmap_127[7:0]) +
	( 12'sd 1838) * $signed(input_fmap_128[7:0]) +
	( 13'sd 2999) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31679) * $signed(input_fmap_130[7:0]) +
	( 16'sd 26255) * $signed(input_fmap_131[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12427) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11958) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17251) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13383) * $signed(input_fmap_137[7:0]) +
	( 15'sd 13908) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18439) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1966) * $signed(input_fmap_140[7:0]) +
	( 14'sd 7612) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_142[7:0]) +
	( 15'sd 9172) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13472) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7955) * $signed(input_fmap_145[7:0]) +
	( 16'sd 32707) * $signed(input_fmap_146[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17949) * $signed(input_fmap_148[7:0]) +
	( 12'sd 1677) * $signed(input_fmap_149[7:0]) +
	( 14'sd 7157) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14894) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20446) * $signed(input_fmap_152[7:0]) +
	( 15'sd 15681) * $signed(input_fmap_153[7:0]) +
	( 16'sd 17283) * $signed(input_fmap_154[7:0]) +
	( 14'sd 4655) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15155) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11016) * $signed(input_fmap_157[7:0]) +
	( 15'sd 10676) * $signed(input_fmap_158[7:0]) +
	( 16'sd 30989) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22326) * $signed(input_fmap_160[7:0]) +
	( 16'sd 18697) * $signed(input_fmap_161[7:0]) +
	( 15'sd 9745) * $signed(input_fmap_162[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10290) * $signed(input_fmap_164[7:0]) +
	( 16'sd 24721) * $signed(input_fmap_165[7:0]) +
	( 15'sd 14861) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24039) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14418) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17478) * $signed(input_fmap_169[7:0]) +
	( 16'sd 19440) * $signed(input_fmap_170[7:0]) +
	( 16'sd 22010) * $signed(input_fmap_171[7:0]) +
	( 16'sd 29927) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12736) * $signed(input_fmap_173[7:0]) +
	( 13'sd 2288) * $signed(input_fmap_174[7:0]) +
	( 16'sd 26365) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_176[7:0]) +
	( 15'sd 12903) * $signed(input_fmap_177[7:0]) +
	( 16'sd 24105) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6775) * $signed(input_fmap_180[7:0]) +
	( 16'sd 27889) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6830) * $signed(input_fmap_182[7:0]) +
	( 15'sd 10539) * $signed(input_fmap_183[7:0]) +
	( 14'sd 4974) * $signed(input_fmap_184[7:0]) +
	( 16'sd 23667) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12576) * $signed(input_fmap_186[7:0]) +
	( 15'sd 14916) * $signed(input_fmap_187[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19087) * $signed(input_fmap_189[7:0]) +
	( 13'sd 2621) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26819) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27886) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29515) * $signed(input_fmap_193[7:0]) +
	( 14'sd 6648) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17261) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17169) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26839) * $signed(input_fmap_197[7:0]) +
	( 16'sd 30814) * $signed(input_fmap_198[7:0]) +
	( 14'sd 4284) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3907) * $signed(input_fmap_200[7:0]) +
	( 15'sd 14996) * $signed(input_fmap_201[7:0]) +
	( 10'sd 348) * $signed(input_fmap_202[7:0]) +
	( 16'sd 26589) * $signed(input_fmap_203[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28514) * $signed(input_fmap_205[7:0]) +
	( 14'sd 5360) * $signed(input_fmap_206[7:0]) +
	( 16'sd 25131) * $signed(input_fmap_207[7:0]) +
	( 14'sd 5450) * $signed(input_fmap_208[7:0]) +
	( 15'sd 9101) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_210[7:0]) +
	( 15'sd 13203) * $signed(input_fmap_211[7:0]) +
	( 15'sd 8752) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28185) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17468) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25027) * $signed(input_fmap_215[7:0]) +
	( 15'sd 10477) * $signed(input_fmap_216[7:0]) +
	( 15'sd 13782) * $signed(input_fmap_217[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17488) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14050) * $signed(input_fmap_220[7:0]) +
	( 16'sd 22869) * $signed(input_fmap_221[7:0]) +
	( 16'sd 27506) * $signed(input_fmap_222[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_223[7:0]) +
	( 16'sd 24409) * $signed(input_fmap_224[7:0]) +
	( 15'sd 12804) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14395) * $signed(input_fmap_226[7:0]) +
	( 15'sd 15564) * $signed(input_fmap_227[7:0]) +
	( 14'sd 6894) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_229[7:0]) +
	( 15'sd 10675) * $signed(input_fmap_230[7:0]) +
	( 15'sd 15379) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20937) * $signed(input_fmap_232[7:0]) +
	( 16'sd 22568) * $signed(input_fmap_233[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21647) * $signed(input_fmap_235[7:0]) +
	( 15'sd 15039) * $signed(input_fmap_236[7:0]) +
	( 16'sd 31574) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12238) * $signed(input_fmap_238[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_239[7:0]) +
	( 10'sd 313) * $signed(input_fmap_240[7:0]) +
	( 16'sd 19583) * $signed(input_fmap_241[7:0]) +
	( 16'sd 19907) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23902) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19143) * $signed(input_fmap_245[7:0]) +
	( 16'sd 21042) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13517) * $signed(input_fmap_247[7:0]) +
	( 6'sd 31) * $signed(input_fmap_248[7:0]) +
	( 14'sd 5661) * $signed(input_fmap_249[7:0]) +
	( 15'sd 13873) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13040) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2691) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29181) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_254[7:0]) +
	( 16'sd 25732) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_54;
assign conv_mac_54 = 
	( 16'sd 30962) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17174) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17542) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20607) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25189) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1361) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26081) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25596) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29948) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29051) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12459) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11113) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10970) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14766) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10372) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4829) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3080) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8648) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4692) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24028) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10861) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6611) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13180) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14415) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28941) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15077) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30584) * $signed(input_fmap_32[7:0]) +
	( 11'sd 1015) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7347) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17530) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30735) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13019) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20105) * $signed(input_fmap_38[7:0]) +
	( 11'sd 840) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21196) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21700) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8673) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16914) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9257) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14342) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21365) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29075) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28025) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31360) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10630) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21536) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14229) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11830) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20886) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18351) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9198) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15316) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30799) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16261) * $signed(input_fmap_59[7:0]) +
	( 9'sd 185) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9216) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14754) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17971) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29091) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21912) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24812) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13821) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12456) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7870) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32100) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12199) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12189) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13339) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32730) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15925) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2662) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10158) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26180) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23425) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4539) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32136) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2380) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31477) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32754) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17013) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4775) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3153) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2680) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22571) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24584) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30031) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27071) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9247) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20968) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12359) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13175) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12189) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28916) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18967) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20340) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1054) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12898) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1561) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22883) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25862) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30443) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16947) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31284) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6548) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6006) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32412) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31594) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24829) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15378) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17697) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21823) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29567) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19181) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17046) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7575) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18458) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5540) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18178) * $signed(input_fmap_132[7:0]) +
	( 16'sd 32525) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24919) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19989) * $signed(input_fmap_135[7:0]) +
	( 16'sd 27634) * $signed(input_fmap_136[7:0]) +
	( 14'sd 7367) * $signed(input_fmap_137[7:0]) +
	( 14'sd 5602) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27920) * $signed(input_fmap_139[7:0]) +
	( 16'sd 25107) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5190) * $signed(input_fmap_141[7:0]) +
	( 14'sd 5979) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1928) * $signed(input_fmap_143[7:0]) +
	( 15'sd 8348) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21494) * $signed(input_fmap_145[7:0]) +
	( 16'sd 28404) * $signed(input_fmap_146[7:0]) +
	( 12'sd 1044) * $signed(input_fmap_147[7:0]) +
	( 16'sd 24838) * $signed(input_fmap_148[7:0]) +
	( 16'sd 29736) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25545) * $signed(input_fmap_150[7:0]) +
	( 8'sd 113) * $signed(input_fmap_151[7:0]) +
	( 15'sd 16075) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17749) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22122) * $signed(input_fmap_154[7:0]) +
	( 16'sd 31378) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7197) * $signed(input_fmap_156[7:0]) +
	( 15'sd 9001) * $signed(input_fmap_157[7:0]) +
	( 16'sd 19745) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26258) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_160[7:0]) +
	( 16'sd 21830) * $signed(input_fmap_161[7:0]) +
	( 16'sd 23277) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27022) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_164[7:0]) +
	( 16'sd 20560) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_166[7:0]) +
	( 16'sd 28231) * $signed(input_fmap_167[7:0]) +
	( 16'sd 31267) * $signed(input_fmap_168[7:0]) +
	( 16'sd 22951) * $signed(input_fmap_169[7:0]) +
	( 16'sd 16729) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18931) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1579) * $signed(input_fmap_172[7:0]) +
	( 13'sd 3126) * $signed(input_fmap_173[7:0]) +
	( 14'sd 4769) * $signed(input_fmap_174[7:0]) +
	( 15'sd 14723) * $signed(input_fmap_175[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_176[7:0]) +
	( 15'sd 13559) * $signed(input_fmap_177[7:0]) +
	( 15'sd 13409) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20552) * $signed(input_fmap_179[7:0]) +
	( 10'sd 422) * $signed(input_fmap_180[7:0]) +
	( 15'sd 8893) * $signed(input_fmap_181[7:0]) +
	( 16'sd 24275) * $signed(input_fmap_182[7:0]) +
	( 16'sd 18194) * $signed(input_fmap_183[7:0]) +
	( 12'sd 1462) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7875) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3405) * $signed(input_fmap_186[7:0]) +
	( 16'sd 19487) * $signed(input_fmap_187[7:0]) +
	( 15'sd 8804) * $signed(input_fmap_188[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_189[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_190[7:0]) +
	( 15'sd 15694) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12649) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26304) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26366) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19019) * $signed(input_fmap_195[7:0]) +
	( 13'sd 2552) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14455) * $signed(input_fmap_197[7:0]) +
	( 16'sd 21425) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12570) * $signed(input_fmap_199[7:0]) +
	( 16'sd 22187) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13486) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11178) * $signed(input_fmap_202[7:0]) +
	( 15'sd 8562) * $signed(input_fmap_203[7:0]) +
	( 16'sd 16412) * $signed(input_fmap_204[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_206[7:0]) +
	( 13'sd 2297) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17780) * $signed(input_fmap_208[7:0]) +
	( 16'sd 31510) * $signed(input_fmap_209[7:0]) +
	( 15'sd 8362) * $signed(input_fmap_210[7:0]) +
	( 16'sd 31475) * $signed(input_fmap_211[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2132) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30751) * $signed(input_fmap_214[7:0]) +
	( 11'sd 793) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4122) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25861) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_218[7:0]) +
	( 15'sd 8257) * $signed(input_fmap_219[7:0]) +
	( 14'sd 5526) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13904) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14487) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14260) * $signed(input_fmap_223[7:0]) +
	( 10'sd 360) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26053) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22738) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_227[7:0]) +
	( 16'sd 32530) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23864) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7642) * $signed(input_fmap_230[7:0]) +
	( 16'sd 32676) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29925) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21124) * $signed(input_fmap_233[7:0]) +
	( 15'sd 11917) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7080) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23492) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19454) * $signed(input_fmap_237[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_238[7:0]) +
	( 15'sd 11635) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18105) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18606) * $signed(input_fmap_241[7:0]) +
	( 14'sd 6497) * $signed(input_fmap_242[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_243[7:0]) +
	( 16'sd 21315) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7660) * $signed(input_fmap_245[7:0]) +
	( 14'sd 7111) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21263) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26637) * $signed(input_fmap_248[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_249[7:0]) +
	( 16'sd 27681) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28238) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3591) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9164) * $signed(input_fmap_254[7:0]) +
	( 16'sd 17857) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_55;
assign conv_mac_55 = 
	( 16'sd 23112) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25345) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5270) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29337) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27272) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31450) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17285) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17890) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26226) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28169) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26531) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32333) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32720) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2361) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23425) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5216) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15309) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26560) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17162) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28604) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27898) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2215) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18723) * $signed(input_fmap_23[7:0]) +
	( 10'sd 426) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31898) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21241) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1965) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8792) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27274) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_31[7:0]) +
	( 11'sd 693) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18980) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24234) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26483) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24085) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6117) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20248) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17754) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30066) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11554) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11409) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23113) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13931) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8229) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3958) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14555) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10817) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14974) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1469) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8752) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31777) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14654) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16555) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28582) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29396) * $signed(input_fmap_62[7:0]) +
	( 10'sd 299) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12410) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6990) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19509) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31711) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24274) * $signed(input_fmap_68[7:0]) +
	( 7'sd 34) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11634) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21450) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15483) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29954) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1332) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17838) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30807) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27572) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26648) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2713) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2558) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23977) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19637) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31438) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22722) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32390) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29762) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5334) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21015) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10776) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5644) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26545) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14520) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29411) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25015) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31009) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1501) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16963) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7247) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17319) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29297) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1037) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16877) * $signed(input_fmap_106[7:0]) +
	( 14'sd 8186) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15377) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14881) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16536) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21271) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4530) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4561) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16392) * $signed(input_fmap_115[7:0]) +
	( 11'sd 908) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2549) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13467) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9464) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24858) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1454) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14510) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11017) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4899) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4564) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8519) * $signed(input_fmap_127[7:0]) +
	( 14'sd 6680) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17857) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10665) * $signed(input_fmap_130[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_131[7:0]) +
	( 16'sd 31115) * $signed(input_fmap_132[7:0]) +
	( 16'sd 17629) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31694) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25558) * $signed(input_fmap_136[7:0]) +
	( 16'sd 28733) * $signed(input_fmap_137[7:0]) +
	( 16'sd 20794) * $signed(input_fmap_138[7:0]) +
	( 16'sd 19764) * $signed(input_fmap_139[7:0]) +
	( 16'sd 25214) * $signed(input_fmap_140[7:0]) +
	( 10'sd 256) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25816) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4238) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5571) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28138) * $signed(input_fmap_145[7:0]) +
	( 16'sd 23059) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14127) * $signed(input_fmap_147[7:0]) +
	( 16'sd 19119) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2064) * $signed(input_fmap_149[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_150[7:0]) +
	( 15'sd 15997) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31385) * $signed(input_fmap_152[7:0]) +
	( 16'sd 19785) * $signed(input_fmap_153[7:0]) +
	( 16'sd 28363) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23767) * $signed(input_fmap_155[7:0]) +
	( 14'sd 6788) * $signed(input_fmap_156[7:0]) +
	( 11'sd 580) * $signed(input_fmap_157[7:0]) +
	( 16'sd 23032) * $signed(input_fmap_158[7:0]) +
	( 16'sd 30166) * $signed(input_fmap_159[7:0]) +
	( 16'sd 16641) * $signed(input_fmap_160[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4843) * $signed(input_fmap_162[7:0]) +
	( 14'sd 7119) * $signed(input_fmap_163[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_164[7:0]) +
	( 16'sd 21888) * $signed(input_fmap_165[7:0]) +
	( 16'sd 21200) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17525) * $signed(input_fmap_167[7:0]) +
	( 16'sd 19005) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17335) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28491) * $signed(input_fmap_170[7:0]) +
	( 16'sd 21773) * $signed(input_fmap_171[7:0]) +
	( 15'sd 13379) * $signed(input_fmap_172[7:0]) +
	( 16'sd 24060) * $signed(input_fmap_173[7:0]) +
	( 11'sd 523) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_175[7:0]) +
	( 16'sd 32002) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7148) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_178[7:0]) +
	( 15'sd 11518) * $signed(input_fmap_179[7:0]) +
	( 13'sd 2664) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25275) * $signed(input_fmap_181[7:0]) +
	( 15'sd 11271) * $signed(input_fmap_182[7:0]) +
	( 11'sd 741) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14359) * $signed(input_fmap_184[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_185[7:0]) +
	( 16'sd 20254) * $signed(input_fmap_186[7:0]) +
	( 14'sd 7353) * $signed(input_fmap_187[7:0]) +
	( 15'sd 11479) * $signed(input_fmap_188[7:0]) +
	( 16'sd 27072) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13778) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23801) * $signed(input_fmap_191[7:0]) +
	( 15'sd 8803) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19320) * $signed(input_fmap_193[7:0]) +
	( 16'sd 32631) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27092) * $signed(input_fmap_195[7:0]) +
	( 13'sd 3208) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26130) * $signed(input_fmap_197[7:0]) +
	( 14'sd 4365) * $signed(input_fmap_198[7:0]) +
	( 15'sd 13345) * $signed(input_fmap_199[7:0]) +
	( 16'sd 30225) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22014) * $signed(input_fmap_201[7:0]) +
	( 16'sd 24225) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13230) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6310) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24996) * $signed(input_fmap_205[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_206[7:0]) +
	( 16'sd 22669) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4457) * $signed(input_fmap_208[7:0]) +
	( 14'sd 6055) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10996) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15743) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26286) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5256) * $signed(input_fmap_213[7:0]) +
	( 16'sd 32405) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_215[7:0]) +
	( 15'sd 15229) * $signed(input_fmap_216[7:0]) +
	( 16'sd 28330) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21840) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_220[7:0]) +
	( 15'sd 10549) * $signed(input_fmap_221[7:0]) +
	( 16'sd 21715) * $signed(input_fmap_222[7:0]) +
	( 15'sd 13631) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6240) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14274) * $signed(input_fmap_225[7:0]) +
	( 16'sd 16799) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5565) * $signed(input_fmap_227[7:0]) +
	( 15'sd 16084) * $signed(input_fmap_228[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_229[7:0]) +
	( 16'sd 26844) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13562) * $signed(input_fmap_231[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_232[7:0]) +
	( 14'sd 4946) * $signed(input_fmap_233[7:0]) +
	( 13'sd 2507) * $signed(input_fmap_234[7:0]) +
	( 16'sd 31973) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2872) * $signed(input_fmap_236[7:0]) +
	( 16'sd 22938) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22104) * $signed(input_fmap_238[7:0]) +
	( 11'sd 748) * $signed(input_fmap_239[7:0]) +
	( 16'sd 28428) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20256) * $signed(input_fmap_241[7:0]) +
	( 16'sd 21645) * $signed(input_fmap_242[7:0]) +
	( 16'sd 16887) * $signed(input_fmap_243[7:0]) +
	( 15'sd 16003) * $signed(input_fmap_244[7:0]) +
	( 15'sd 9127) * $signed(input_fmap_245[7:0]) +
	( 15'sd 8641) * $signed(input_fmap_246[7:0]) +
	( 13'sd 2609) * $signed(input_fmap_247[7:0]) +
	( 15'sd 9513) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24041) * $signed(input_fmap_249[7:0]) +
	( 10'sd 382) * $signed(input_fmap_250[7:0]) +
	( 16'sd 23212) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2418) * $signed(input_fmap_252[7:0]) +
	( 16'sd 20786) * $signed(input_fmap_253[7:0]) +
	( 14'sd 7615) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26416) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_56;
assign conv_mac_56 = 
	( 16'sd 30146) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26960) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1371) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23855) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24559) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22286) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3989) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7116) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16046) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18142) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8896) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7191) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20676) * $signed(input_fmap_14[7:0]) +
	( 10'sd 432) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18524) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4437) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9310) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7796) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26416) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25806) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16746) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5009) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29658) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30274) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28499) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18494) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25075) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6981) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25757) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20779) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26875) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17443) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15630) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16911) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25071) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17512) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17652) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_41[7:0]) +
	( 9'sd 246) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25653) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21037) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18555) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19930) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4836) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27823) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32138) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12782) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7184) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19032) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14824) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10373) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24813) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3475) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17516) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7680) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21247) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25849) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31352) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4333) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17143) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14387) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4131) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31565) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16568) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24403) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17615) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18394) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23674) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6414) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_77[7:0]) +
	( 12'sd 1654) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6324) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17399) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14508) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17159) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28180) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27513) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24939) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23982) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11285) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21388) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21000) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16951) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14732) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26645) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20505) * $signed(input_fmap_96[7:0]) +
	( 11'sd 561) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22798) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19270) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13146) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4927) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22700) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15535) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26360) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24621) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24337) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12940) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24123) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17321) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12714) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17789) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26076) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32165) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18982) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25556) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1036) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13699) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23029) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23172) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7992) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15524) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5399) * $signed(input_fmap_123[7:0]) +
	( 11'sd 519) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4734) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29151) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30311) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10420) * $signed(input_fmap_129[7:0]) +
	( 16'sd 23449) * $signed(input_fmap_130[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_131[7:0]) +
	( 14'sd 4831) * $signed(input_fmap_132[7:0]) +
	( 14'sd 4508) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31674) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_135[7:0]) +
	( 16'sd 20326) * $signed(input_fmap_136[7:0]) +
	( 15'sd 8304) * $signed(input_fmap_137[7:0]) +
	( 16'sd 28320) * $signed(input_fmap_138[7:0]) +
	( 11'sd 904) * $signed(input_fmap_139[7:0]) +
	( 16'sd 23642) * $signed(input_fmap_140[7:0]) +
	( 16'sd 25009) * $signed(input_fmap_141[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1128) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22019) * $signed(input_fmap_144[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29270) * $signed(input_fmap_146[7:0]) +
	( 14'sd 6085) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_148[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_149[7:0]) +
	( 16'sd 20280) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18848) * $signed(input_fmap_151[7:0]) +
	( 16'sd 26372) * $signed(input_fmap_152[7:0]) +
	( 10'sd 343) * $signed(input_fmap_153[7:0]) +
	( 15'sd 12786) * $signed(input_fmap_154[7:0]) +
	( 16'sd 31435) * $signed(input_fmap_155[7:0]) +
	( 14'sd 4578) * $signed(input_fmap_156[7:0]) +
	( 15'sd 8925) * $signed(input_fmap_157[7:0]) +
	( 16'sd 27224) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_160[7:0]) +
	( 16'sd 24003) * $signed(input_fmap_161[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_163[7:0]) +
	( 16'sd 27979) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30334) * $signed(input_fmap_165[7:0]) +
	( 14'sd 6116) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7857) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29132) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_169[7:0]) +
	( 14'sd 6810) * $signed(input_fmap_170[7:0]) +
	( 16'sd 22716) * $signed(input_fmap_171[7:0]) +
	( 16'sd 26532) * $signed(input_fmap_172[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11976) * $signed(input_fmap_174[7:0]) +
	( 16'sd 20085) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21655) * $signed(input_fmap_176[7:0]) +
	( 15'sd 11716) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1946) * $signed(input_fmap_178[7:0]) +
	( 16'sd 27804) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28276) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18973) * $signed(input_fmap_181[7:0]) +
	( 15'sd 13610) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27924) * $signed(input_fmap_183[7:0]) +
	( 14'sd 5321) * $signed(input_fmap_184[7:0]) +
	( 16'sd 30223) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2829) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1030) * $signed(input_fmap_187[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_188[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_189[7:0]) +
	( 13'sd 2413) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29577) * $signed(input_fmap_191[7:0]) +
	( 15'sd 9143) * $signed(input_fmap_192[7:0]) +
	( 16'sd 21828) * $signed(input_fmap_193[7:0]) +
	( 15'sd 10151) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1316) * $signed(input_fmap_195[7:0]) +
	( 16'sd 16811) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15229) * $signed(input_fmap_197[7:0]) +
	( 15'sd 8525) * $signed(input_fmap_198[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_199[7:0]) +
	( 16'sd 21349) * $signed(input_fmap_200[7:0]) +
	( 16'sd 20909) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_202[7:0]) +
	( 15'sd 14100) * $signed(input_fmap_203[7:0]) +
	( 16'sd 28991) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2884) * $signed(input_fmap_205[7:0]) +
	( 15'sd 15081) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12380) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8284) * $signed(input_fmap_208[7:0]) +
	( 16'sd 25459) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10430) * $signed(input_fmap_210[7:0]) +
	( 14'sd 7434) * $signed(input_fmap_211[7:0]) +
	( 14'sd 5883) * $signed(input_fmap_212[7:0]) +
	( 16'sd 31295) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1369) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25859) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20677) * $signed(input_fmap_216[7:0]) +
	( 16'sd 21753) * $signed(input_fmap_217[7:0]) +
	( 14'sd 4164) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12441) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25753) * $signed(input_fmap_220[7:0]) +
	( 14'sd 4354) * $signed(input_fmap_221[7:0]) +
	( 16'sd 32442) * $signed(input_fmap_222[7:0]) +
	( 16'sd 26118) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3797) * $signed(input_fmap_225[7:0]) +
	( 16'sd 21288) * $signed(input_fmap_226[7:0]) +
	( 15'sd 16090) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25094) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29167) * $signed(input_fmap_229[7:0]) +
	( 16'sd 24505) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1800) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18036) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11604) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13044) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_235[7:0]) +
	( 11'sd 853) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2869) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16530) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23654) * $signed(input_fmap_239[7:0]) +
	( 16'sd 24977) * $signed(input_fmap_240[7:0]) +
	( 15'sd 9716) * $signed(input_fmap_241[7:0]) +
	( 14'sd 6828) * $signed(input_fmap_242[7:0]) +
	( 15'sd 12752) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13742) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7344) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14330) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12667) * $signed(input_fmap_247[7:0]) +
	( 16'sd 24493) * $signed(input_fmap_248[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12772) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6655) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6488) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6209) * $signed(input_fmap_253[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_254[7:0]) +
	( 12'sd 2047) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_57;
assign conv_mac_57 = 
	( 16'sd 28532) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14568) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3954) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9917) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15765) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28403) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12110) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31269) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13137) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10784) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32163) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7322) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31935) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18684) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21664) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20105) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29510) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25371) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31254) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18144) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13806) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20522) * $signed(input_fmap_26[7:0]) +
	( 11'sd 695) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11811) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22107) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25544) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10685) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4242) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29628) * $signed(input_fmap_33[7:0]) +
	( 16'sd 32517) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27102) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6030) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8424) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20398) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7120) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6019) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23230) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4277) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1277) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13833) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7801) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8370) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5650) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21313) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14639) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7512) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2486) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16756) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15038) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15659) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32214) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27661) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17030) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30428) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5402) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10516) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18191) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4299) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19296) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15113) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10778) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18115) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27635) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11277) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16748) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13419) * $signed(input_fmap_79[7:0]) +
	( 11'sd 801) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16006) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11014) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14305) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15081) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30206) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4143) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8456) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9459) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7477) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31163) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27993) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8981) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17583) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10954) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24653) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17118) * $signed(input_fmap_97[7:0]) +
	( 6'sd 21) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18381) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24580) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23410) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12693) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9400) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10942) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18693) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32535) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4672) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6153) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2358) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23482) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5491) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13574) * $signed(input_fmap_116[7:0]) +
	( 10'sd 305) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8201) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9266) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24715) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13437) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28027) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31851) * $signed(input_fmap_124[7:0]) +
	( 10'sd 319) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22648) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27795) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9464) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5889) * $signed(input_fmap_129[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15573) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5330) * $signed(input_fmap_132[7:0]) +
	( 16'sd 32494) * $signed(input_fmap_133[7:0]) +
	( 15'sd 8398) * $signed(input_fmap_134[7:0]) +
	( 15'sd 16205) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7539) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12807) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9974) * $signed(input_fmap_138[7:0]) +
	( 15'sd 15658) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26968) * $signed(input_fmap_140[7:0]) +
	( 16'sd 27589) * $signed(input_fmap_141[7:0]) +
	( 10'sd 423) * $signed(input_fmap_142[7:0]) +
	( 15'sd 15742) * $signed(input_fmap_143[7:0]) +
	( 15'sd 10889) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9946) * $signed(input_fmap_146[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6733) * $signed(input_fmap_148[7:0]) +
	( 15'sd 13873) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27983) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23257) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30363) * $signed(input_fmap_152[7:0]) +
	( 16'sd 19905) * $signed(input_fmap_153[7:0]) +
	( 15'sd 8230) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27874) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28560) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6322) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4876) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20003) * $signed(input_fmap_159[7:0]) +
	( 13'sd 3563) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_161[7:0]) +
	( 16'sd 17150) * $signed(input_fmap_162[7:0]) +
	( 12'sd 1113) * $signed(input_fmap_163[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9456) * $signed(input_fmap_165[7:0]) +
	( 16'sd 24184) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26457) * $signed(input_fmap_167[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_168[7:0]) +
	( 15'sd 8748) * $signed(input_fmap_169[7:0]) +
	( 16'sd 30326) * $signed(input_fmap_170[7:0]) +
	( 15'sd 13527) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_172[7:0]) +
	( 14'sd 6833) * $signed(input_fmap_173[7:0]) +
	( 16'sd 17051) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21904) * $signed(input_fmap_175[7:0]) +
	( 9'sd 234) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29919) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15984) * $signed(input_fmap_178[7:0]) +
	( 15'sd 11797) * $signed(input_fmap_179[7:0]) +
	( 15'sd 12413) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3124) * $signed(input_fmap_181[7:0]) +
	( 16'sd 20594) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27016) * $signed(input_fmap_183[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_184[7:0]) +
	( 16'sd 28994) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6718) * $signed(input_fmap_186[7:0]) +
	( 14'sd 7509) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32490) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_189[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_190[7:0]) +
	( 14'sd 6023) * $signed(input_fmap_191[7:0]) +
	( 14'sd 8088) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_193[7:0]) +
	( 13'sd 4086) * $signed(input_fmap_194[7:0]) +
	( 16'sd 30509) * $signed(input_fmap_195[7:0]) +
	( 16'sd 18797) * $signed(input_fmap_196[7:0]) +
	( 16'sd 27118) * $signed(input_fmap_197[7:0]) +
	( 16'sd 26394) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_199[7:0]) +
	( 16'sd 21188) * $signed(input_fmap_200[7:0]) +
	( 15'sd 16022) * $signed(input_fmap_201[7:0]) +
	( 15'sd 10234) * $signed(input_fmap_202[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_205[7:0]) +
	( 16'sd 23958) * $signed(input_fmap_206[7:0]) +
	( 15'sd 10130) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18365) * $signed(input_fmap_208[7:0]) +
	( 15'sd 12316) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11206) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28171) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19930) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6385) * $signed(input_fmap_213[7:0]) +
	( 16'sd 32385) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7122) * $signed(input_fmap_215[7:0]) +
	( 16'sd 31444) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24857) * $signed(input_fmap_217[7:0]) +
	( 15'sd 15942) * $signed(input_fmap_218[7:0]) +
	( 16'sd 23200) * $signed(input_fmap_219[7:0]) +
	( 15'sd 12414) * $signed(input_fmap_220[7:0]) +
	( 16'sd 22293) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3148) * $signed(input_fmap_222[7:0]) +
	( 16'sd 20289) * $signed(input_fmap_223[7:0]) +
	( 14'sd 4851) * $signed(input_fmap_224[7:0]) +
	( 14'sd 8158) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31466) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20002) * $signed(input_fmap_227[7:0]) +
	( 14'sd 6364) * $signed(input_fmap_228[7:0]) +
	( 16'sd 22055) * $signed(input_fmap_229[7:0]) +
	( 13'sd 3664) * $signed(input_fmap_230[7:0]) +
	( 14'sd 5378) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14154) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28150) * $signed(input_fmap_233[7:0]) +
	( 16'sd 24186) * $signed(input_fmap_234[7:0]) +
	( 12'sd 1360) * $signed(input_fmap_235[7:0]) +
	( 16'sd 20005) * $signed(input_fmap_236[7:0]) +
	( 16'sd 26103) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12849) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9362) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31895) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32077) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29790) * $signed(input_fmap_242[7:0]) +
	( 16'sd 19810) * $signed(input_fmap_243[7:0]) +
	( 16'sd 21813) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30306) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17723) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_247[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_248[7:0]) +
	( 16'sd 31317) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24683) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4761) * $signed(input_fmap_251[7:0]) +
	( 16'sd 23108) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11792) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9453) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5826) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_58;
assign conv_mac_58 = 
	( 16'sd 17347) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32013) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28003) * $signed(input_fmap_2[7:0]) +
	( 15'sd 16164) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11205) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25570) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27609) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7217) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15549) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29307) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26011) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17821) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17922) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22672) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24327) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18961) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12376) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18104) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28233) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20926) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12859) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18676) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9770) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8780) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14009) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8417) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8293) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9897) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31664) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2261) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28219) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20331) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13200) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3864) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22341) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9140) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30559) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22182) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12058) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20236) * $signed(input_fmap_42[7:0]) +
	( 11'sd 905) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6675) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16082) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13774) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11403) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26718) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19668) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9584) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22402) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3046) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5868) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20780) * $signed(input_fmap_55[7:0]) +
	( 10'sd 307) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12201) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19522) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13124) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19173) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26407) * $signed(input_fmap_61[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2510) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27710) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17966) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3211) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14720) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5080) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30110) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17600) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22758) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29657) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26931) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16101) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6456) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30305) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18005) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8038) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32743) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5180) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21289) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22817) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31971) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7099) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16196) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22897) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6760) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29145) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16271) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22072) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9873) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19340) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13675) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11657) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23089) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26856) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16769) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24972) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20563) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18260) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13235) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31504) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27341) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13216) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19769) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25828) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20020) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31142) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3880) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4151) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32487) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6834) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29575) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19613) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25389) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23119) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25628) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18621) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1167) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13063) * $signed(input_fmap_126[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_127[7:0]) +
	( 12'sd 1468) * $signed(input_fmap_128[7:0]) +
	( 16'sd 29018) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18686) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_131[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_132[7:0]) +
	( 16'sd 24169) * $signed(input_fmap_133[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_134[7:0]) +
	( 11'sd 722) * $signed(input_fmap_135[7:0]) +
	( 16'sd 20115) * $signed(input_fmap_136[7:0]) +
	( 16'sd 20930) * $signed(input_fmap_137[7:0]) +
	( 15'sd 12912) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24744) * $signed(input_fmap_139[7:0]) +
	( 16'sd 32670) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12514) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31354) * $signed(input_fmap_142[7:0]) +
	( 13'sd 2610) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19433) * $signed(input_fmap_144[7:0]) +
	( 16'sd 20519) * $signed(input_fmap_145[7:0]) +
	( 16'sd 31779) * $signed(input_fmap_146[7:0]) +
	( 16'sd 26328) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17300) * $signed(input_fmap_148[7:0]) +
	( 16'sd 20550) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24637) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29918) * $signed(input_fmap_152[7:0]) +
	( 14'sd 5415) * $signed(input_fmap_153[7:0]) +
	( 16'sd 29517) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28708) * $signed(input_fmap_155[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_156[7:0]) +
	( 16'sd 28318) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18018) * $signed(input_fmap_158[7:0]) +
	( 16'sd 22258) * $signed(input_fmap_159[7:0]) +
	( 16'sd 25277) * $signed(input_fmap_160[7:0]) +
	( 14'sd 7894) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21198) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27312) * $signed(input_fmap_163[7:0]) +
	( 16'sd 28240) * $signed(input_fmap_164[7:0]) +
	( 15'sd 16314) * $signed(input_fmap_165[7:0]) +
	( 16'sd 29368) * $signed(input_fmap_166[7:0]) +
	( 16'sd 28600) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4597) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21652) * $signed(input_fmap_169[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_170[7:0]) +
	( 16'sd 26409) * $signed(input_fmap_171[7:0]) +
	( 16'sd 18242) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23136) * $signed(input_fmap_173[7:0]) +
	( 16'sd 25871) * $signed(input_fmap_174[7:0]) +
	( 16'sd 22463) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30060) * $signed(input_fmap_177[7:0]) +
	( 14'sd 7221) * $signed(input_fmap_178[7:0]) +
	( 15'sd 13793) * $signed(input_fmap_179[7:0]) +
	( 16'sd 22170) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6165) * $signed(input_fmap_181[7:0]) +
	( 16'sd 20870) * $signed(input_fmap_182[7:0]) +
	( 15'sd 8653) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31704) * $signed(input_fmap_184[7:0]) +
	( 16'sd 29709) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13660) * $signed(input_fmap_186[7:0]) +
	( 15'sd 14080) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_188[7:0]) +
	( 16'sd 16632) * $signed(input_fmap_189[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_190[7:0]) +
	( 12'sd 1485) * $signed(input_fmap_191[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26675) * $signed(input_fmap_193[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24439) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19615) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1721) * $signed(input_fmap_197[7:0]) +
	( 15'sd 11085) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1752) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_200[7:0]) +
	( 14'sd 4403) * $signed(input_fmap_201[7:0]) +
	( 16'sd 28385) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21229) * $signed(input_fmap_203[7:0]) +
	( 16'sd 18179) * $signed(input_fmap_204[7:0]) +
	( 16'sd 21466) * $signed(input_fmap_205[7:0]) +
	( 16'sd 24357) * $signed(input_fmap_206[7:0]) +
	( 13'sd 2112) * $signed(input_fmap_207[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_208[7:0]) +
	( 10'sd 497) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3034) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6976) * $signed(input_fmap_211[7:0]) +
	( 16'sd 22429) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24011) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14419) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10686) * $signed(input_fmap_215[7:0]) +
	( 16'sd 27391) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19650) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8761) * $signed(input_fmap_218[7:0]) +
	( 16'sd 18965) * $signed(input_fmap_219[7:0]) +
	( 15'sd 8592) * $signed(input_fmap_220[7:0]) +
	( 13'sd 2570) * $signed(input_fmap_221[7:0]) +
	( 14'sd 6284) * $signed(input_fmap_222[7:0]) +
	( 16'sd 29504) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14885) * $signed(input_fmap_224[7:0]) +
	( 16'sd 30172) * $signed(input_fmap_225[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27240) * $signed(input_fmap_227[7:0]) +
	( 15'sd 14071) * $signed(input_fmap_228[7:0]) +
	( 16'sd 16754) * $signed(input_fmap_229[7:0]) +
	( 11'sd 1007) * $signed(input_fmap_230[7:0]) +
	( 15'sd 11276) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7661) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10628) * $signed(input_fmap_233[7:0]) +
	( 15'sd 11441) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22251) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25301) * $signed(input_fmap_236[7:0]) +
	( 13'sd 3610) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27267) * $signed(input_fmap_238[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_239[7:0]) +
	( 15'sd 13471) * $signed(input_fmap_240[7:0]) +
	( 16'sd 16510) * $signed(input_fmap_241[7:0]) +
	( 11'sd 954) * $signed(input_fmap_242[7:0]) +
	( 15'sd 9051) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6050) * $signed(input_fmap_244[7:0]) +
	( 16'sd 17056) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10372) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12025) * $signed(input_fmap_247[7:0]) +
	( 15'sd 11151) * $signed(input_fmap_248[7:0]) +
	( 16'sd 19040) * $signed(input_fmap_249[7:0]) +
	( 11'sd 725) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2756) * $signed(input_fmap_251[7:0]) +
	( 15'sd 9611) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25592) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9814) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24047) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_59;
assign conv_mac_59 = 
	( 15'sd 15980) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7155) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8548) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28354) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15053) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6420) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13975) * $signed(input_fmap_7[7:0]) +
	( 15'sd 8966) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15801) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3808) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6325) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30321) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19264) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19250) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23078) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30856) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1742) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21207) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27451) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4391) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30537) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21761) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12958) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9621) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10138) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20594) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14619) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17823) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16928) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18127) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17723) * $signed(input_fmap_33[7:0]) +
	( 9'sd 246) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8309) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29910) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17364) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13146) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2305) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30823) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17809) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18165) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27935) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27385) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27218) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9622) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9675) * $signed(input_fmap_52[7:0]) +
	( 11'sd 703) * $signed(input_fmap_53[7:0]) +
	( 10'sd 338) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21164) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32407) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13302) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7604) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18621) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11213) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17362) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11606) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25231) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29643) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12778) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28220) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14418) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21494) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1245) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5029) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20356) * $signed(input_fmap_71[7:0]) +
	( 8'sd 98) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27422) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14872) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12204) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3240) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17428) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23917) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16010) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8884) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2421) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27328) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10439) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16842) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21036) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29556) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9602) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22829) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15409) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1229) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14847) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13886) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18428) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24552) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1726) * $signed(input_fmap_101[7:0]) +
	( 11'sd 736) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22131) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3393) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22049) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27697) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9433) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21340) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20630) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26999) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2618) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12601) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5032) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28345) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20759) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14848) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14316) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1837) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21809) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1346) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26925) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26662) * $signed(input_fmap_127[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_128[7:0]) +
	( 16'sd 26273) * $signed(input_fmap_129[7:0]) +
	( 12'sd 2038) * $signed(input_fmap_130[7:0]) +
	( 14'sd 4257) * $signed(input_fmap_131[7:0]) +
	( 16'sd 26445) * $signed(input_fmap_132[7:0]) +
	( 16'sd 20104) * $signed(input_fmap_133[7:0]) +
	( 15'sd 14128) * $signed(input_fmap_134[7:0]) +
	( 10'sd 324) * $signed(input_fmap_135[7:0]) +
	( 14'sd 6005) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26402) * $signed(input_fmap_137[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_138[7:0]) +
	( 14'sd 6128) * $signed(input_fmap_139[7:0]) +
	( 10'sd 339) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3366) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11077) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26103) * $signed(input_fmap_143[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26876) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21992) * $signed(input_fmap_146[7:0]) +
	( 14'sd 7585) * $signed(input_fmap_147[7:0]) +
	( 16'sd 25542) * $signed(input_fmap_148[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_149[7:0]) +
	( 15'sd 13320) * $signed(input_fmap_150[7:0]) +
	( 10'sd 384) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2535) * $signed(input_fmap_152[7:0]) +
	( 15'sd 13480) * $signed(input_fmap_153[7:0]) +
	( 15'sd 16188) * $signed(input_fmap_154[7:0]) +
	( 15'sd 15136) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24711) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25100) * $signed(input_fmap_157[7:0]) +
	( 14'sd 5034) * $signed(input_fmap_158[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_160[7:0]) +
	( 15'sd 12974) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2123) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27486) * $signed(input_fmap_163[7:0]) +
	( 16'sd 20991) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11774) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3517) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7792) * $signed(input_fmap_167[7:0]) +
	( 15'sd 16331) * $signed(input_fmap_168[7:0]) +
	( 15'sd 9472) * $signed(input_fmap_169[7:0]) +
	( 16'sd 32268) * $signed(input_fmap_170[7:0]) +
	( 13'sd 4051) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12640) * $signed(input_fmap_172[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_173[7:0]) +
	( 16'sd 30017) * $signed(input_fmap_174[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_175[7:0]) +
	( 16'sd 31619) * $signed(input_fmap_176[7:0]) +
	( 14'sd 4522) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14954) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25773) * $signed(input_fmap_179[7:0]) +
	( 13'sd 2171) * $signed(input_fmap_180[7:0]) +
	( 12'sd 1734) * $signed(input_fmap_181[7:0]) +
	( 13'sd 3286) * $signed(input_fmap_182[7:0]) +
	( 15'sd 13691) * $signed(input_fmap_183[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5113) * $signed(input_fmap_185[7:0]) +
	( 16'sd 21379) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9110) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13153) * $signed(input_fmap_188[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13976) * $signed(input_fmap_190[7:0]) +
	( 15'sd 16023) * $signed(input_fmap_191[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15974) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3244) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22949) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5649) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26352) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10818) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14822) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15900) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9574) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7726) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25590) * $signed(input_fmap_203[7:0]) +
	( 16'sd 27036) * $signed(input_fmap_204[7:0]) +
	( 16'sd 19840) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9122) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_207[7:0]) +
	( 16'sd 24546) * $signed(input_fmap_208[7:0]) +
	( 16'sd 25971) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19626) * $signed(input_fmap_210[7:0]) +
	( 12'sd 1528) * $signed(input_fmap_211[7:0]) +
	( 15'sd 9174) * $signed(input_fmap_212[7:0]) +
	( 16'sd 21940) * $signed(input_fmap_213[7:0]) +
	( 14'sd 6987) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22251) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28658) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30371) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13884) * $signed(input_fmap_218[7:0]) +
	( 16'sd 31373) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28157) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14374) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15881) * $signed(input_fmap_223[7:0]) +
	( 16'sd 29008) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13437) * $signed(input_fmap_225[7:0]) +
	( 16'sd 28128) * $signed(input_fmap_226[7:0]) +
	( 14'sd 4712) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1293) * $signed(input_fmap_228[7:0]) +
	( 15'sd 11190) * $signed(input_fmap_229[7:0]) +
	( 16'sd 20517) * $signed(input_fmap_230[7:0]) +
	( 15'sd 12103) * $signed(input_fmap_231[7:0]) +
	( 16'sd 23721) * $signed(input_fmap_232[7:0]) +
	( 15'sd 12437) * $signed(input_fmap_233[7:0]) +
	( 16'sd 24078) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5467) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11638) * $signed(input_fmap_237[7:0]) +
	( 15'sd 11276) * $signed(input_fmap_238[7:0]) +
	( 15'sd 14445) * $signed(input_fmap_239[7:0]) +
	( 13'sd 3001) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5135) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28930) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2134) * $signed(input_fmap_243[7:0]) +
	( 16'sd 27428) * $signed(input_fmap_244[7:0]) +
	( 14'sd 4212) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22252) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27842) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4753) * $signed(input_fmap_248[7:0]) +
	( 15'sd 11626) * $signed(input_fmap_249[7:0]) +
	( 16'sd 27815) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_251[7:0]) +
	( 16'sd 19101) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_253[7:0]) +
	( 16'sd 30354) * $signed(input_fmap_254[7:0]) +
	( 16'sd 19305) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_60;
assign conv_mac_60 = 
	( 16'sd 22404) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7168) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2804) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19449) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21678) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10066) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24785) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25781) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18917) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21866) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20277) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7024) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27556) * $signed(input_fmap_12[7:0]) +
	( 11'sd 968) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15538) * $signed(input_fmap_15[7:0]) +
	( 8'sd 98) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22729) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8572) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14170) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2527) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14189) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1379) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32266) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22200) * $signed(input_fmap_25[7:0]) +
	( 11'sd 703) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6738) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29979) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29605) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18006) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24904) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5466) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24246) * $signed(input_fmap_34[7:0]) +
	( 11'sd 811) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32592) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1807) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10024) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17363) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11513) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5643) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7639) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14832) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14083) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25237) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12002) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27001) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31615) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8708) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11978) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30554) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31492) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27320) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29606) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5407) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21422) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18235) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22963) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17521) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7894) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5503) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22400) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15601) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31380) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30642) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13983) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4598) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7791) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13314) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24073) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2136) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13806) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3214) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27501) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21062) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26601) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26183) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7498) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9650) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14762) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23660) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13646) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3832) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12246) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4201) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30917) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5795) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20333) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25018) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11438) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3009) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10014) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18374) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29698) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27016) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2669) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32247) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16197) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27630) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30180) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11171) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13053) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3010) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3639) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5118) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21498) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19342) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29989) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23204) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26301) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4435) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28749) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28940) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3083) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4228) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2260) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10999) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18547) * $signed(input_fmap_130[7:0]) +
	( 13'sd 2879) * $signed(input_fmap_131[7:0]) +
	( 16'sd 31430) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28117) * $signed(input_fmap_133[7:0]) +
	( 16'sd 30890) * $signed(input_fmap_134[7:0]) +
	( 14'sd 8097) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4779) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4956) * $signed(input_fmap_137[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_138[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30373) * $signed(input_fmap_140[7:0]) +
	( 16'sd 28174) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6679) * $signed(input_fmap_142[7:0]) +
	( 16'sd 24819) * $signed(input_fmap_143[7:0]) +
	( 15'sd 8879) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22009) * $signed(input_fmap_145[7:0]) +
	( 16'sd 31571) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30194) * $signed(input_fmap_147[7:0]) +
	( 16'sd 19142) * $signed(input_fmap_148[7:0]) +
	( 15'sd 8538) * $signed(input_fmap_149[7:0]) +
	( 16'sd 30684) * $signed(input_fmap_150[7:0]) +
	( 16'sd 22945) * $signed(input_fmap_151[7:0]) +
	( 15'sd 11176) * $signed(input_fmap_152[7:0]) +
	( 15'sd 15336) * $signed(input_fmap_153[7:0]) +
	( 16'sd 29971) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20756) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25426) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24304) * $signed(input_fmap_157[7:0]) +
	( 15'sd 14632) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_159[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_160[7:0]) +
	( 15'sd 13174) * $signed(input_fmap_161[7:0]) +
	( 16'sd 31651) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8402) * $signed(input_fmap_163[7:0]) +
	( 16'sd 30471) * $signed(input_fmap_164[7:0]) +
	( 15'sd 15366) * $signed(input_fmap_165[7:0]) +
	( 16'sd 23739) * $signed(input_fmap_166[7:0]) +
	( 16'sd 28064) * $signed(input_fmap_167[7:0]) +
	( 16'sd 25757) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30491) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20770) * $signed(input_fmap_170[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_171[7:0]) +
	( 15'sd 8381) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19700) * $signed(input_fmap_173[7:0]) +
	( 15'sd 13117) * $signed(input_fmap_174[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15841) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1806) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22448) * $signed(input_fmap_178[7:0]) +
	( 16'sd 27623) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23257) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15271) * $signed(input_fmap_181[7:0]) +
	( 16'sd 21841) * $signed(input_fmap_182[7:0]) +
	( 15'sd 9428) * $signed(input_fmap_183[7:0]) +
	( 16'sd 23974) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22379) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2697) * $signed(input_fmap_186[7:0]) +
	( 16'sd 21941) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31616) * $signed(input_fmap_188[7:0]) +
	( 16'sd 32498) * $signed(input_fmap_189[7:0]) +
	( 16'sd 18196) * $signed(input_fmap_190[7:0]) +
	( 13'sd 2951) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20564) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9124) * $signed(input_fmap_193[7:0]) +
	( 16'sd 19170) * $signed(input_fmap_194[7:0]) +
	( 15'sd 16341) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15186) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11885) * $signed(input_fmap_197[7:0]) +
	( 14'sd 6594) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6004) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16397) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_202[7:0]) +
	( 16'sd 22583) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2375) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12944) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28102) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7268) * $signed(input_fmap_207[7:0]) +
	( 16'sd 20081) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7734) * $signed(input_fmap_209[7:0]) +
	( 16'sd 32215) * $signed(input_fmap_210[7:0]) +
	( 16'sd 29354) * $signed(input_fmap_211[7:0]) +
	( 14'sd 7844) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5666) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30027) * $signed(input_fmap_214[7:0]) +
	( 15'sd 14677) * $signed(input_fmap_215[7:0]) +
	( 16'sd 27074) * $signed(input_fmap_216[7:0]) +
	( 15'sd 14019) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5613) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3018) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19143) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25765) * $signed(input_fmap_221[7:0]) +
	( 16'sd 24805) * $signed(input_fmap_222[7:0]) +
	( 14'sd 8147) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7924) * $signed(input_fmap_224[7:0]) +
	( 14'sd 4896) * $signed(input_fmap_225[7:0]) +
	( 16'sd 26328) * $signed(input_fmap_226[7:0]) +
	( 16'sd 16956) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26440) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10793) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6505) * $signed(input_fmap_230[7:0]) +
	( 14'sd 5368) * $signed(input_fmap_231[7:0]) +
	( 16'sd 22153) * $signed(input_fmap_232[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13879) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12929) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28764) * $signed(input_fmap_236[7:0]) +
	( 15'sd 12217) * $signed(input_fmap_237[7:0]) +
	( 16'sd 18050) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21975) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31765) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18787) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5075) * $signed(input_fmap_242[7:0]) +
	( 16'sd 30521) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13531) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7360) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14667) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3942) * $signed(input_fmap_247[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_248[7:0]) +
	( 15'sd 8626) * $signed(input_fmap_249[7:0]) +
	( 14'sd 4976) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2259) * $signed(input_fmap_251[7:0]) +
	( 16'sd 23635) * $signed(input_fmap_252[7:0]) +
	( 15'sd 9204) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5248) * $signed(input_fmap_254[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_61;
assign conv_mac_61 = 
	( 15'sd 10469) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3058) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12978) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18050) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25100) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1753) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30675) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7640) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4129) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2420) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16775) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23602) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4791) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26798) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2168) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12920) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20233) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29670) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13791) * $signed(input_fmap_19[7:0]) +
	( 9'sd 254) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11025) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1460) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31550) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21197) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14138) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6249) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32582) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25785) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10159) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13632) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23932) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29160) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8511) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12554) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26471) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1119) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21871) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2554) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25836) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1141) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30653) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8558) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32139) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4973) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1935) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19782) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18215) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22464) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19121) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4119) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21573) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18453) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27535) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1923) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26356) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26682) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30134) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9408) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10355) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15593) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28593) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23020) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3721) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9691) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18915) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26327) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14991) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21166) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2338) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16478) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14206) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22534) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29693) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27264) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32568) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2623) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10726) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2697) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16815) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30391) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16509) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23787) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24129) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16816) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3639) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2713) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8279) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27303) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8515) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8717) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23632) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26908) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4101) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_103[7:0]) +
	( 10'sd 466) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28515) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11853) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15998) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20891) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11069) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19424) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2095) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3046) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26169) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31843) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23111) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9058) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31075) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5700) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21087) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25586) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28423) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22335) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4929) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5542) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5631) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4251) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15630) * $signed(input_fmap_128[7:0]) +
	( 16'sd 29440) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19897) * $signed(input_fmap_130[7:0]) +
	( 16'sd 32726) * $signed(input_fmap_131[7:0]) +
	( 16'sd 17103) * $signed(input_fmap_132[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26908) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13005) * $signed(input_fmap_136[7:0]) +
	( 16'sd 30828) * $signed(input_fmap_137[7:0]) +
	( 15'sd 8522) * $signed(input_fmap_138[7:0]) +
	( 15'sd 16242) * $signed(input_fmap_139[7:0]) +
	( 15'sd 8986) * $signed(input_fmap_140[7:0]) +
	( 16'sd 28858) * $signed(input_fmap_141[7:0]) +
	( 14'sd 5296) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5921) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9421) * $signed(input_fmap_144[7:0]) +
	( 14'sd 8191) * $signed(input_fmap_145[7:0]) +
	( 14'sd 6458) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8194) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17622) * $signed(input_fmap_148[7:0]) +
	( 15'sd 10987) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15675) * $signed(input_fmap_150[7:0]) +
	( 16'sd 16770) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29487) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4561) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25772) * $signed(input_fmap_154[7:0]) +
	( 13'sd 3418) * $signed(input_fmap_155[7:0]) +
	( 14'sd 4113) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22065) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20513) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14679) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17958) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23077) * $signed(input_fmap_161[7:0]) +
	( 9'sd 159) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13667) * $signed(input_fmap_164[7:0]) +
	( 16'sd 26713) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8475) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_167[7:0]) +
	( 16'sd 22756) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21194) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11148) * $signed(input_fmap_170[7:0]) +
	( 15'sd 13096) * $signed(input_fmap_171[7:0]) +
	( 16'sd 20547) * $signed(input_fmap_172[7:0]) +
	( 14'sd 7498) * $signed(input_fmap_173[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_174[7:0]) +
	( 15'sd 13471) * $signed(input_fmap_175[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_176[7:0]) +
	( 16'sd 21186) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17176) * $signed(input_fmap_178[7:0]) +
	( 16'sd 24714) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15260) * $signed(input_fmap_180[7:0]) +
	( 16'sd 20040) * $signed(input_fmap_181[7:0]) +
	( 15'sd 9218) * $signed(input_fmap_182[7:0]) +
	( 16'sd 23712) * $signed(input_fmap_183[7:0]) +
	( 16'sd 19210) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11803) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23672) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5896) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12264) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_189[7:0]) +
	( 11'sd 863) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29952) * $signed(input_fmap_191[7:0]) +
	( 14'sd 7962) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15421) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21714) * $signed(input_fmap_194[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_195[7:0]) +
	( 15'sd 9452) * $signed(input_fmap_196[7:0]) +
	( 16'sd 23557) * $signed(input_fmap_197[7:0]) +
	( 15'sd 16278) * $signed(input_fmap_198[7:0]) +
	( 16'sd 19724) * $signed(input_fmap_199[7:0]) +
	( 16'sd 21893) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11045) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8813) * $signed(input_fmap_202[7:0]) +
	( 16'sd 31599) * $signed(input_fmap_203[7:0]) +
	( 10'sd 509) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24860) * $signed(input_fmap_205[7:0]) +
	( 14'sd 5801) * $signed(input_fmap_206[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_207[7:0]) +
	( 16'sd 27943) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23660) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18744) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12581) * $signed(input_fmap_211[7:0]) +
	( 11'sd 880) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9942) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1206) * $signed(input_fmap_214[7:0]) +
	( 16'sd 16523) * $signed(input_fmap_215[7:0]) +
	( 16'sd 30874) * $signed(input_fmap_216[7:0]) +
	( 15'sd 8237) * $signed(input_fmap_217[7:0]) +
	( 16'sd 27707) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10739) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19770) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19921) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14368) * $signed(input_fmap_222[7:0]) +
	( 16'sd 21041) * $signed(input_fmap_223[7:0]) +
	( 16'sd 24531) * $signed(input_fmap_224[7:0]) +
	( 14'sd 7138) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30685) * $signed(input_fmap_226[7:0]) +
	( 10'sd 310) * $signed(input_fmap_227[7:0]) +
	( 11'sd 823) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23151) * $signed(input_fmap_229[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_230[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9784) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21780) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_234[7:0]) +
	( 16'sd 27119) * $signed(input_fmap_235[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_236[7:0]) +
	( 16'sd 30703) * $signed(input_fmap_237[7:0]) +
	( 16'sd 32454) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13412) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18146) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30115) * $signed(input_fmap_241[7:0]) +
	( 13'sd 2547) * $signed(input_fmap_242[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22382) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19388) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1881) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11206) * $signed(input_fmap_247[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25388) * $signed(input_fmap_249[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_250[7:0]) +
	( 16'sd 31813) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30401) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28105) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19528) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_62;
assign conv_mac_62 = 
	( 16'sd 23133) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23361) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20827) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7737) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30728) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5135) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15874) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27897) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31259) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29949) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3947) * $signed(input_fmap_11[7:0]) +
	( 16'sd 16424) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14102) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14345) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31977) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2858) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11046) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11194) * $signed(input_fmap_19[7:0]) +
	( 10'sd 376) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22531) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18767) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9362) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27401) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11031) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30687) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6215) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18303) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11769) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4722) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_35[7:0]) +
	( 11'sd 648) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16483) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14133) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6265) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16191) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1860) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24176) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13687) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26581) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26481) * $signed(input_fmap_46[7:0]) +
	( 11'sd 570) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8730) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25868) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22017) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1850) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19642) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32695) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15978) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26664) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31675) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22465) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22224) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8457) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21823) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3571) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32304) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28051) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21878) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5087) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26406) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23069) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15316) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30582) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10500) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27492) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15389) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23069) * $signed(input_fmap_78[7:0]) +
	( 11'sd 575) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22959) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10454) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10575) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18571) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7734) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23283) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11865) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15831) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27237) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30498) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18773) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15469) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24361) * $signed(input_fmap_93[7:0]) +
	( 12'sd 2014) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28985) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28696) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22403) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5939) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32728) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25879) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10331) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27751) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17282) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5899) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21681) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9061) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7066) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12187) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1173) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30655) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19215) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1296) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30409) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12535) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2650) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2979) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24892) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30266) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7224) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6454) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16485) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11398) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2354) * $signed(input_fmap_127[7:0]) +
	( 16'sd 21903) * $signed(input_fmap_128[7:0]) +
	( 10'sd 386) * $signed(input_fmap_129[7:0]) +
	( 14'sd 5511) * $signed(input_fmap_130[7:0]) +
	( 11'sd 597) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1596) * $signed(input_fmap_132[7:0]) +
	( 12'sd 1642) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18968) * $signed(input_fmap_134[7:0]) +
	( 16'sd 22631) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23430) * $signed(input_fmap_136[7:0]) +
	( 16'sd 29215) * $signed(input_fmap_137[7:0]) +
	( 16'sd 25129) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18861) * $signed(input_fmap_139[7:0]) +
	( 16'sd 23118) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5149) * $signed(input_fmap_141[7:0]) +
	( 16'sd 32578) * $signed(input_fmap_142[7:0]) +
	( 15'sd 8766) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4430) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_146[7:0]) +
	( 16'sd 25680) * $signed(input_fmap_147[7:0]) +
	( 15'sd 9873) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_149[7:0]) +
	( 14'sd 7522) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_151[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11315) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10245) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12262) * $signed(input_fmap_155[7:0]) +
	( 15'sd 11270) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13554) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25576) * $signed(input_fmap_158[7:0]) +
	( 15'sd 10846) * $signed(input_fmap_159[7:0]) +
	( 14'sd 4744) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19313) * $signed(input_fmap_161[7:0]) +
	( 15'sd 12993) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2117) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9940) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14604) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31900) * $signed(input_fmap_166[7:0]) +
	( 15'sd 15449) * $signed(input_fmap_167[7:0]) +
	( 16'sd 25988) * $signed(input_fmap_168[7:0]) +
	( 16'sd 24402) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5729) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30951) * $signed(input_fmap_171[7:0]) +
	( 16'sd 30053) * $signed(input_fmap_172[7:0]) +
	( 12'sd 2003) * $signed(input_fmap_173[7:0]) +
	( 11'sd 712) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25392) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_177[7:0]) +
	( 15'sd 13239) * $signed(input_fmap_178[7:0]) +
	( 15'sd 8887) * $signed(input_fmap_179[7:0]) +
	( 16'sd 31458) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28670) * $signed(input_fmap_181[7:0]) +
	( 16'sd 24890) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25674) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8748) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11604) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2386) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11405) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29077) * $signed(input_fmap_188[7:0]) +
	( 15'sd 12232) * $signed(input_fmap_189[7:0]) +
	( 10'sd 399) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31045) * $signed(input_fmap_191[7:0]) +
	( 15'sd 13079) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5150) * $signed(input_fmap_193[7:0]) +
	( 16'sd 31852) * $signed(input_fmap_194[7:0]) +
	( 16'sd 21200) * $signed(input_fmap_195[7:0]) +
	( 16'sd 23987) * $signed(input_fmap_196[7:0]) +
	( 16'sd 17617) * $signed(input_fmap_197[7:0]) +
	( 15'sd 12906) * $signed(input_fmap_198[7:0]) +
	( 16'sd 17892) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13736) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15267) * $signed(input_fmap_201[7:0]) +
	( 15'sd 15348) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19481) * $signed(input_fmap_203[7:0]) +
	( 13'sd 3247) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30071) * $signed(input_fmap_205[7:0]) +
	( 16'sd 22046) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5389) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4414) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19138) * $signed(input_fmap_209[7:0]) +
	( 15'sd 8220) * $signed(input_fmap_210[7:0]) +
	( 16'sd 18150) * $signed(input_fmap_211[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_212[7:0]) +
	( 16'sd 22168) * $signed(input_fmap_213[7:0]) +
	( 16'sd 22039) * $signed(input_fmap_214[7:0]) +
	( 15'sd 13539) * $signed(input_fmap_215[7:0]) +
	( 15'sd 9870) * $signed(input_fmap_216[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_217[7:0]) +
	( 15'sd 14705) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20569) * $signed(input_fmap_219[7:0]) +
	( 15'sd 11533) * $signed(input_fmap_220[7:0]) +
	( 13'sd 2339) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12897) * $signed(input_fmap_222[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12752) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2217) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11908) * $signed(input_fmap_226[7:0]) +
	( 16'sd 28891) * $signed(input_fmap_227[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26087) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30629) * $signed(input_fmap_230[7:0]) +
	( 14'sd 4891) * $signed(input_fmap_231[7:0]) +
	( 16'sd 28968) * $signed(input_fmap_232[7:0]) +
	( 14'sd 7786) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_234[7:0]) +
	( 16'sd 18986) * $signed(input_fmap_235[7:0]) +
	( 14'sd 6206) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6715) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22452) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31303) * $signed(input_fmap_239[7:0]) +
	( 14'sd 5610) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15071) * $signed(input_fmap_241[7:0]) +
	( 15'sd 13704) * $signed(input_fmap_242[7:0]) +
	( 11'sd 687) * $signed(input_fmap_243[7:0]) +
	( 15'sd 10247) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2651) * $signed(input_fmap_245[7:0]) +
	( 16'sd 26509) * $signed(input_fmap_246[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_247[7:0]) +
	( 16'sd 19534) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12721) * $signed(input_fmap_249[7:0]) +
	( 14'sd 8095) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15572) * $signed(input_fmap_251[7:0]) +
	( 16'sd 29177) * $signed(input_fmap_252[7:0]) +
	( 16'sd 23856) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5753) * $signed(input_fmap_254[7:0]) +
	( 16'sd 31003) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_63;
assign conv_mac_63 = 
	( 16'sd 31510) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13497) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3939) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10078) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23054) * $signed(input_fmap_8[7:0]) +
	( 10'sd 390) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10155) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31786) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29102) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9964) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22858) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28538) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23328) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1907) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14646) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2384) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13319) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10751) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3050) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10796) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7831) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22421) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5751) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16990) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16405) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4959) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5005) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13555) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3853) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15805) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8327) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26681) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26725) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23144) * $signed(input_fmap_42[7:0]) +
	( 11'sd 681) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2704) * $signed(input_fmap_44[7:0]) +
	( 8'sd 94) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15852) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30354) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26117) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18690) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19404) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27094) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7262) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8278) * $signed(input_fmap_56[7:0]) +
	( 11'sd 1023) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14330) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22368) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3298) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7571) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3121) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1208) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1082) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24486) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27002) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3138) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25042) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16130) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18300) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21637) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27415) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21644) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27736) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27111) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22421) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5464) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5745) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31257) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23860) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24482) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13438) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25483) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5119) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25178) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19613) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30304) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18525) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18905) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17168) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24123) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21239) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28385) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3962) * $signed(input_fmap_97[7:0]) +
	( 11'sd 543) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25529) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7419) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14120) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13974) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32740) * $signed(input_fmap_104[7:0]) +
	( 15'sd 16213) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9392) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12302) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12772) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4886) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9716) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17800) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26819) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22953) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25598) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6403) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4717) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21330) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32470) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8930) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32565) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13139) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29013) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11132) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28317) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13590) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29151) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5708) * $signed(input_fmap_129[7:0]) +
	( 13'sd 2784) * $signed(input_fmap_130[7:0]) +
	( 14'sd 4124) * $signed(input_fmap_131[7:0]) +
	( 16'sd 16837) * $signed(input_fmap_132[7:0]) +
	( 11'sd 749) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4952) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20139) * $signed(input_fmap_135[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_136[7:0]) +
	( 16'sd 23212) * $signed(input_fmap_137[7:0]) +
	( 15'sd 13305) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3802) * $signed(input_fmap_139[7:0]) +
	( 11'sd 572) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5138) * $signed(input_fmap_141[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_142[7:0]) +
	( 14'sd 6073) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28580) * $signed(input_fmap_144[7:0]) +
	( 14'sd 5215) * $signed(input_fmap_145[7:0]) +
	( 16'sd 30802) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18687) * $signed(input_fmap_147[7:0]) +
	( 16'sd 18709) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17996) * $signed(input_fmap_149[7:0]) +
	( 12'sd 1111) * $signed(input_fmap_150[7:0]) +
	( 16'sd 29612) * $signed(input_fmap_151[7:0]) +
	( 16'sd 26961) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1863) * $signed(input_fmap_153[7:0]) +
	( 16'sd 17143) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19287) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28599) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27396) * $signed(input_fmap_157[7:0]) +
	( 15'sd 13912) * $signed(input_fmap_158[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24171) * $signed(input_fmap_160[7:0]) +
	( 16'sd 17020) * $signed(input_fmap_161[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_162[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13674) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23237) * $signed(input_fmap_165[7:0]) +
	( 15'sd 15781) * $signed(input_fmap_166[7:0]) +
	( 16'sd 27779) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26508) * $signed(input_fmap_168[7:0]) +
	( 16'sd 19534) * $signed(input_fmap_169[7:0]) +
	( 15'sd 16107) * $signed(input_fmap_170[7:0]) +
	( 11'sd 651) * $signed(input_fmap_171[7:0]) +
	( 12'sd 2001) * $signed(input_fmap_172[7:0]) +
	( 10'sd 482) * $signed(input_fmap_173[7:0]) +
	( 16'sd 24555) * $signed(input_fmap_174[7:0]) +
	( 15'sd 8243) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15652) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22844) * $signed(input_fmap_177[7:0]) +
	( 15'sd 11540) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2256) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28479) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15768) * $signed(input_fmap_181[7:0]) +
	( 16'sd 25403) * $signed(input_fmap_182[7:0]) +
	( 14'sd 6838) * $signed(input_fmap_183[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26915) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4137) * $signed(input_fmap_186[7:0]) +
	( 16'sd 17836) * $signed(input_fmap_187[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_188[7:0]) +
	( 12'sd 1770) * $signed(input_fmap_189[7:0]) +
	( 16'sd 24974) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19667) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31684) * $signed(input_fmap_192[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_193[7:0]) +
	( 15'sd 15158) * $signed(input_fmap_194[7:0]) +
	( 15'sd 15102) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15013) * $signed(input_fmap_196[7:0]) +
	( 13'sd 3707) * $signed(input_fmap_197[7:0]) +
	( 16'sd 25762) * $signed(input_fmap_198[7:0]) +
	( 15'sd 13641) * $signed(input_fmap_199[7:0]) +
	( 14'sd 4697) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12769) * $signed(input_fmap_201[7:0]) +
	( 16'sd 25380) * $signed(input_fmap_202[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_203[7:0]) +
	( 15'sd 10386) * $signed(input_fmap_204[7:0]) +
	( 16'sd 23559) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3995) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5013) * $signed(input_fmap_207[7:0]) +
	( 16'sd 27518) * $signed(input_fmap_208[7:0]) +
	( 10'sd 511) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10488) * $signed(input_fmap_210[7:0]) +
	( 15'sd 11436) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12778) * $signed(input_fmap_213[7:0]) +
	( 16'sd 27608) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9280) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4381) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25518) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5280) * $signed(input_fmap_218[7:0]) +
	( 16'sd 27308) * $signed(input_fmap_219[7:0]) +
	( 14'sd 6560) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13873) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2519) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22710) * $signed(input_fmap_223[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32361) * $signed(input_fmap_226[7:0]) +
	( 16'sd 29441) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4457) * $signed(input_fmap_228[7:0]) +
	( 14'sd 5232) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7201) * $signed(input_fmap_230[7:0]) +
	( 11'sd 697) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15680) * $signed(input_fmap_232[7:0]) +
	( 16'sd 25531) * $signed(input_fmap_233[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_234[7:0]) +
	( 16'sd 17491) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10058) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19386) * $signed(input_fmap_237[7:0]) +
	( 12'sd 1972) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22099) * $signed(input_fmap_239[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_240[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_241[7:0]) +
	( 16'sd 25234) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25438) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18871) * $signed(input_fmap_244[7:0]) +
	( 16'sd 27298) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31858) * $signed(input_fmap_246[7:0]) +
	( 16'sd 29070) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1542) * $signed(input_fmap_248[7:0]) +
	( 16'sd 31482) * $signed(input_fmap_249[7:0]) +
	( 14'sd 8000) * $signed(input_fmap_250[7:0]) +
	( 16'sd 16899) * $signed(input_fmap_251[7:0]) +
	( 8'sd 100) * $signed(input_fmap_252[7:0]) +
	( 16'sd 23534) * $signed(input_fmap_253[7:0]) +
	( 15'sd 11375) * $signed(input_fmap_254[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_64;
assign conv_mac_64 = 
	( 15'sd 12355) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16810) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_2[7:0]) +
	( 15'sd 16112) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19574) * $signed(input_fmap_4[7:0]) +
	( 11'sd 986) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2894) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13756) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22063) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5581) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24270) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17249) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19135) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14314) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6354) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32594) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28579) * $signed(input_fmap_20[7:0]) +
	( 10'sd 265) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21082) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4457) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18026) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7260) * $signed(input_fmap_27[7:0]) +
	( 8'sd 76) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2524) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28280) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1027) * $signed(input_fmap_33[7:0]) +
	( 11'sd 952) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8242) * $signed(input_fmap_35[7:0]) +
	( 11'sd 780) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25749) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14483) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23546) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21655) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2182) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22831) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1920) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3364) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32588) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26831) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20481) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23493) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15824) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20378) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26962) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27198) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22204) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1602) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30208) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3357) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31681) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29956) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15938) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11418) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19831) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16982) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25820) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4139) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28574) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2719) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15607) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_70[7:0]) +
	( 11'sd 842) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26595) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30688) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7974) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12401) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5728) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24240) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16024) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28492) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1744) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19325) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14766) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25763) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26202) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20626) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20406) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12805) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20458) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14488) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17970) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11353) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19570) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32471) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19175) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15917) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28813) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3327) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1210) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17795) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7958) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11050) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19543) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12144) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21220) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10953) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28706) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8658) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11994) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20452) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25471) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24319) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1793) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26704) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11400) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7937) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23379) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16855) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20856) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19504) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24971) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10875) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31922) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27418) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30572) * $signed(input_fmap_130[7:0]) +
	( 16'sd 25652) * $signed(input_fmap_131[7:0]) +
	( 14'sd 6171) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31200) * $signed(input_fmap_133[7:0]) +
	( 16'sd 20312) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21450) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_136[7:0]) +
	( 16'sd 28983) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27908) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31719) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3710) * $signed(input_fmap_140[7:0]) +
	( 15'sd 15697) * $signed(input_fmap_141[7:0]) +
	( 13'sd 3518) * $signed(input_fmap_142[7:0]) +
	( 14'sd 6623) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4505) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7657) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9693) * $signed(input_fmap_146[7:0]) +
	( 14'sd 6984) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4599) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2188) * $signed(input_fmap_149[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_150[7:0]) +
	( 14'sd 7361) * $signed(input_fmap_151[7:0]) +
	( 16'sd 26786) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11398) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20391) * $signed(input_fmap_156[7:0]) +
	( 16'sd 32025) * $signed(input_fmap_157[7:0]) +
	( 16'sd 32660) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32014) * $signed(input_fmap_159[7:0]) +
	( 16'sd 32272) * $signed(input_fmap_160[7:0]) +
	( 16'sd 21646) * $signed(input_fmap_161[7:0]) +
	( 14'sd 6595) * $signed(input_fmap_162[7:0]) +
	( 16'sd 23984) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11327) * $signed(input_fmap_164[7:0]) +
	( 16'sd 32504) * $signed(input_fmap_165[7:0]) +
	( 14'sd 5313) * $signed(input_fmap_166[7:0]) +
	( 16'sd 22887) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9155) * $signed(input_fmap_168[7:0]) +
	( 14'sd 4839) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5302) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24338) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4632) * $signed(input_fmap_172[7:0]) +
	( 15'sd 10981) * $signed(input_fmap_173[7:0]) +
	( 15'sd 12271) * $signed(input_fmap_174[7:0]) +
	( 15'sd 10117) * $signed(input_fmap_175[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_176[7:0]) +
	( 15'sd 8205) * $signed(input_fmap_177[7:0]) +
	( 16'sd 18908) * $signed(input_fmap_178[7:0]) +
	( 16'sd 17632) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6281) * $signed(input_fmap_180[7:0]) +
	( 15'sd 10813) * $signed(input_fmap_181[7:0]) +
	( 13'sd 3034) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_183[7:0]) +
	( 13'sd 3363) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22815) * $signed(input_fmap_185[7:0]) +
	( 15'sd 10304) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27368) * $signed(input_fmap_187[7:0]) +
	( 16'sd 20705) * $signed(input_fmap_188[7:0]) +
	( 15'sd 8744) * $signed(input_fmap_189[7:0]) +
	( 16'sd 25135) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26014) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29017) * $signed(input_fmap_192[7:0]) +
	( 16'sd 16901) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21562) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17694) * $signed(input_fmap_195[7:0]) +
	( 13'sd 2084) * $signed(input_fmap_196[7:0]) +
	( 16'sd 29277) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18797) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24181) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25277) * $signed(input_fmap_200[7:0]) +
	( 16'sd 24779) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8224) * $signed(input_fmap_202[7:0]) +
	( 8'sd 96) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5328) * $signed(input_fmap_204[7:0]) +
	( 16'sd 26735) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2372) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28600) * $signed(input_fmap_207[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_208[7:0]) +
	( 16'sd 28852) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19726) * $signed(input_fmap_210[7:0]) +
	( 12'sd 1372) * $signed(input_fmap_211[7:0]) +
	( 7'sd 44) * $signed(input_fmap_212[7:0]) +
	( 16'sd 16730) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15066) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23232) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4608) * $signed(input_fmap_216[7:0]) +
	( 11'sd 657) * $signed(input_fmap_217[7:0]) +
	( 16'sd 17595) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10101) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22713) * $signed(input_fmap_220[7:0]) +
	( 15'sd 9306) * $signed(input_fmap_221[7:0]) +
	( 14'sd 6618) * $signed(input_fmap_222[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_223[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_224[7:0]) +
	( 15'sd 11611) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32113) * $signed(input_fmap_226[7:0]) +
	( 12'sd 1876) * $signed(input_fmap_227[7:0]) +
	( 14'sd 8135) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20435) * $signed(input_fmap_229[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_230[7:0]) +
	( 16'sd 26731) * $signed(input_fmap_231[7:0]) +
	( 16'sd 28456) * $signed(input_fmap_232[7:0]) +
	( 16'sd 19359) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14899) * $signed(input_fmap_234[7:0]) +
	( 11'sd 941) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2717) * $signed(input_fmap_237[7:0]) +
	( 16'sd 32743) * $signed(input_fmap_238[7:0]) +
	( 13'sd 3938) * $signed(input_fmap_239[7:0]) +
	( 16'sd 28825) * $signed(input_fmap_240[7:0]) +
	( 16'sd 16490) * $signed(input_fmap_241[7:0]) +
	( 15'sd 10977) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2417) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2638) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3557) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28972) * $signed(input_fmap_246[7:0]) +
	( 16'sd 29197) * $signed(input_fmap_247[7:0]) +
	( 15'sd 14441) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_249[7:0]) +
	( 16'sd 29115) * $signed(input_fmap_250[7:0]) +
	( 15'sd 10912) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2361) * $signed(input_fmap_252[7:0]) +
	( 9'sd 218) * $signed(input_fmap_253[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_254[7:0]) +
	( 10'sd 328) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_65;
assign conv_mac_65 = 
	( 14'sd 6014) * $signed(input_fmap_0[7:0]) +
	( 11'sd 741) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29625) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23894) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5184) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9478) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31028) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28752) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12528) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20986) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14290) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20891) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10377) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19456) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18500) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17737) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14689) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9462) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3848) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1984) * $signed(input_fmap_20[7:0]) +
	( 16'sd 29830) * $signed(input_fmap_21[7:0]) +
	( 10'sd 300) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8833) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20197) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31295) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7237) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27080) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25770) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2748) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31750) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18922) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29179) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20710) * $signed(input_fmap_34[7:0]) +
	( 13'sd 4064) * $signed(input_fmap_35[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17887) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14332) * $signed(input_fmap_38[7:0]) +
	( 14'sd 8112) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27357) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17217) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10646) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5245) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4785) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29569) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16812) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5795) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11302) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28876) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27900) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18972) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28320) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3047) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24077) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13103) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15987) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12984) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7010) * $signed(input_fmap_62[7:0]) +
	( 11'sd 582) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2838) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32728) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31987) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21755) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6586) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24980) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20326) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17714) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29301) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28315) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11074) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31676) * $signed(input_fmap_75[7:0]) +
	( 11'sd 768) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3272) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17457) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17978) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13821) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11835) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11250) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3057) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7592) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2314) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16880) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16200) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14128) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5767) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31065) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3303) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11503) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18692) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13762) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30233) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23615) * $signed(input_fmap_101[7:0]) +
	( 9'sd 232) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10393) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12260) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32139) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21053) * $signed(input_fmap_106[7:0]) +
	( 11'sd 842) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5114) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28044) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20449) * $signed(input_fmap_110[7:0]) +
	( 11'sd 822) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5627) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1797) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22096) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17003) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2784) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9067) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24455) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27916) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10205) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23981) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21461) * $signed(input_fmap_122[7:0]) +
	( 13'sd 4013) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27981) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29984) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27059) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19352) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4772) * $signed(input_fmap_128[7:0]) +
	( 15'sd 8664) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19662) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23154) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10818) * $signed(input_fmap_132[7:0]) +
	( 16'sd 30781) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1132) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23224) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8919) * $signed(input_fmap_136[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32377) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20349) * $signed(input_fmap_139[7:0]) +
	( 11'sd 868) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20943) * $signed(input_fmap_141[7:0]) +
	( 16'sd 18918) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5050) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17719) * $signed(input_fmap_145[7:0]) +
	( 15'sd 10152) * $signed(input_fmap_146[7:0]) +
	( 15'sd 16243) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26314) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2885) * $signed(input_fmap_149[7:0]) +
	( 11'sd 1006) * $signed(input_fmap_150[7:0]) +
	( 16'sd 32389) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23985) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14578) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25825) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10178) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18995) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31577) * $signed(input_fmap_157[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12721) * $signed(input_fmap_159[7:0]) +
	( 16'sd 25101) * $signed(input_fmap_160[7:0]) +
	( 16'sd 18157) * $signed(input_fmap_161[7:0]) +
	( 15'sd 8603) * $signed(input_fmap_162[7:0]) +
	( 15'sd 11878) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1565) * $signed(input_fmap_164[7:0]) +
	( 16'sd 16583) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9214) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13377) * $signed(input_fmap_167[7:0]) +
	( 16'sd 27737) * $signed(input_fmap_168[7:0]) +
	( 15'sd 9313) * $signed(input_fmap_169[7:0]) +
	( 16'sd 26205) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15242) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22112) * $signed(input_fmap_172[7:0]) +
	( 15'sd 14970) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10944) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1120) * $signed(input_fmap_175[7:0]) +
	( 16'sd 25318) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_177[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_178[7:0]) +
	( 16'sd 16741) * $signed(input_fmap_179[7:0]) +
	( 16'sd 30664) * $signed(input_fmap_180[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_181[7:0]) +
	( 16'sd 18726) * $signed(input_fmap_182[7:0]) +
	( 15'sd 11992) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13428) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25238) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4558) * $signed(input_fmap_186[7:0]) +
	( 16'sd 29715) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21905) * $signed(input_fmap_188[7:0]) +
	( 15'sd 16047) * $signed(input_fmap_189[7:0]) +
	( 16'sd 26469) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19261) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28365) * $signed(input_fmap_192[7:0]) +
	( 16'sd 25321) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9175) * $signed(input_fmap_194[7:0]) +
	( 14'sd 7419) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24807) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32507) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29154) * $signed(input_fmap_198[7:0]) +
	( 13'sd 2359) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6455) * $signed(input_fmap_200[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_201[7:0]) +
	( 16'sd 23356) * $signed(input_fmap_202[7:0]) +
	( 16'sd 17257) * $signed(input_fmap_203[7:0]) +
	( 16'sd 29237) * $signed(input_fmap_204[7:0]) +
	( 16'sd 25216) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_206[7:0]) +
	( 15'sd 8630) * $signed(input_fmap_207[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_208[7:0]) +
	( 16'sd 28382) * $signed(input_fmap_209[7:0]) +
	( 16'sd 25480) * $signed(input_fmap_210[7:0]) +
	( 16'sd 21445) * $signed(input_fmap_211[7:0]) +
	( 16'sd 28742) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23940) * $signed(input_fmap_213[7:0]) +
	( 15'sd 16210) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11868) * $signed(input_fmap_215[7:0]) +
	( 15'sd 13076) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24508) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5800) * $signed(input_fmap_218[7:0]) +
	( 15'sd 9669) * $signed(input_fmap_219[7:0]) +
	( 16'sd 27669) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12082) * $signed(input_fmap_221[7:0]) +
	( 11'sd 830) * $signed(input_fmap_222[7:0]) +
	( 14'sd 5350) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6836) * $signed(input_fmap_224[7:0]) +
	( 16'sd 22345) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6006) * $signed(input_fmap_226[7:0]) +
	( 15'sd 11430) * $signed(input_fmap_227[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_228[7:0]) +
	( 16'sd 28609) * $signed(input_fmap_229[7:0]) +
	( 16'sd 24611) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18309) * $signed(input_fmap_231[7:0]) +
	( 14'sd 5864) * $signed(input_fmap_232[7:0]) +
	( 14'sd 7017) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3850) * $signed(input_fmap_234[7:0]) +
	( 15'sd 9190) * $signed(input_fmap_235[7:0]) +
	( 16'sd 32003) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10979) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17498) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22591) * $signed(input_fmap_239[7:0]) +
	( 15'sd 13879) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3067) * $signed(input_fmap_241[7:0]) +
	( 15'sd 12842) * $signed(input_fmap_242[7:0]) +
	( 15'sd 15505) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24353) * $signed(input_fmap_244[7:0]) +
	( 9'sd 161) * $signed(input_fmap_245[7:0]) +
	( 16'sd 27070) * $signed(input_fmap_246[7:0]) +
	( 15'sd 16014) * $signed(input_fmap_247[7:0]) +
	( 10'sd 467) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25500) * $signed(input_fmap_249[7:0]) +
	( 16'sd 19075) * $signed(input_fmap_250[7:0]) +
	( 16'sd 17800) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26117) * $signed(input_fmap_252[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_253[7:0]) +
	( 11'sd 678) * $signed(input_fmap_254[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_66;
assign conv_mac_66 = 
	( 15'sd 11257) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30042) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22209) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29118) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3548) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30273) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2861) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25899) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16832) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7829) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1503) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24726) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13079) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19659) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28212) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7667) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6796) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26359) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27994) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20195) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27920) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1673) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15167) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5021) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31794) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9103) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20767) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8298) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22627) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23245) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30457) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8872) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1347) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29725) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11969) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9417) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1455) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30784) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2290) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10260) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7695) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29441) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15228) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31560) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17949) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21753) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32201) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6554) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28227) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16891) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4905) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23149) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31268) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21919) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23221) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3961) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20163) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4209) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27644) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25514) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27890) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11678) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8445) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27555) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18381) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7646) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17858) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27775) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23279) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27173) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26591) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22043) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15263) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24244) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12649) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32512) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22179) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6993) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12996) * $signed(input_fmap_93[7:0]) +
	( 11'sd 1000) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16371) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29285) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24817) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10157) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13431) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14226) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17868) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17967) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31970) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17221) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32752) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13689) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32316) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_109[7:0]) +
	( 10'sd 435) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32576) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20365) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13709) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7767) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11776) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21998) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21597) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10963) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18246) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4930) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19575) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16540) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7761) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29921) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25824) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15246) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30429) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14316) * $signed(input_fmap_129[7:0]) +
	( 14'sd 7163) * $signed(input_fmap_130[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_131[7:0]) +
	( 13'sd 2247) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22464) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1795) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18355) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8591) * $signed(input_fmap_136[7:0]) +
	( 16'sd 20108) * $signed(input_fmap_137[7:0]) +
	( 14'sd 4736) * $signed(input_fmap_138[7:0]) +
	( 9'sd 252) * $signed(input_fmap_139[7:0]) +
	( 10'sd 338) * $signed(input_fmap_140[7:0]) +
	( 16'sd 32767) * $signed(input_fmap_141[7:0]) +
	( 16'sd 18482) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5513) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18900) * $signed(input_fmap_144[7:0]) +
	( 16'sd 32267) * $signed(input_fmap_145[7:0]) +
	( 15'sd 8728) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19378) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4912) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7813) * $signed(input_fmap_149[7:0]) +
	( 16'sd 29997) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30852) * $signed(input_fmap_151[7:0]) +
	( 16'sd 19705) * $signed(input_fmap_152[7:0]) +
	( 14'sd 6422) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30482) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19955) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20190) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11612) * $signed(input_fmap_158[7:0]) +
	( 16'sd 28661) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17677) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28181) * $signed(input_fmap_161[7:0]) +
	( 16'sd 18657) * $signed(input_fmap_162[7:0]) +
	( 15'sd 10298) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3244) * $signed(input_fmap_164[7:0]) +
	( 14'sd 5035) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12194) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20737) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5462) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6629) * $signed(input_fmap_169[7:0]) +
	( 13'sd 3448) * $signed(input_fmap_170[7:0]) +
	( 16'sd 27134) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22678) * $signed(input_fmap_172[7:0]) +
	( 15'sd 10671) * $signed(input_fmap_173[7:0]) +
	( 11'sd 887) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7607) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18230) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27807) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25348) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_180[7:0]) +
	( 12'sd 1576) * $signed(input_fmap_181[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_182[7:0]) +
	( 16'sd 19664) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8691) * $signed(input_fmap_184[7:0]) +
	( 15'sd 10331) * $signed(input_fmap_185[7:0]) +
	( 16'sd 27642) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11719) * $signed(input_fmap_187[7:0]) +
	( 10'sd 331) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25074) * $signed(input_fmap_189[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_190[7:0]) +
	( 11'sd 700) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19284) * $signed(input_fmap_192[7:0]) +
	( 12'sd 1105) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12287) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14238) * $signed(input_fmap_195[7:0]) +
	( 16'sd 29821) * $signed(input_fmap_196[7:0]) +
	( 13'sd 3989) * $signed(input_fmap_197[7:0]) +
	( 15'sd 15550) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10287) * $signed(input_fmap_199[7:0]) +
	( 15'sd 11325) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3160) * $signed(input_fmap_201[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_202[7:0]) +
	( 14'sd 7937) * $signed(input_fmap_203[7:0]) +
	( 16'sd 24882) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6053) * $signed(input_fmap_205[7:0]) +
	( 16'sd 16442) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3624) * $signed(input_fmap_207[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_208[7:0]) +
	( 13'sd 2818) * $signed(input_fmap_209[7:0]) +
	( 13'sd 2319) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26160) * $signed(input_fmap_211[7:0]) +
	( 16'sd 23829) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28676) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15958) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6708) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19997) * $signed(input_fmap_216[7:0]) +
	( 16'sd 21684) * $signed(input_fmap_217[7:0]) +
	( 16'sd 18132) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20943) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_220[7:0]) +
	( 14'sd 7458) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28251) * $signed(input_fmap_222[7:0]) +
	( 16'sd 16537) * $signed(input_fmap_223[7:0]) +
	( 16'sd 24570) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20152) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30261) * $signed(input_fmap_226[7:0]) +
	( 16'sd 29998) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19124) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10154) * $signed(input_fmap_229[7:0]) +
	( 11'sd 689) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_231[7:0]) +
	( 16'sd 23228) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23444) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14136) * $signed(input_fmap_234[7:0]) +
	( 14'sd 4512) * $signed(input_fmap_235[7:0]) +
	( 16'sd 18693) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11821) * $signed(input_fmap_237[7:0]) +
	( 16'sd 29846) * $signed(input_fmap_238[7:0]) +
	( 15'sd 10005) * $signed(input_fmap_239[7:0]) +
	( 14'sd 4688) * $signed(input_fmap_240[7:0]) +
	( 15'sd 16333) * $signed(input_fmap_241[7:0]) +
	( 14'sd 7898) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10478) * $signed(input_fmap_243[7:0]) +
	( 15'sd 16237) * $signed(input_fmap_244[7:0]) +
	( 11'sd 516) * $signed(input_fmap_245[7:0]) +
	( 14'sd 6058) * $signed(input_fmap_246[7:0]) +
	( 16'sd 22503) * $signed(input_fmap_247[7:0]) +
	( 16'sd 16571) * $signed(input_fmap_248[7:0]) +
	( 11'sd 800) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19567) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10174) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11243) * $signed(input_fmap_253[7:0]) +
	( 15'sd 14010) * $signed(input_fmap_254[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_67;
assign conv_mac_67 = 
	( 16'sd 23292) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27101) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8203) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7372) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29274) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30644) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27398) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24644) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19785) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2236) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18242) * $signed(input_fmap_10[7:0]) +
	( 10'sd 366) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28589) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13110) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11591) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21190) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3439) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14633) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6515) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21277) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25311) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1893) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13830) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25946) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11444) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2178) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28434) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22390) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32324) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21767) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8341) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21996) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6906) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9021) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16749) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27393) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23209) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9169) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15959) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5825) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25739) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21922) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7856) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27421) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22019) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26819) * $signed(input_fmap_48[7:0]) +
	( 10'sd 388) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22306) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6282) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27205) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22464) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9783) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5516) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10037) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2347) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23275) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30096) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18655) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26733) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20743) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18141) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16395) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19183) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13553) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14035) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7837) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12132) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30189) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30487) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30860) * $signed(input_fmap_75[7:0]) +
	( 11'sd 823) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3301) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8695) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26284) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25327) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22574) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2769) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11852) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17588) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11341) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20507) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12781) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10753) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31796) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1239) * $signed(input_fmap_92[7:0]) +
	( 11'sd 681) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10208) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26543) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26287) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5235) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15623) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20338) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26685) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1038) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20163) * $signed(input_fmap_102[7:0]) +
	( 13'sd 4019) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8199) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13230) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12857) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2959) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23114) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9806) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15366) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10134) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1541) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16520) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18226) * $signed(input_fmap_116[7:0]) +
	( 11'sd 530) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13773) * $signed(input_fmap_118[7:0]) +
	( 15'sd 16352) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14717) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31023) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2311) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11771) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19406) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18233) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27590) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32317) * $signed(input_fmap_127[7:0]) +
	( 16'sd 21893) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7805) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12527) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20793) * $signed(input_fmap_131[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31126) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21788) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20891) * $signed(input_fmap_135[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6974) * $signed(input_fmap_137[7:0]) +
	( 16'sd 20007) * $signed(input_fmap_138[7:0]) +
	( 16'sd 30392) * $signed(input_fmap_139[7:0]) +
	( 16'sd 21351) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_143[7:0]) +
	( 12'sd 1932) * $signed(input_fmap_144[7:0]) +
	( 15'sd 9604) * $signed(input_fmap_145[7:0]) +
	( 16'sd 28959) * $signed(input_fmap_146[7:0]) +
	( 16'sd 22518) * $signed(input_fmap_147[7:0]) +
	( 11'sd 836) * $signed(input_fmap_148[7:0]) +
	( 14'sd 5506) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18455) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14534) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29800) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1156) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11451) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28497) * $signed(input_fmap_155[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_156[7:0]) +
	( 15'sd 10081) * $signed(input_fmap_157[7:0]) +
	( 15'sd 13279) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26531) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_160[7:0]) +
	( 14'sd 7701) * $signed(input_fmap_161[7:0]) +
	( 14'sd 5678) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_163[7:0]) +
	( 15'sd 14468) * $signed(input_fmap_164[7:0]) +
	( 16'sd 32085) * $signed(input_fmap_165[7:0]) +
	( 12'sd 1815) * $signed(input_fmap_166[7:0]) +
	( 15'sd 14078) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17404) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_169[7:0]) +
	( 16'sd 26682) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7044) * $signed(input_fmap_171[7:0]) +
	( 16'sd 23717) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27048) * $signed(input_fmap_173[7:0]) +
	( 15'sd 9116) * $signed(input_fmap_174[7:0]) +
	( 15'sd 10302) * $signed(input_fmap_175[7:0]) +
	( 16'sd 32009) * $signed(input_fmap_176[7:0]) +
	( 16'sd 20148) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15613) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_179[7:0]) +
	( 16'sd 19331) * $signed(input_fmap_180[7:0]) +
	( 15'sd 8631) * $signed(input_fmap_181[7:0]) +
	( 15'sd 9389) * $signed(input_fmap_182[7:0]) +
	( 16'sd 16500) * $signed(input_fmap_183[7:0]) +
	( 16'sd 25990) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11029) * $signed(input_fmap_185[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22685) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32460) * $signed(input_fmap_188[7:0]) +
	( 15'sd 16370) * $signed(input_fmap_189[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_190[7:0]) +
	( 14'sd 6723) * $signed(input_fmap_191[7:0]) +
	( 14'sd 8124) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12055) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23335) * $signed(input_fmap_194[7:0]) +
	( 14'sd 6502) * $signed(input_fmap_195[7:0]) +
	( 16'sd 26299) * $signed(input_fmap_196[7:0]) +
	( 16'sd 27503) * $signed(input_fmap_197[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_198[7:0]) +
	( 13'sd 2510) * $signed(input_fmap_199[7:0]) +
	( 12'sd 1298) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1383) * $signed(input_fmap_201[7:0]) +
	( 15'sd 16176) * $signed(input_fmap_202[7:0]) +
	( 16'sd 32721) * $signed(input_fmap_203[7:0]) +
	( 16'sd 30089) * $signed(input_fmap_204[7:0]) +
	( 16'sd 22424) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31576) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5527) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15104) * $signed(input_fmap_208[7:0]) +
	( 16'sd 30533) * $signed(input_fmap_209[7:0]) +
	( 16'sd 27134) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20273) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29119) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6094) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7471) * $signed(input_fmap_214[7:0]) +
	( 16'sd 20680) * $signed(input_fmap_215[7:0]) +
	( 16'sd 31097) * $signed(input_fmap_216[7:0]) +
	( 16'sd 20796) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10189) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_219[7:0]) +
	( 16'sd 32311) * $signed(input_fmap_220[7:0]) +
	( 13'sd 3184) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25406) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19345) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27332) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_226[7:0]) +
	( 15'sd 11519) * $signed(input_fmap_227[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10591) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28115) * $signed(input_fmap_230[7:0]) +
	( 14'sd 5311) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_232[7:0]) +
	( 16'sd 31910) * $signed(input_fmap_233[7:0]) +
	( 16'sd 16833) * $signed(input_fmap_234[7:0]) +
	( 16'sd 31096) * $signed(input_fmap_235[7:0]) +
	( 16'sd 19849) * $signed(input_fmap_236[7:0]) +
	( 12'sd 1859) * $signed(input_fmap_237[7:0]) +
	( 14'sd 6981) * $signed(input_fmap_238[7:0]) +
	( 16'sd 29590) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6568) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18439) * $signed(input_fmap_241[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13432) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12348) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28749) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14528) * $signed(input_fmap_246[7:0]) +
	( 11'sd 728) * $signed(input_fmap_247[7:0]) +
	( 16'sd 16623) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12048) * $signed(input_fmap_249[7:0]) +
	( 16'sd 19953) * $signed(input_fmap_250[7:0]) +
	( 15'sd 10322) * $signed(input_fmap_251[7:0]) +
	( 16'sd 16385) * $signed(input_fmap_252[7:0]) +
	( 10'sd 333) * $signed(input_fmap_253[7:0]) +
	( 7'sd 34) * $signed(input_fmap_254[7:0]) +
	( 16'sd 31927) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_68;
assign conv_mac_68 = 
	( 16'sd 17549) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26870) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30304) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21098) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27291) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3211) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32444) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1524) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18970) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4391) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28674) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11263) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13676) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2590) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22348) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_18[7:0]) +
	( 10'sd 331) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11393) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17261) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2405) * $signed(input_fmap_22[7:0]) +
	( 11'sd 870) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9122) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24639) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7163) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24843) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22039) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15816) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3836) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4498) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23660) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19334) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29310) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20763) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6981) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16728) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23620) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18663) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21948) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3504) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7782) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3355) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_44[7:0]) +
	( 11'sd 602) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20617) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1141) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11542) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5086) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10656) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27073) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4644) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2870) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7698) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3720) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27360) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28575) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10210) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11526) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9645) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11490) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28961) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30329) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13832) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11659) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11305) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14799) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5937) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24672) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30806) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22438) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7263) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23420) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32120) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17134) * $signed(input_fmap_76[7:0]) +
	( 9'sd 193) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21110) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4247) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8084) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1560) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16264) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3864) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7593) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28813) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32094) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3931) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25255) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12674) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24460) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26008) * $signed(input_fmap_92[7:0]) +
	( 11'sd 980) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25067) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21787) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6825) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24818) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13404) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10134) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13653) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10175) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23476) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29732) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16944) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13657) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17743) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19911) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17820) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28357) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27203) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3818) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10154) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19301) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3011) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6345) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21064) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19535) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15674) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9881) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24417) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16923) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_127[7:0]) +
	( 15'sd 11094) * $signed(input_fmap_128[7:0]) +
	( 13'sd 2938) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1687) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3241) * $signed(input_fmap_131[7:0]) +
	( 15'sd 9712) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16785) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31357) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23518) * $signed(input_fmap_135[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11247) * $signed(input_fmap_137[7:0]) +
	( 16'sd 28024) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28407) * $signed(input_fmap_139[7:0]) +
	( 16'sd 22161) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29824) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8702) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10859) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6148) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21912) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9746) * $signed(input_fmap_146[7:0]) +
	( 15'sd 12573) * $signed(input_fmap_147[7:0]) +
	( 14'sd 7802) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4392) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23592) * $signed(input_fmap_150[7:0]) +
	( 16'sd 32384) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20056) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31544) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31897) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12439) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25279) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27808) * $signed(input_fmap_157[7:0]) +
	( 16'sd 31595) * $signed(input_fmap_158[7:0]) +
	( 9'sd 247) * $signed(input_fmap_159[7:0]) +
	( 15'sd 12013) * $signed(input_fmap_160[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14427) * $signed(input_fmap_162[7:0]) +
	( 15'sd 10337) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3056) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11287) * $signed(input_fmap_165[7:0]) +
	( 16'sd 16564) * $signed(input_fmap_166[7:0]) +
	( 14'sd 8186) * $signed(input_fmap_167[7:0]) +
	( 16'sd 16437) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11317) * $signed(input_fmap_169[7:0]) +
	( 16'sd 29917) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11762) * $signed(input_fmap_172[7:0]) +
	( 16'sd 21603) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17231) * $signed(input_fmap_175[7:0]) +
	( 15'sd 12610) * $signed(input_fmap_176[7:0]) +
	( 15'sd 9519) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_179[7:0]) +
	( 16'sd 31513) * $signed(input_fmap_180[7:0]) +
	( 16'sd 19312) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29300) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29341) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_185[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5418) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21822) * $signed(input_fmap_188[7:0]) +
	( 16'sd 28348) * $signed(input_fmap_189[7:0]) +
	( 15'sd 8806) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31285) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14602) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30315) * $signed(input_fmap_193[7:0]) +
	( 16'sd 17601) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13110) * $signed(input_fmap_195[7:0]) +
	( 13'sd 3299) * $signed(input_fmap_196[7:0]) +
	( 15'sd 12043) * $signed(input_fmap_197[7:0]) +
	( 14'sd 4155) * $signed(input_fmap_198[7:0]) +
	( 9'sd 223) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8823) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15689) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11759) * $signed(input_fmap_202[7:0]) +
	( 13'sd 3863) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19163) * $signed(input_fmap_204[7:0]) +
	( 13'sd 3338) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6796) * $signed(input_fmap_206[7:0]) +
	( 16'sd 26378) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7745) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5799) * $signed(input_fmap_210[7:0]) +
	( 15'sd 13214) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29480) * $signed(input_fmap_212[7:0]) +
	( 14'sd 7381) * $signed(input_fmap_213[7:0]) +
	( 16'sd 24144) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11944) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5874) * $signed(input_fmap_216[7:0]) +
	( 12'sd 2033) * $signed(input_fmap_217[7:0]) +
	( 16'sd 17962) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20906) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26035) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27657) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5276) * $signed(input_fmap_222[7:0]) +
	( 13'sd 3293) * $signed(input_fmap_223[7:0]) +
	( 16'sd 24079) * $signed(input_fmap_224[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_225[7:0]) +
	( 16'sd 16816) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27818) * $signed(input_fmap_227[7:0]) +
	( 16'sd 32338) * $signed(input_fmap_228[7:0]) +
	( 15'sd 12557) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_230[7:0]) +
	( 15'sd 15791) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9066) * $signed(input_fmap_232[7:0]) +
	( 16'sd 16812) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18439) * $signed(input_fmap_234[7:0]) +
	( 13'sd 2499) * $signed(input_fmap_235[7:0]) +
	( 16'sd 19367) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29389) * $signed(input_fmap_237[7:0]) +
	( 14'sd 7925) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13456) * $signed(input_fmap_239[7:0]) +
	( 16'sd 29044) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23799) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28412) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28482) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2109) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7696) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15774) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15518) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10400) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2819) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9364) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4233) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27473) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1763) * $signed(input_fmap_254[7:0]) +
	( 16'sd 18069) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_69;
assign conv_mac_69 = 
	( 16'sd 20335) * $signed(input_fmap_0[7:0]) +
	( 11'sd 707) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1269) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25802) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20515) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13001) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23844) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25335) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20280) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20126) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5727) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13866) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31007) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26379) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18225) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10922) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2461) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26443) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5483) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21547) * $signed(input_fmap_21[7:0]) +
	( 10'sd 477) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5753) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7426) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19507) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10981) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25601) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14572) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9517) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6579) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15842) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16757) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30806) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27645) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3454) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29758) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30660) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7232) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18844) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11317) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23941) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29069) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27502) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25564) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25408) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25486) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15763) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18019) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12671) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26954) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25378) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10261) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23116) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28195) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15267) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30434) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29349) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8354) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26850) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17586) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30861) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18592) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9337) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32581) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18752) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32606) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31066) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3617) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22946) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25045) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11378) * $signed(input_fmap_80[7:0]) +
	( 14'sd 8111) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31204) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23933) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27206) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28355) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9780) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13204) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31381) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25868) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16559) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25419) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26719) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27140) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17878) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19747) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2881) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22893) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13233) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3681) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16358) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18223) * $signed(input_fmap_102[7:0]) +
	( 10'sd 468) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15321) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19049) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26205) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29483) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18993) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24134) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14089) * $signed(input_fmap_111[7:0]) +
	( 11'sd 655) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13695) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3842) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4134) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18195) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19300) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23677) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18139) * $signed(input_fmap_119[7:0]) +
	( 10'sd 415) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14461) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12284) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14646) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6363) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21514) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21535) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28473) * $signed(input_fmap_127[7:0]) +
	( 14'sd 7374) * $signed(input_fmap_128[7:0]) +
	( 16'sd 30730) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27854) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5359) * $signed(input_fmap_131[7:0]) +
	( 13'sd 2751) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_133[7:0]) +
	( 15'sd 10793) * $signed(input_fmap_134[7:0]) +
	( 14'sd 6279) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30907) * $signed(input_fmap_136[7:0]) +
	( 14'sd 8044) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_138[7:0]) +
	( 15'sd 12807) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1808) * $signed(input_fmap_140[7:0]) +
	( 15'sd 14313) * $signed(input_fmap_141[7:0]) +
	( 15'sd 10360) * $signed(input_fmap_142[7:0]) +
	( 15'sd 8931) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13232) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2442) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29548) * $signed(input_fmap_146[7:0]) +
	( 16'sd 25740) * $signed(input_fmap_147[7:0]) +
	( 11'sd 799) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_149[7:0]) +
	( 12'sd 1775) * $signed(input_fmap_150[7:0]) +
	( 16'sd 16865) * $signed(input_fmap_151[7:0]) +
	( 11'sd 901) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2417) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10150) * $signed(input_fmap_154[7:0]) +
	( 13'sd 2178) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_156[7:0]) +
	( 16'sd 32532) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20713) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32652) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21613) * $signed(input_fmap_160[7:0]) +
	( 16'sd 32618) * $signed(input_fmap_161[7:0]) +
	( 15'sd 16024) * $signed(input_fmap_162[7:0]) +
	( 15'sd 13214) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10897) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12271) * $signed(input_fmap_165[7:0]) +
	( 16'sd 23530) * $signed(input_fmap_166[7:0]) +
	( 16'sd 27447) * $signed(input_fmap_167[7:0]) +
	( 11'sd 582) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17972) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1714) * $signed(input_fmap_172[7:0]) +
	( 15'sd 11812) * $signed(input_fmap_173[7:0]) +
	( 16'sd 18239) * $signed(input_fmap_174[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1354) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27599) * $signed(input_fmap_178[7:0]) +
	( 16'sd 32742) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4569) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28969) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16441) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17868) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24178) * $signed(input_fmap_184[7:0]) +
	( 16'sd 20172) * $signed(input_fmap_185[7:0]) +
	( 16'sd 32375) * $signed(input_fmap_186[7:0]) +
	( 15'sd 8771) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4845) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19794) * $signed(input_fmap_189[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_190[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19671) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29387) * $signed(input_fmap_193[7:0]) +
	( 15'sd 11923) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_195[7:0]) +
	( 16'sd 18599) * $signed(input_fmap_196[7:0]) +
	( 16'sd 28523) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24653) * $signed(input_fmap_198[7:0]) +
	( 13'sd 2308) * $signed(input_fmap_199[7:0]) +
	( 15'sd 9601) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22212) * $signed(input_fmap_201[7:0]) +
	( 14'sd 8001) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24483) * $signed(input_fmap_203[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_204[7:0]) +
	( 15'sd 13381) * $signed(input_fmap_205[7:0]) +
	( 16'sd 19750) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29911) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28485) * $signed(input_fmap_208[7:0]) +
	( 16'sd 32691) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4654) * $signed(input_fmap_210[7:0]) +
	( 13'sd 2678) * $signed(input_fmap_211[7:0]) +
	( 15'sd 13137) * $signed(input_fmap_212[7:0]) +
	( 16'sd 30815) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29296) * $signed(input_fmap_215[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_216[7:0]) +
	( 16'sd 29061) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7648) * $signed(input_fmap_218[7:0]) +
	( 16'sd 31104) * $signed(input_fmap_219[7:0]) +
	( 16'sd 16658) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23894) * $signed(input_fmap_221[7:0]) +
	( 16'sd 22849) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_223[7:0]) +
	( 14'sd 4478) * $signed(input_fmap_224[7:0]) +
	( 10'sd 358) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14655) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13745) * $signed(input_fmap_227[7:0]) +
	( 11'sd 584) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15417) * $signed(input_fmap_230[7:0]) +
	( 16'sd 23342) * $signed(input_fmap_231[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_232[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_233[7:0]) +
	( 15'sd 9117) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29771) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27035) * $signed(input_fmap_236[7:0]) +
	( 13'sd 3596) * $signed(input_fmap_237[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_238[7:0]) +
	( 15'sd 14372) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23233) * $signed(input_fmap_240[7:0]) +
	( 15'sd 10971) * $signed(input_fmap_241[7:0]) +
	( 15'sd 14874) * $signed(input_fmap_242[7:0]) +
	( 15'sd 15078) * $signed(input_fmap_243[7:0]) +
	( 16'sd 23686) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28620) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19221) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20284) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4399) * $signed(input_fmap_248[7:0]) +
	( 16'sd 31647) * $signed(input_fmap_249[7:0]) +
	( 16'sd 18277) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21766) * $signed(input_fmap_251[7:0]) +
	( 10'sd 399) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6102) * $signed(input_fmap_253[7:0]) +
	( 14'sd 6201) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14085) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_70;
assign conv_mac_70 = 
	( 16'sd 16645) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29005) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19032) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6223) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16802) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20879) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7254) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20877) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3894) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29525) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8822) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8922) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8307) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13033) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13207) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25743) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30387) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6345) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11437) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28868) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19606) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21301) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22634) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3654) * $signed(input_fmap_25[7:0]) +
	( 7'sd 37) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30927) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14875) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9836) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3033) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25553) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4897) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27194) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17518) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12055) * $signed(input_fmap_36[7:0]) +
	( 11'sd 690) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28544) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30188) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4995) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6267) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27484) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3033) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15498) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32263) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13543) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4736) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28375) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17339) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1692) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14566) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21990) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31501) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5939) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13552) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15872) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26166) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16042) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6136) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26159) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13090) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13891) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30474) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18169) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30545) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5681) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18607) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24266) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28620) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28448) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9057) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20778) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30928) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3154) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4925) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27365) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27679) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26843) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31201) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3951) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22533) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32256) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10761) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4294) * $signed(input_fmap_93[7:0]) +
	( 14'sd 8126) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10977) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20514) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4273) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2300) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5911) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6102) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11138) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1245) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7873) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23219) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9675) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19095) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4838) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17849) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8653) * $signed(input_fmap_112[7:0]) +
	( 11'sd 888) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13959) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16874) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29211) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22587) * $signed(input_fmap_121[7:0]) +
	( 8'sd 107) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10563) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5830) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29590) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12710) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27889) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13171) * $signed(input_fmap_128[7:0]) +
	( 14'sd 6961) * $signed(input_fmap_129[7:0]) +
	( 15'sd 9512) * $signed(input_fmap_130[7:0]) +
	( 16'sd 22462) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11201) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21683) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25129) * $signed(input_fmap_134[7:0]) +
	( 16'sd 24854) * $signed(input_fmap_135[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15821) * $signed(input_fmap_137[7:0]) +
	( 12'sd 1796) * $signed(input_fmap_138[7:0]) +
	( 16'sd 25389) * $signed(input_fmap_139[7:0]) +
	( 16'sd 16921) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10708) * $signed(input_fmap_141[7:0]) +
	( 15'sd 10677) * $signed(input_fmap_142[7:0]) +
	( 14'sd 8131) * $signed(input_fmap_143[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2915) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15589) * $signed(input_fmap_146[7:0]) +
	( 15'sd 12739) * $signed(input_fmap_147[7:0]) +
	( 16'sd 27683) * $signed(input_fmap_148[7:0]) +
	( 16'sd 22263) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31515) * $signed(input_fmap_150[7:0]) +
	( 16'sd 31402) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2675) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23045) * $signed(input_fmap_154[7:0]) +
	( 12'sd 1477) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7063) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31907) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11108) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_159[7:0]) +
	( 15'sd 9356) * $signed(input_fmap_160[7:0]) +
	( 15'sd 10073) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27223) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_163[7:0]) +
	( 12'sd 2007) * $signed(input_fmap_164[7:0]) +
	( 14'sd 5832) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4983) * $signed(input_fmap_166[7:0]) +
	( 16'sd 19393) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4276) * $signed(input_fmap_168[7:0]) +
	( 14'sd 8068) * $signed(input_fmap_169[7:0]) +
	( 16'sd 27397) * $signed(input_fmap_170[7:0]) +
	( 16'sd 17741) * $signed(input_fmap_171[7:0]) +
	( 14'sd 5447) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29050) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7524) * $signed(input_fmap_174[7:0]) +
	( 16'sd 27769) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27766) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1854) * $signed(input_fmap_177[7:0]) +
	( 14'sd 6032) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20182) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21971) * $signed(input_fmap_180[7:0]) +
	( 15'sd 9101) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_182[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_183[7:0]) +
	( 10'sd 505) * $signed(input_fmap_184[7:0]) +
	( 15'sd 14816) * $signed(input_fmap_185[7:0]) +
	( 16'sd 24294) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11062) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11766) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17005) * $signed(input_fmap_190[7:0]) +
	( 15'sd 11579) * $signed(input_fmap_191[7:0]) +
	( 16'sd 23440) * $signed(input_fmap_192[7:0]) +
	( 16'sd 25537) * $signed(input_fmap_193[7:0]) +
	( 16'sd 28513) * $signed(input_fmap_194[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_195[7:0]) +
	( 14'sd 8017) * $signed(input_fmap_196[7:0]) +
	( 16'sd 17731) * $signed(input_fmap_197[7:0]) +
	( 16'sd 30459) * $signed(input_fmap_198[7:0]) +
	( 16'sd 19711) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29861) * $signed(input_fmap_200[7:0]) +
	( 14'sd 4730) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7876) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_203[7:0]) +
	( 14'sd 7470) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30044) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13493) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22458) * $signed(input_fmap_208[7:0]) +
	( 14'sd 8014) * $signed(input_fmap_209[7:0]) +
	( 16'sd 21971) * $signed(input_fmap_210[7:0]) +
	( 16'sd 31086) * $signed(input_fmap_211[7:0]) +
	( 9'sd 235) * $signed(input_fmap_212[7:0]) +
	( 16'sd 16830) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17534) * $signed(input_fmap_215[7:0]) +
	( 16'sd 21444) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10125) * $signed(input_fmap_217[7:0]) +
	( 13'sd 3534) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21805) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4165) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1938) * $signed(input_fmap_221[7:0]) +
	( 16'sd 32269) * $signed(input_fmap_222[7:0]) +
	( 16'sd 27254) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14039) * $signed(input_fmap_224[7:0]) +
	( 14'sd 7633) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31404) * $signed(input_fmap_226[7:0]) +
	( 16'sd 16991) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25946) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8828) * $signed(input_fmap_229[7:0]) +
	( 16'sd 16640) * $signed(input_fmap_230[7:0]) +
	( 15'sd 8789) * $signed(input_fmap_231[7:0]) +
	( 16'sd 17027) * $signed(input_fmap_232[7:0]) +
	( 16'sd 32013) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15420) * $signed(input_fmap_234[7:0]) +
	( 15'sd 8553) * $signed(input_fmap_235[7:0]) +
	( 15'sd 14518) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19003) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13517) * $signed(input_fmap_239[7:0]) +
	( 11'sd 658) * $signed(input_fmap_240[7:0]) +
	( 12'sd 1197) * $signed(input_fmap_241[7:0]) +
	( 16'sd 31988) * $signed(input_fmap_242[7:0]) +
	( 16'sd 19670) * $signed(input_fmap_243[7:0]) +
	( 16'sd 27749) * $signed(input_fmap_244[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14787) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17549) * $signed(input_fmap_247[7:0]) +
	( 13'sd 2740) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30994) * $signed(input_fmap_249[7:0]) +
	( 16'sd 16893) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15278) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12921) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11878) * $signed(input_fmap_253[7:0]) +
	( 13'sd 4062) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11052) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_71;
assign conv_mac_71 = 
	( 16'sd 27338) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29228) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26044) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15369) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2726) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6716) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6611) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28312) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29690) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12612) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30996) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22557) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32251) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3131) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14672) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22374) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29618) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30317) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5331) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4904) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3816) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20033) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12028) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27243) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8857) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15890) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1468) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10236) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28806) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6546) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32115) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22191) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2751) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1047) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32204) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23324) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25254) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27063) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12150) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20449) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19338) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18217) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12312) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7178) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2187) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24133) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6443) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11743) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18235) * $signed(input_fmap_54[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2560) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27165) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1628) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10901) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31676) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30762) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22318) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30155) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11166) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23372) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31521) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32450) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15560) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30205) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14664) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21639) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8302) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1519) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30021) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24099) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26075) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3338) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21547) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13632) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32162) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11121) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9438) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20835) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13987) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28668) * $signed(input_fmap_86[7:0]) +
	( 11'sd 965) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20151) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23608) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23958) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25329) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5509) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14424) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28657) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28464) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8879) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13465) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10259) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6161) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16965) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23670) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2151) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22483) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16931) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28339) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13075) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18636) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15889) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20203) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2169) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7379) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30468) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19592) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5301) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15758) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1235) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2512) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29780) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20828) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5188) * $signed(input_fmap_126[7:0]) +
	( 11'sd 1020) * $signed(input_fmap_127[7:0]) +
	( 14'sd 5147) * $signed(input_fmap_128[7:0]) +
	( 16'sd 22837) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14396) * $signed(input_fmap_130[7:0]) +
	( 15'sd 12725) * $signed(input_fmap_131[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_132[7:0]) +
	( 14'sd 8094) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1973) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32765) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8421) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4582) * $signed(input_fmap_137[7:0]) +
	( 15'sd 8917) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14237) * $signed(input_fmap_139[7:0]) +
	( 16'sd 31235) * $signed(input_fmap_140[7:0]) +
	( 16'sd 30751) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22934) * $signed(input_fmap_142[7:0]) +
	( 15'sd 11889) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28744) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25737) * $signed(input_fmap_145[7:0]) +
	( 16'sd 22959) * $signed(input_fmap_146[7:0]) +
	( 16'sd 28125) * $signed(input_fmap_147[7:0]) +
	( 16'sd 31156) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4550) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5035) * $signed(input_fmap_150[7:0]) +
	( 15'sd 11287) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21032) * $signed(input_fmap_152[7:0]) +
	( 16'sd 19809) * $signed(input_fmap_153[7:0]) +
	( 16'sd 21977) * $signed(input_fmap_154[7:0]) +
	( 14'sd 4997) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17962) * $signed(input_fmap_156[7:0]) +
	( 16'sd 28560) * $signed(input_fmap_157[7:0]) +
	( 16'sd 26540) * $signed(input_fmap_158[7:0]) +
	( 16'sd 23061) * $signed(input_fmap_159[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_160[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26135) * $signed(input_fmap_162[7:0]) +
	( 16'sd 25021) * $signed(input_fmap_163[7:0]) +
	( 16'sd 27478) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23223) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31236) * $signed(input_fmap_166[7:0]) +
	( 15'sd 8536) * $signed(input_fmap_167[7:0]) +
	( 15'sd 16127) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30354) * $signed(input_fmap_169[7:0]) +
	( 15'sd 12491) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24862) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3583) * $signed(input_fmap_172[7:0]) +
	( 16'sd 24040) * $signed(input_fmap_173[7:0]) +
	( 16'sd 22187) * $signed(input_fmap_174[7:0]) +
	( 15'sd 14138) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_177[7:0]) +
	( 16'sd 28872) * $signed(input_fmap_178[7:0]) +
	( 16'sd 23769) * $signed(input_fmap_179[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_180[7:0]) +
	( 15'sd 10393) * $signed(input_fmap_181[7:0]) +
	( 16'sd 28477) * $signed(input_fmap_182[7:0]) +
	( 16'sd 24793) * $signed(input_fmap_183[7:0]) +
	( 14'sd 7559) * $signed(input_fmap_184[7:0]) +
	( 15'sd 9209) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13116) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22076) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_188[7:0]) +
	( 16'sd 23514) * $signed(input_fmap_189[7:0]) +
	( 13'sd 3636) * $signed(input_fmap_190[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29524) * $signed(input_fmap_192[7:0]) +
	( 13'sd 2848) * $signed(input_fmap_193[7:0]) +
	( 16'sd 31033) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19989) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24649) * $signed(input_fmap_196[7:0]) +
	( 16'sd 23562) * $signed(input_fmap_197[7:0]) +
	( 15'sd 15354) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24953) * $signed(input_fmap_199[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21634) * $signed(input_fmap_201[7:0]) +
	( 16'sd 16494) * $signed(input_fmap_202[7:0]) +
	( 15'sd 9708) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2491) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24599) * $signed(input_fmap_205[7:0]) +
	( 16'sd 22129) * $signed(input_fmap_206[7:0]) +
	( 13'sd 2220) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12314) * $signed(input_fmap_208[7:0]) +
	( 16'sd 16997) * $signed(input_fmap_209[7:0]) +
	( 14'sd 8051) * $signed(input_fmap_210[7:0]) +
	( 12'sd 1806) * $signed(input_fmap_211[7:0]) +
	( 16'sd 31971) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2806) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30525) * $signed(input_fmap_214[7:0]) +
	( 16'sd 32470) * $signed(input_fmap_215[7:0]) +
	( 14'sd 6394) * $signed(input_fmap_216[7:0]) +
	( 16'sd 21050) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22024) * $signed(input_fmap_218[7:0]) +
	( 16'sd 29078) * $signed(input_fmap_219[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_220[7:0]) +
	( 16'sd 31414) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15307) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12131) * $signed(input_fmap_223[7:0]) +
	( 16'sd 31111) * $signed(input_fmap_224[7:0]) +
	( 14'sd 7537) * $signed(input_fmap_225[7:0]) +
	( 16'sd 23449) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22676) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4960) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17525) * $signed(input_fmap_229[7:0]) +
	( 15'sd 11057) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3518) * $signed(input_fmap_231[7:0]) +
	( 16'sd 32348) * $signed(input_fmap_232[7:0]) +
	( 16'sd 29693) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3278) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14738) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28093) * $signed(input_fmap_236[7:0]) +
	( 15'sd 15688) * $signed(input_fmap_237[7:0]) +
	( 16'sd 21413) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13439) * $signed(input_fmap_239[7:0]) +
	( 16'sd 32408) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30750) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27512) * $signed(input_fmap_242[7:0]) +
	( 13'sd 3024) * $signed(input_fmap_243[7:0]) +
	( 16'sd 25155) * $signed(input_fmap_244[7:0]) +
	( 12'sd 1739) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22213) * $signed(input_fmap_246[7:0]) +
	( 15'sd 14248) * $signed(input_fmap_247[7:0]) +
	( 15'sd 16191) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3231) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9510) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19340) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20907) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24458) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10504) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_72;
assign conv_mac_72 = 
	( 15'sd 15659) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11626) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11058) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18527) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16482) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3875) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24150) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13028) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6397) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30074) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27393) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3038) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28229) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1079) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20867) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13831) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14483) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15306) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6293) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6832) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3977) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10971) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12424) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7780) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13956) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24766) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14015) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13380) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26579) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6927) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21128) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28108) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18946) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19705) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30244) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_37[7:0]) +
	( 14'sd 8063) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17538) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29699) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23477) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30294) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11552) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28336) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28961) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27261) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20174) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13082) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8897) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31390) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6367) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26854) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21038) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19670) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23641) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12337) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21390) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28395) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2631) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10368) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10326) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18757) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2616) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11908) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19574) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15856) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12627) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22217) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21979) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10988) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15765) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28218) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32591) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23590) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10986) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13208) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29193) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14566) * $signed(input_fmap_84[7:0]) +
	( 10'sd 471) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30681) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27683) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20051) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21999) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19393) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28477) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21035) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5701) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23525) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21451) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17590) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19136) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21614) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9060) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9609) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30109) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5653) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23999) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32560) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7033) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24011) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2243) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6326) * $signed(input_fmap_110[7:0]) +
	( 6'sd 19) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1274) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18065) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20880) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6995) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7070) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6698) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15501) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9099) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11591) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3675) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25032) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26665) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7786) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23277) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2824) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18459) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19425) * $signed(input_fmap_129[7:0]) +
	( 10'sd 505) * $signed(input_fmap_130[7:0]) +
	( 16'sd 28847) * $signed(input_fmap_131[7:0]) +
	( 9'sd 148) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11424) * $signed(input_fmap_133[7:0]) +
	( 16'sd 17673) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19082) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25697) * $signed(input_fmap_136[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_137[7:0]) +
	( 13'sd 3892) * $signed(input_fmap_138[7:0]) +
	( 15'sd 13996) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18687) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25961) * $signed(input_fmap_142[7:0]) +
	( 16'sd 27642) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22762) * $signed(input_fmap_144[7:0]) +
	( 16'sd 16779) * $signed(input_fmap_145[7:0]) +
	( 13'sd 2561) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21382) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21160) * $signed(input_fmap_148[7:0]) +
	( 16'sd 19720) * $signed(input_fmap_149[7:0]) +
	( 9'sd 202) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3568) * $signed(input_fmap_151[7:0]) +
	( 15'sd 9523) * $signed(input_fmap_152[7:0]) +
	( 15'sd 16082) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24675) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7279) * $signed(input_fmap_155[7:0]) +
	( 14'sd 8009) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24084) * $signed(input_fmap_157[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32696) * $signed(input_fmap_159[7:0]) +
	( 12'sd 2034) * $signed(input_fmap_160[7:0]) +
	( 16'sd 18493) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4597) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3940) * $signed(input_fmap_163[7:0]) +
	( 16'sd 26760) * $signed(input_fmap_164[7:0]) +
	( 11'sd 1003) * $signed(input_fmap_165[7:0]) +
	( 16'sd 27226) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7836) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29705) * $signed(input_fmap_168[7:0]) +
	( 14'sd 5473) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_170[7:0]) +
	( 15'sd 10455) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11827) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5352) * $signed(input_fmap_173[7:0]) +
	( 11'sd 1016) * $signed(input_fmap_174[7:0]) +
	( 10'sd 291) * $signed(input_fmap_175[7:0]) +
	( 10'sd 258) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7736) * $signed(input_fmap_177[7:0]) +
	( 16'sd 29709) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18499) * $signed(input_fmap_179[7:0]) +
	( 16'sd 25091) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19313) * $signed(input_fmap_182[7:0]) +
	( 16'sd 22065) * $signed(input_fmap_183[7:0]) +
	( 16'sd 29611) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26629) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12023) * $signed(input_fmap_186[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_187[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25836) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20645) * $signed(input_fmap_190[7:0]) +
	( 16'sd 28925) * $signed(input_fmap_191[7:0]) +
	( 16'sd 16959) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15052) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12624) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25139) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11547) * $signed(input_fmap_196[7:0]) +
	( 14'sd 6463) * $signed(input_fmap_197[7:0]) +
	( 16'sd 21458) * $signed(input_fmap_198[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6426) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16819) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14827) * $signed(input_fmap_202[7:0]) +
	( 15'sd 14651) * $signed(input_fmap_203[7:0]) +
	( 14'sd 8170) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_205[7:0]) +
	( 12'sd 1194) * $signed(input_fmap_206[7:0]) +
	( 14'sd 8047) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17915) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3848) * $signed(input_fmap_209[7:0]) +
	( 15'sd 14683) * $signed(input_fmap_210[7:0]) +
	( 16'sd 29866) * $signed(input_fmap_211[7:0]) +
	( 14'sd 6328) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12145) * $signed(input_fmap_213[7:0]) +
	( 15'sd 12102) * $signed(input_fmap_214[7:0]) +
	( 16'sd 18558) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24838) * $signed(input_fmap_216[7:0]) +
	( 16'sd 18449) * $signed(input_fmap_217[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14648) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28475) * $signed(input_fmap_221[7:0]) +
	( 14'sd 6766) * $signed(input_fmap_222[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_223[7:0]) +
	( 13'sd 3829) * $signed(input_fmap_224[7:0]) +
	( 16'sd 19997) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32206) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6437) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25350) * $signed(input_fmap_228[7:0]) +
	( 16'sd 30014) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27279) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20204) * $signed(input_fmap_231[7:0]) +
	( 16'sd 25956) * $signed(input_fmap_232[7:0]) +
	( 15'sd 16196) * $signed(input_fmap_233[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_235[7:0]) +
	( 16'sd 16791) * $signed(input_fmap_236[7:0]) +
	( 14'sd 4131) * $signed(input_fmap_237[7:0]) +
	( 14'sd 6988) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26849) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26017) * $signed(input_fmap_240[7:0]) +
	( 16'sd 31737) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29915) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23231) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19697) * $signed(input_fmap_244[7:0]) +
	( 16'sd 31432) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_246[7:0]) +
	( 16'sd 26657) * $signed(input_fmap_247[7:0]) +
	( 16'sd 16674) * $signed(input_fmap_248[7:0]) +
	( 7'sd 41) * $signed(input_fmap_249[7:0]) +
	( 16'sd 18697) * $signed(input_fmap_250[7:0]) +
	( 16'sd 25365) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_252[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10587) * $signed(input_fmap_254[7:0]) +
	( 16'sd 16522) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_73;
assign conv_mac_73 = 
	( 15'sd 12382) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24693) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8428) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31609) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17174) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26239) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6465) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3212) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18603) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24701) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9028) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9917) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16918) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2154) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9944) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14729) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7826) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28043) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32399) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24240) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19834) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12212) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16658) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27943) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12060) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15381) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19500) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24743) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3465) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20671) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6273) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26829) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22590) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28737) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19382) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20964) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10354) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24660) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2836) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28431) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9885) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5936) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31019) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13378) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11446) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18368) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21799) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20674) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17599) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16030) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12059) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8150) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4531) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4814) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7519) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15928) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23739) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21017) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4402) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15031) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24317) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11605) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27475) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18128) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25559) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3752) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7446) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26717) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32189) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9626) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30840) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29868) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17977) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18996) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15481) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25431) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6018) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28562) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20953) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19663) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9601) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3605) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19379) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3599) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14936) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15058) * $signed(input_fmap_99[7:0]) +
	( 11'sd 784) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15705) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31231) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19448) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22949) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20949) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8793) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18228) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17478) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11298) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2368) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3765) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20684) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3876) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32399) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25136) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17710) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5251) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5095) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22108) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8523) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9447) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4620) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6699) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18132) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19439) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19799) * $signed(input_fmap_130[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8323) * $signed(input_fmap_132[7:0]) +
	( 15'sd 15272) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5004) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20992) * $signed(input_fmap_135[7:0]) +
	( 16'sd 19677) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4179) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27156) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28768) * $signed(input_fmap_139[7:0]) +
	( 15'sd 12239) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24085) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27255) * $signed(input_fmap_142[7:0]) +
	( 16'sd 21361) * $signed(input_fmap_143[7:0]) +
	( 12'sd 1038) * $signed(input_fmap_144[7:0]) +
	( 14'sd 6808) * $signed(input_fmap_145[7:0]) +
	( 16'sd 28449) * $signed(input_fmap_146[7:0]) +
	( 16'sd 32523) * $signed(input_fmap_147[7:0]) +
	( 16'sd 31469) * $signed(input_fmap_148[7:0]) +
	( 16'sd 24623) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18796) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23731) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23242) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23628) * $signed(input_fmap_153[7:0]) +
	( 15'sd 12822) * $signed(input_fmap_154[7:0]) +
	( 16'sd 31386) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28214) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22096) * $signed(input_fmap_157[7:0]) +
	( 11'sd 571) * $signed(input_fmap_158[7:0]) +
	( 15'sd 15159) * $signed(input_fmap_159[7:0]) +
	( 14'sd 7301) * $signed(input_fmap_160[7:0]) +
	( 16'sd 25904) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10190) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22216) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11700) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4422) * $signed(input_fmap_166[7:0]) +
	( 11'sd 701) * $signed(input_fmap_167[7:0]) +
	( 16'sd 22396) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3818) * $signed(input_fmap_169[7:0]) +
	( 15'sd 12710) * $signed(input_fmap_170[7:0]) +
	( 16'sd 27364) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15559) * $signed(input_fmap_172[7:0]) +
	( 16'sd 25131) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14949) * $signed(input_fmap_174[7:0]) +
	( 16'sd 29678) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15839) * $signed(input_fmap_176[7:0]) +
	( 14'sd 4422) * $signed(input_fmap_177[7:0]) +
	( 16'sd 19045) * $signed(input_fmap_178[7:0]) +
	( 15'sd 10814) * $signed(input_fmap_179[7:0]) +
	( 15'sd 8922) * $signed(input_fmap_180[7:0]) +
	( 16'sd 21948) * $signed(input_fmap_181[7:0]) +
	( 11'sd 698) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29830) * $signed(input_fmap_183[7:0]) +
	( 8'sd 91) * $signed(input_fmap_184[7:0]) +
	( 16'sd 29887) * $signed(input_fmap_185[7:0]) +
	( 16'sd 22205) * $signed(input_fmap_186[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_187[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7375) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17651) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20479) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15312) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20093) * $signed(input_fmap_193[7:0]) +
	( 16'sd 22180) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22596) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_196[7:0]) +
	( 16'sd 16904) * $signed(input_fmap_197[7:0]) +
	( 16'sd 26698) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13103) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15644) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21145) * $signed(input_fmap_203[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_204[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29135) * $signed(input_fmap_206[7:0]) +
	( 16'sd 31709) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11940) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22770) * $signed(input_fmap_209[7:0]) +
	( 15'sd 12885) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20008) * $signed(input_fmap_211[7:0]) +
	( 15'sd 13839) * $signed(input_fmap_212[7:0]) +
	( 16'sd 20853) * $signed(input_fmap_213[7:0]) +
	( 15'sd 16237) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25105) * $signed(input_fmap_215[7:0]) +
	( 13'sd 2502) * $signed(input_fmap_216[7:0]) +
	( 13'sd 4038) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8885) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17642) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_220[7:0]) +
	( 16'sd 31920) * $signed(input_fmap_221[7:0]) +
	( 16'sd 29535) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8313) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17005) * $signed(input_fmap_224[7:0]) +
	( 10'sd 295) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29502) * $signed(input_fmap_226[7:0]) +
	( 16'sd 25576) * $signed(input_fmap_227[7:0]) +
	( 16'sd 30150) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_229[7:0]) +
	( 16'sd 21113) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13805) * $signed(input_fmap_231[7:0]) +
	( 16'sd 27881) * $signed(input_fmap_232[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_233[7:0]) +
	( 16'sd 31066) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12614) * $signed(input_fmap_235[7:0]) +
	( 13'sd 3393) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20641) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3307) * $signed(input_fmap_238[7:0]) +
	( 16'sd 30654) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22121) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23912) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26817) * $signed(input_fmap_242[7:0]) +
	( 16'sd 24741) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20059) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19715) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23792) * $signed(input_fmap_246[7:0]) +
	( 15'sd 16060) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13246) * $signed(input_fmap_248[7:0]) +
	( 16'sd 22568) * $signed(input_fmap_249[7:0]) +
	( 14'sd 4455) * $signed(input_fmap_250[7:0]) +
	( 16'sd 20793) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20181) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29961) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11121) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_74;
assign conv_mac_74 = 
	( 15'sd 13213) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16547) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29781) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2669) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14697) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17301) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28587) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21820) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8527) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17188) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31952) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23199) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30002) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32344) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15891) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23451) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8987) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12368) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23235) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15535) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20274) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9904) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3664) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21708) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28968) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12198) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21810) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20179) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17391) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14423) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32081) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22174) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10820) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29082) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32516) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32755) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18248) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13972) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13824) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31731) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30248) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4683) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26539) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31483) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13990) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1473) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23306) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26452) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9855) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14662) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26757) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26162) * $signed(input_fmap_66[7:0]) +
	( 10'sd 281) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13625) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25114) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1501) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10494) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14268) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6745) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23685) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5269) * $signed(input_fmap_75[7:0]) +
	( 16'sd 28320) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32653) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11838) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8293) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18831) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28304) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13265) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12173) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8431) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29850) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14497) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2811) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18571) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13557) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14325) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30118) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31395) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19760) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7499) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18620) * $signed(input_fmap_97[7:0]) +
	( 13'sd 4031) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30212) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1353) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8356) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6769) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23838) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19510) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21951) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28133) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23897) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9703) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8806) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25883) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6156) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28262) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6198) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32061) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27042) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20643) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17132) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18151) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11651) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27679) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9351) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31017) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2737) * $signed(input_fmap_128[7:0]) +
	( 16'sd 16996) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6583) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5357) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8955) * $signed(input_fmap_132[7:0]) +
	( 16'sd 24528) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25327) * $signed(input_fmap_134[7:0]) +
	( 15'sd 11518) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4331) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6982) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29119) * $signed(input_fmap_138[7:0]) +
	( 15'sd 10811) * $signed(input_fmap_139[7:0]) +
	( 16'sd 25608) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20563) * $signed(input_fmap_141[7:0]) +
	( 16'sd 18737) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12638) * $signed(input_fmap_143[7:0]) +
	( 15'sd 15786) * $signed(input_fmap_144[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18387) * $signed(input_fmap_146[7:0]) +
	( 15'sd 10711) * $signed(input_fmap_147[7:0]) +
	( 15'sd 8612) * $signed(input_fmap_148[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_149[7:0]) +
	( 16'sd 20972) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4408) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7563) * $signed(input_fmap_152[7:0]) +
	( 14'sd 5272) * $signed(input_fmap_153[7:0]) +
	( 16'sd 27760) * $signed(input_fmap_154[7:0]) +
	( 16'sd 32598) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_156[7:0]) +
	( 13'sd 4015) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1274) * $signed(input_fmap_158[7:0]) +
	( 15'sd 13179) * $signed(input_fmap_159[7:0]) +
	( 15'sd 14844) * $signed(input_fmap_160[7:0]) +
	( 11'sd 783) * $signed(input_fmap_161[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20247) * $signed(input_fmap_163[7:0]) +
	( 16'sd 28966) * $signed(input_fmap_164[7:0]) +
	( 16'sd 31179) * $signed(input_fmap_165[7:0]) +
	( 14'sd 7359) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9133) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3603) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31772) * $signed(input_fmap_170[7:0]) +
	( 14'sd 4722) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_172[7:0]) +
	( 13'sd 2882) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26605) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_175[7:0]) +
	( 14'sd 4721) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19886) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10270) * $signed(input_fmap_178[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29059) * $signed(input_fmap_180[7:0]) +
	( 15'sd 12118) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12895) * $signed(input_fmap_182[7:0]) +
	( 15'sd 11419) * $signed(input_fmap_183[7:0]) +
	( 14'sd 6684) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3894) * $signed(input_fmap_185[7:0]) +
	( 12'sd 1316) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18653) * $signed(input_fmap_187[7:0]) +
	( 16'sd 27676) * $signed(input_fmap_188[7:0]) +
	( 16'sd 31346) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23542) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29317) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27680) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12386) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27075) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25260) * $signed(input_fmap_196[7:0]) +
	( 14'sd 6597) * $signed(input_fmap_197[7:0]) +
	( 16'sd 32320) * $signed(input_fmap_198[7:0]) +
	( 16'sd 19660) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25946) * $signed(input_fmap_200[7:0]) +
	( 16'sd 30051) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5952) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5742) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30387) * $signed(input_fmap_205[7:0]) +
	( 15'sd 10369) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28242) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28428) * $signed(input_fmap_208[7:0]) +
	( 16'sd 30523) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5306) * $signed(input_fmap_210[7:0]) +
	( 13'sd 2091) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12207) * $signed(input_fmap_212[7:0]) +
	( 10'sd 439) * $signed(input_fmap_213[7:0]) +
	( 16'sd 32702) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1477) * $signed(input_fmap_215[7:0]) +
	( 15'sd 9788) * $signed(input_fmap_216[7:0]) +
	( 16'sd 28946) * $signed(input_fmap_217[7:0]) +
	( 16'sd 17717) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12057) * $signed(input_fmap_219[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_221[7:0]) +
	( 16'sd 31845) * $signed(input_fmap_222[7:0]) +
	( 15'sd 16222) * $signed(input_fmap_223[7:0]) +
	( 15'sd 10441) * $signed(input_fmap_224[7:0]) +
	( 16'sd 16803) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32735) * $signed(input_fmap_226[7:0]) +
	( 16'sd 21425) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23497) * $signed(input_fmap_229[7:0]) +
	( 16'sd 22451) * $signed(input_fmap_230[7:0]) +
	( 16'sd 27653) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14527) * $signed(input_fmap_232[7:0]) +
	( 16'sd 26914) * $signed(input_fmap_233[7:0]) +
	( 15'sd 12204) * $signed(input_fmap_234[7:0]) +
	( 11'sd 945) * $signed(input_fmap_235[7:0]) +
	( 13'sd 3697) * $signed(input_fmap_236[7:0]) +
	( 16'sd 26762) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_238[7:0]) +
	( 14'sd 4358) * $signed(input_fmap_239[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32107) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26828) * $signed(input_fmap_242[7:0]) +
	( 16'sd 24346) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2154) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7057) * $signed(input_fmap_245[7:0]) +
	( 15'sd 16249) * $signed(input_fmap_246[7:0]) +
	( 16'sd 25047) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3810) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25781) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32208) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13301) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26227) * $signed(input_fmap_254[7:0]) +
	( 13'sd 2286) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_75;
assign conv_mac_75 = 
	( 16'sd 26247) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10027) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25476) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3833) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4993) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12942) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29065) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13520) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22567) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4442) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20333) * $signed(input_fmap_13[7:0]) +
	( 9'sd 215) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10853) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5164) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9966) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20138) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12670) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14184) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32485) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14850) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6321) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18414) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16277) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13298) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1794) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27763) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6213) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24725) * $signed(input_fmap_34[7:0]) +
	( 11'sd 904) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14806) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26742) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19575) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16709) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12184) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20094) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11343) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31843) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22411) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12922) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24234) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18933) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20813) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15934) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26696) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1881) * $signed(input_fmap_53[7:0]) +
	( 9'sd 171) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22902) * $signed(input_fmap_55[7:0]) +
	( 15'sd 16120) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23580) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32561) * $signed(input_fmap_58[7:0]) +
	( 11'sd 886) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32358) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5365) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26442) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27504) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29868) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28248) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15206) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20114) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23414) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30456) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17000) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13842) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10853) * $signed(input_fmap_72[7:0]) +
	( 15'sd 13380) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32232) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31975) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29433) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14037) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25289) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13445) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17499) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10783) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6979) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3349) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30360) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13671) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2229) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2479) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2541) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21502) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10865) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14946) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1959) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29261) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1507) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31476) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14291) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24136) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3051) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16570) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28130) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29431) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20073) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26563) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9854) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1668) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25773) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16530) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32597) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23230) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30128) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30669) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20792) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5821) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26670) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21801) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1777) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13962) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27236) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10216) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21690) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20498) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13562) * $signed(input_fmap_128[7:0]) +
	( 15'sd 12658) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18829) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14322) * $signed(input_fmap_131[7:0]) +
	( 14'sd 7529) * $signed(input_fmap_132[7:0]) +
	( 15'sd 13979) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5676) * $signed(input_fmap_134[7:0]) +
	( 15'sd 12522) * $signed(input_fmap_135[7:0]) +
	( 16'sd 19117) * $signed(input_fmap_136[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10329) * $signed(input_fmap_138[7:0]) +
	( 14'sd 6581) * $signed(input_fmap_139[7:0]) +
	( 14'sd 8161) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10384) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28429) * $signed(input_fmap_142[7:0]) +
	( 16'sd 27432) * $signed(input_fmap_143[7:0]) +
	( 13'sd 4047) * $signed(input_fmap_144[7:0]) +
	( 14'sd 6700) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29507) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3904) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22351) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17234) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27506) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14096) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1954) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6703) * $signed(input_fmap_154[7:0]) +
	( 16'sd 24409) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7962) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24700) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17662) * $signed(input_fmap_158[7:0]) +
	( 15'sd 13853) * $signed(input_fmap_159[7:0]) +
	( 15'sd 15071) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1862) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26686) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22109) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1051) * $signed(input_fmap_164[7:0]) +
	( 15'sd 16382) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12108) * $signed(input_fmap_166[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_167[7:0]) +
	( 16'sd 22131) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10261) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11692) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20605) * $signed(input_fmap_171[7:0]) +
	( 13'sd 2399) * $signed(input_fmap_172[7:0]) +
	( 15'sd 8303) * $signed(input_fmap_173[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_174[7:0]) +
	( 15'sd 12392) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29473) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22985) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31436) * $signed(input_fmap_178[7:0]) +
	( 16'sd 30443) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6793) * $signed(input_fmap_181[7:0]) +
	( 12'sd 1436) * $signed(input_fmap_182[7:0]) +
	( 16'sd 26998) * $signed(input_fmap_183[7:0]) +
	( 15'sd 10315) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25836) * $signed(input_fmap_185[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27752) * $signed(input_fmap_187[7:0]) +
	( 16'sd 27695) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19758) * $signed(input_fmap_189[7:0]) +
	( 15'sd 12455) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14002) * $signed(input_fmap_191[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22981) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27398) * $signed(input_fmap_194[7:0]) +
	( 14'sd 4289) * $signed(input_fmap_195[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15940) * $signed(input_fmap_197[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5214) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5372) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21076) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19920) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12275) * $signed(input_fmap_203[7:0]) +
	( 14'sd 8144) * $signed(input_fmap_204[7:0]) +
	( 14'sd 4278) * $signed(input_fmap_205[7:0]) +
	( 16'sd 24463) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12103) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25758) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14299) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10454) * $signed(input_fmap_210[7:0]) +
	( 14'sd 4669) * $signed(input_fmap_211[7:0]) +
	( 13'sd 3660) * $signed(input_fmap_212[7:0]) +
	( 15'sd 14678) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23003) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5175) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28726) * $signed(input_fmap_216[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_217[7:0]) +
	( 16'sd 20831) * $signed(input_fmap_218[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22644) * $signed(input_fmap_220[7:0]) +
	( 16'sd 21811) * $signed(input_fmap_221[7:0]) +
	( 16'sd 30610) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25612) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27096) * $signed(input_fmap_224[7:0]) +
	( 15'sd 12450) * $signed(input_fmap_225[7:0]) +
	( 15'sd 8550) * $signed(input_fmap_226[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_227[7:0]) +
	( 16'sd 30228) * $signed(input_fmap_228[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_229[7:0]) +
	( 16'sd 19138) * $signed(input_fmap_230[7:0]) +
	( 16'sd 27157) * $signed(input_fmap_231[7:0]) +
	( 16'sd 31887) * $signed(input_fmap_232[7:0]) +
	( 15'sd 8740) * $signed(input_fmap_233[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_234[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_235[7:0]) +
	( 14'sd 6797) * $signed(input_fmap_236[7:0]) +
	( 16'sd 21801) * $signed(input_fmap_237[7:0]) +
	( 10'sd 353) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20066) * $signed(input_fmap_239[7:0]) +
	( 14'sd 5328) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23653) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5860) * $signed(input_fmap_242[7:0]) +
	( 16'sd 20459) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19809) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24229) * $signed(input_fmap_245[7:0]) +
	( 8'sd 80) * $signed(input_fmap_246[7:0]) +
	( 14'sd 7393) * $signed(input_fmap_247[7:0]) +
	( 15'sd 14561) * $signed(input_fmap_248[7:0]) +
	( 8'sd 125) * $signed(input_fmap_249[7:0]) +
	( 13'sd 2100) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4662) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13359) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5266) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2897) * $signed(input_fmap_254[7:0]) +
	( 16'sd 18977) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_76;
assign conv_mac_76 = 
	( 16'sd 31419) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10714) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9456) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10543) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16010) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28819) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8746) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17087) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5807) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23670) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19264) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5951) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2761) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1393) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5295) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26966) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22514) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28542) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28478) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5435) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1943) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8939) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7199) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10484) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4837) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15151) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13927) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27488) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2596) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2680) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28938) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25575) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4423) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21950) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15421) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22305) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1502) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19598) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29968) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9259) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15027) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28902) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32166) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28566) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29410) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31244) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24725) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22978) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5013) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20679) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29713) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19457) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18255) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22644) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3739) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32115) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22810) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24627) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6266) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31990) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10064) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28015) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18806) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28511) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31708) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12262) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20667) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25346) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17384) * $signed(input_fmap_77[7:0]) +
	( 14'sd 8058) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29042) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9451) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24796) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17413) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5406) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30778) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11126) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2809) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25481) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3456) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17061) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21196) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10558) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31958) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26434) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18680) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32747) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9458) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11931) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13577) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17446) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7404) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13412) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21162) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18279) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23180) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30397) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21012) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25085) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29585) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30237) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20694) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2948) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19240) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18877) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24621) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15542) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22612) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23596) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30525) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5536) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25944) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19402) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3150) * $signed(input_fmap_127[7:0]) +
	( 15'sd 14794) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31065) * $signed(input_fmap_130[7:0]) +
	( 14'sd 4621) * $signed(input_fmap_131[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28047) * $signed(input_fmap_133[7:0]) +
	( 16'sd 23111) * $signed(input_fmap_134[7:0]) +
	( 15'sd 9591) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13429) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13686) * $signed(input_fmap_137[7:0]) +
	( 14'sd 8013) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14692) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10926) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8975) * $signed(input_fmap_142[7:0]) +
	( 16'sd 24523) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11507) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17733) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27753) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19598) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6740) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_149[7:0]) +
	( 15'sd 12944) * $signed(input_fmap_150[7:0]) +
	( 16'sd 22014) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21194) * $signed(input_fmap_152[7:0]) +
	( 16'sd 26732) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10812) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10469) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17415) * $signed(input_fmap_156[7:0]) +
	( 14'sd 4109) * $signed(input_fmap_157[7:0]) +
	( 16'sd 26128) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5886) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24939) * $signed(input_fmap_160[7:0]) +
	( 16'sd 17163) * $signed(input_fmap_161[7:0]) +
	( 16'sd 25193) * $signed(input_fmap_162[7:0]) +
	( 9'sd 165) * $signed(input_fmap_163[7:0]) +
	( 16'sd 22916) * $signed(input_fmap_164[7:0]) +
	( 14'sd 7117) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2841) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23372) * $signed(input_fmap_167[7:0]) +
	( 16'sd 31491) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3713) * $signed(input_fmap_169[7:0]) +
	( 12'sd 2039) * $signed(input_fmap_170[7:0]) +
	( 16'sd 27061) * $signed(input_fmap_171[7:0]) +
	( 16'sd 32047) * $signed(input_fmap_172[7:0]) +
	( 16'sd 32762) * $signed(input_fmap_173[7:0]) +
	( 16'sd 17300) * $signed(input_fmap_174[7:0]) +
	( 15'sd 12923) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27479) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20924) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4622) * $signed(input_fmap_180[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_181[7:0]) +
	( 16'sd 18135) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17676) * $signed(input_fmap_183[7:0]) +
	( 16'sd 19610) * $signed(input_fmap_184[7:0]) +
	( 15'sd 13352) * $signed(input_fmap_185[7:0]) +
	( 15'sd 11665) * $signed(input_fmap_186[7:0]) +
	( 16'sd 24866) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23316) * $signed(input_fmap_188[7:0]) +
	( 15'sd 10868) * $signed(input_fmap_189[7:0]) +
	( 15'sd 16121) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17636) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14189) * $signed(input_fmap_192[7:0]) +
	( 14'sd 4108) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12615) * $signed(input_fmap_194[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25557) * $signed(input_fmap_196[7:0]) +
	( 16'sd 29723) * $signed(input_fmap_197[7:0]) +
	( 15'sd 12220) * $signed(input_fmap_198[7:0]) +
	( 15'sd 13562) * $signed(input_fmap_199[7:0]) +
	( 10'sd 426) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18510) * $signed(input_fmap_201[7:0]) +
	( 16'sd 26357) * $signed(input_fmap_202[7:0]) +
	( 15'sd 8523) * $signed(input_fmap_203[7:0]) +
	( 16'sd 27548) * $signed(input_fmap_204[7:0]) +
	( 16'sd 17638) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3028) * $signed(input_fmap_206[7:0]) +
	( 11'sd 738) * $signed(input_fmap_207[7:0]) +
	( 16'sd 24063) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20303) * $signed(input_fmap_209[7:0]) +
	( 16'sd 17706) * $signed(input_fmap_210[7:0]) +
	( 16'sd 25205) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26869) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24784) * $signed(input_fmap_213[7:0]) +
	( 14'sd 5642) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6543) * $signed(input_fmap_215[7:0]) +
	( 16'sd 30438) * $signed(input_fmap_216[7:0]) +
	( 12'sd 1667) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7413) * $signed(input_fmap_218[7:0]) +
	( 14'sd 4553) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19082) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_221[7:0]) +
	( 16'sd 24734) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1878) * $signed(input_fmap_224[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_225[7:0]) +
	( 15'sd 15945) * $signed(input_fmap_226[7:0]) +
	( 14'sd 4797) * $signed(input_fmap_227[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6146) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29931) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13465) * $signed(input_fmap_231[7:0]) +
	( 16'sd 31063) * $signed(input_fmap_232[7:0]) +
	( 15'sd 8899) * $signed(input_fmap_233[7:0]) +
	( 11'sd 824) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14192) * $signed(input_fmap_235[7:0]) +
	( 16'sd 22675) * $signed(input_fmap_236[7:0]) +
	( 15'sd 12472) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3356) * $signed(input_fmap_238[7:0]) +
	( 13'sd 3105) * $signed(input_fmap_239[7:0]) +
	( 16'sd 32423) * $signed(input_fmap_240[7:0]) +
	( 12'sd 1333) * $signed(input_fmap_241[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23610) * $signed(input_fmap_243[7:0]) +
	( 13'sd 3426) * $signed(input_fmap_244[7:0]) +
	( 10'sd 463) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_246[7:0]) +
	( 16'sd 29363) * $signed(input_fmap_247[7:0]) +
	( 15'sd 15783) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4232) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7732) * $signed(input_fmap_250[7:0]) +
	( 15'sd 8370) * $signed(input_fmap_251[7:0]) +
	( 16'sd 32556) * $signed(input_fmap_252[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_253[7:0]) +
	( 15'sd 15751) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5109) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_77;
assign conv_mac_77 = 
	( 13'sd 3091) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19235) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16206) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9360) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3295) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20876) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11914) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16714) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9514) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3965) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4799) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18265) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21980) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9204) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27725) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12111) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2869) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5832) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9588) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26177) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24326) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27021) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32752) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28608) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26034) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14317) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12861) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23930) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17687) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22724) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15613) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31598) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15969) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31981) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15692) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1905) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11464) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21996) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15356) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29561) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10729) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11286) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9169) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8092) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22971) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24770) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5874) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32567) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6386) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29925) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17183) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6796) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31998) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14093) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13510) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32661) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21835) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30778) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26506) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28851) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32575) * $signed(input_fmap_67[7:0]) +
	( 13'sd 4003) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27452) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29235) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26644) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11267) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5920) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23403) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30932) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1511) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2898) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17298) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17816) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24898) * $signed(input_fmap_80[7:0]) +
	( 11'sd 1000) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3255) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13263) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5506) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1042) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25359) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12627) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29005) * $signed(input_fmap_89[7:0]) +
	( 10'sd 387) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27834) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25787) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30577) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13470) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4105) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7426) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10694) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25640) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8644) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25780) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2740) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10012) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17513) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18451) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7632) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18093) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13477) * $signed(input_fmap_107[7:0]) +
	( 11'sd 532) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5712) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8647) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1488) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6086) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10342) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23354) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21739) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17359) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18883) * $signed(input_fmap_118[7:0]) +
	( 13'sd 4065) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12476) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17188) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27300) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10578) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13588) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20411) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27476) * $signed(input_fmap_127[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_128[7:0]) +
	( 16'sd 22473) * $signed(input_fmap_129[7:0]) +
	( 14'sd 4998) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5189) * $signed(input_fmap_131[7:0]) +
	( 13'sd 2808) * $signed(input_fmap_132[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3915) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32558) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25903) * $signed(input_fmap_136[7:0]) +
	( 16'sd 28323) * $signed(input_fmap_137[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24941) * $signed(input_fmap_139[7:0]) +
	( 16'sd 23370) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18517) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31153) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11790) * $signed(input_fmap_144[7:0]) +
	( 12'sd 1561) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7544) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14806) * $signed(input_fmap_147[7:0]) +
	( 10'sd 316) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18852) * $signed(input_fmap_149[7:0]) +
	( 14'sd 4349) * $signed(input_fmap_150[7:0]) +
	( 16'sd 22141) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30144) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27633) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23334) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22990) * $signed(input_fmap_155[7:0]) +
	( 16'sd 26153) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6749) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11607) * $signed(input_fmap_158[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_159[7:0]) +
	( 14'sd 7616) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31376) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30667) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22397) * $signed(input_fmap_163[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14516) * $signed(input_fmap_165[7:0]) +
	( 16'sd 28376) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9069) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14550) * $signed(input_fmap_168[7:0]) +
	( 16'sd 19486) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23656) * $signed(input_fmap_170[7:0]) +
	( 12'sd 1429) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5587) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7827) * $signed(input_fmap_174[7:0]) +
	( 13'sd 2277) * $signed(input_fmap_175[7:0]) +
	( 16'sd 22580) * $signed(input_fmap_176[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_177[7:0]) +
	( 13'sd 3826) * $signed(input_fmap_178[7:0]) +
	( 15'sd 10673) * $signed(input_fmap_179[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25468) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10833) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5340) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31241) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25468) * $signed(input_fmap_185[7:0]) +
	( 16'sd 32517) * $signed(input_fmap_186[7:0]) +
	( 14'sd 6988) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12030) * $signed(input_fmap_188[7:0]) +
	( 15'sd 15916) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_191[7:0]) +
	( 15'sd 9105) * $signed(input_fmap_192[7:0]) +
	( 16'sd 31828) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14677) * $signed(input_fmap_195[7:0]) +
	( 16'sd 26833) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1925) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5091) * $signed(input_fmap_198[7:0]) +
	( 16'sd 25388) * $signed(input_fmap_199[7:0]) +
	( 15'sd 11152) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3226) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2551) * $signed(input_fmap_202[7:0]) +
	( 15'sd 10279) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12313) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18503) * $signed(input_fmap_205[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_206[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30615) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_209[7:0]) +
	( 15'sd 13109) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17137) * $signed(input_fmap_211[7:0]) +
	( 16'sd 31997) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2592) * $signed(input_fmap_213[7:0]) +
	( 11'sd 766) * $signed(input_fmap_214[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_215[7:0]) +
	( 16'sd 16402) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24254) * $signed(input_fmap_217[7:0]) +
	( 15'sd 12133) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19951) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14461) * $signed(input_fmap_220[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14974) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_223[7:0]) +
	( 15'sd 15059) * $signed(input_fmap_224[7:0]) +
	( 15'sd 9347) * $signed(input_fmap_225[7:0]) +
	( 12'sd 1667) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20599) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31301) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_229[7:0]) +
	( 15'sd 8390) * $signed(input_fmap_230[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_231[7:0]) +
	( 14'sd 4956) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10190) * $signed(input_fmap_233[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5543) * $signed(input_fmap_235[7:0]) +
	( 16'sd 19686) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28278) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13766) * $signed(input_fmap_238[7:0]) +
	( 16'sd 25595) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3647) * $signed(input_fmap_241[7:0]) +
	( 16'sd 32718) * $signed(input_fmap_242[7:0]) +
	( 12'sd 1836) * $signed(input_fmap_243[7:0]) +
	( 16'sd 27435) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28767) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19166) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20104) * $signed(input_fmap_247[7:0]) +
	( 14'sd 7204) * $signed(input_fmap_248[7:0]) +
	( 12'sd 1959) * $signed(input_fmap_249[7:0]) +
	( 16'sd 18946) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7967) * $signed(input_fmap_251[7:0]) +
	( 11'sd 904) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19258) * $signed(input_fmap_254[7:0]) +
	( 14'sd 6260) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_78;
assign conv_mac_78 = 
	( 16'sd 31077) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9786) * $signed(input_fmap_1[7:0]) +
	( 14'sd 8138) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3612) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27781) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24219) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18401) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13113) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28497) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24505) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17462) * $signed(input_fmap_14[7:0]) +
	( 11'sd 987) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27302) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10339) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30143) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14575) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24385) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25148) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20322) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5238) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30771) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1289) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_27[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15999) * $signed(input_fmap_29[7:0]) +
	( 8'sd 76) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20585) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24627) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22863) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30960) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21572) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6430) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8930) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18367) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22641) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23808) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1188) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4731) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21991) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17613) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25251) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19619) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8317) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29197) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7234) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_52[7:0]) +
	( 10'sd 454) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7581) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19086) * $signed(input_fmap_55[7:0]) +
	( 13'sd 4064) * $signed(input_fmap_56[7:0]) +
	( 16'sd 16826) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4212) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10833) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23816) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19517) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18974) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12657) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27085) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14012) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27005) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15891) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8420) * $signed(input_fmap_69[7:0]) +
	( 16'sd 26030) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31983) * $signed(input_fmap_71[7:0]) +
	( 11'sd 973) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28047) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6728) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12390) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20437) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6334) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8182) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20519) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3516) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14237) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2067) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3341) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14607) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29759) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9153) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9111) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25261) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11783) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8718) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22215) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6280) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15662) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8318) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23790) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2502) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19222) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29312) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23444) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19312) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18685) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19399) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19485) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17854) * $signed(input_fmap_109[7:0]) +
	( 10'sd 358) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15743) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32437) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25522) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22801) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19279) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10344) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3888) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16618) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14773) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9686) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19272) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26104) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26477) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32128) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29223) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25955) * $signed(input_fmap_127[7:0]) +
	( 16'sd 32382) * $signed(input_fmap_128[7:0]) +
	( 16'sd 20589) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30702) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20889) * $signed(input_fmap_131[7:0]) +
	( 15'sd 12828) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10852) * $signed(input_fmap_133[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31734) * $signed(input_fmap_135[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27659) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31594) * $signed(input_fmap_138[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_140[7:0]) +
	( 16'sd 26975) * $signed(input_fmap_141[7:0]) +
	( 16'sd 23364) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_143[7:0]) +
	( 16'sd 29886) * $signed(input_fmap_144[7:0]) +
	( 14'sd 4577) * $signed(input_fmap_145[7:0]) +
	( 15'sd 13133) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11249) * $signed(input_fmap_147[7:0]) +
	( 16'sd 18887) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18341) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21157) * $signed(input_fmap_150[7:0]) +
	( 15'sd 8244) * $signed(input_fmap_151[7:0]) +
	( 13'sd 3515) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31855) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22805) * $signed(input_fmap_154[7:0]) +
	( 15'sd 11438) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_156[7:0]) +
	( 13'sd 2149) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28617) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4530) * $signed(input_fmap_159[7:0]) +
	( 16'sd 23988) * $signed(input_fmap_160[7:0]) +
	( 16'sd 16825) * $signed(input_fmap_161[7:0]) +
	( 15'sd 8407) * $signed(input_fmap_162[7:0]) +
	( 16'sd 25664) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6935) * $signed(input_fmap_164[7:0]) +
	( 16'sd 17653) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30975) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30023) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5922) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3395) * $signed(input_fmap_169[7:0]) +
	( 14'sd 6615) * $signed(input_fmap_170[7:0]) +
	( 16'sd 17377) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3318) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19895) * $signed(input_fmap_173[7:0]) +
	( 16'sd 24821) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7331) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_176[7:0]) +
	( 14'sd 8034) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1105) * $signed(input_fmap_178[7:0]) +
	( 15'sd 9429) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4714) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25448) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29248) * $signed(input_fmap_182[7:0]) +
	( 14'sd 4373) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14845) * $signed(input_fmap_184[7:0]) +
	( 16'sd 28695) * $signed(input_fmap_185[7:0]) +
	( 16'sd 27362) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_187[7:0]) +
	( 15'sd 15508) * $signed(input_fmap_188[7:0]) +
	( 16'sd 23411) * $signed(input_fmap_189[7:0]) +
	( 16'sd 24317) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19544) * $signed(input_fmap_192[7:0]) +
	( 16'sd 32272) * $signed(input_fmap_193[7:0]) +
	( 16'sd 28503) * $signed(input_fmap_194[7:0]) +
	( 15'sd 10884) * $signed(input_fmap_195[7:0]) +
	( 16'sd 16598) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11334) * $signed(input_fmap_197[7:0]) +
	( 15'sd 11795) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20796) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5836) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11019) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21679) * $signed(input_fmap_202[7:0]) +
	( 16'sd 28704) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_204[7:0]) +
	( 16'sd 26412) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6718) * $signed(input_fmap_206[7:0]) +
	( 16'sd 31732) * $signed(input_fmap_207[7:0]) +
	( 15'sd 16111) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14824) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15242) * $signed(input_fmap_211[7:0]) +
	( 13'sd 2269) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3468) * $signed(input_fmap_213[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_214[7:0]) +
	( 16'sd 27455) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28076) * $signed(input_fmap_216[7:0]) +
	( 11'sd 719) * $signed(input_fmap_217[7:0]) +
	( 16'sd 17978) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17560) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24468) * $signed(input_fmap_220[7:0]) +
	( 14'sd 7355) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2938) * $signed(input_fmap_222[7:0]) +
	( 16'sd 29815) * $signed(input_fmap_223[7:0]) +
	( 13'sd 2569) * $signed(input_fmap_224[7:0]) +
	( 16'sd 25955) * $signed(input_fmap_225[7:0]) +
	( 16'sd 26484) * $signed(input_fmap_226[7:0]) +
	( 15'sd 16362) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24665) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8677) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18651) * $signed(input_fmap_230[7:0]) +
	( 16'sd 23111) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7074) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14387) * $signed(input_fmap_233[7:0]) +
	( 16'sd 16943) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29587) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14726) * $signed(input_fmap_237[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_238[7:0]) +
	( 15'sd 15037) * $signed(input_fmap_239[7:0]) +
	( 14'sd 4974) * $signed(input_fmap_240[7:0]) +
	( 15'sd 11911) * $signed(input_fmap_241[7:0]) +
	( 15'sd 9777) * $signed(input_fmap_242[7:0]) +
	( 16'sd 24539) * $signed(input_fmap_243[7:0]) +
	( 16'sd 26609) * $signed(input_fmap_244[7:0]) +
	( 16'sd 32150) * $signed(input_fmap_245[7:0]) +
	( 16'sd 24443) * $signed(input_fmap_246[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1967) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15582) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_250[7:0]) +
	( 13'sd 3524) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30988) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11277) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10324) * $signed(input_fmap_254[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_79;
assign conv_mac_79 = 
	( 15'sd 15878) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16009) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15053) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12232) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31977) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22894) * $signed(input_fmap_7[7:0]) +
	( 11'sd 776) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28047) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31430) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10987) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9195) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9053) * $signed(input_fmap_16[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29050) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9983) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28021) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26020) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23907) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20245) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14124) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32595) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7825) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32226) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24709) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3168) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29761) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31487) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30878) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4301) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24243) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23167) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14840) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10477) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4177) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19964) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20196) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29372) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20689) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4380) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9433) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32350) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7746) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9282) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1366) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16918) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9345) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26940) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28990) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15392) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25140) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15047) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11533) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17438) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3346) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22748) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9257) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5303) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20546) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3815) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29589) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23532) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9613) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22555) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1744) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3983) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3085) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2140) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20625) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16598) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26464) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14941) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18375) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15779) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22284) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25703) * $signed(input_fmap_94[7:0]) +
	( 12'sd 2036) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1989) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14870) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6804) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25843) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13609) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30143) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11751) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28903) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14526) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3931) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24067) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23304) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2869) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9006) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30389) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21928) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24701) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11101) * $signed(input_fmap_115[7:0]) +
	( 11'sd 560) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22878) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19929) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8920) * $signed(input_fmap_119[7:0]) +
	( 10'sd 448) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15148) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7434) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17334) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24724) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13524) * $signed(input_fmap_126[7:0]) +
	( 15'sd 16001) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4506) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30424) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13337) * $signed(input_fmap_131[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_132[7:0]) +
	( 15'sd 14618) * $signed(input_fmap_133[7:0]) +
	( 16'sd 20331) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31793) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4577) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27491) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11052) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24608) * $signed(input_fmap_139[7:0]) +
	( 15'sd 13543) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20587) * $signed(input_fmap_141[7:0]) +
	( 15'sd 15607) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17105) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22153) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2260) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1609) * $signed(input_fmap_146[7:0]) +
	( 16'sd 20688) * $signed(input_fmap_147[7:0]) +
	( 15'sd 10656) * $signed(input_fmap_148[7:0]) +
	( 15'sd 8520) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23288) * $signed(input_fmap_150[7:0]) +
	( 16'sd 22479) * $signed(input_fmap_151[7:0]) +
	( 11'sd 750) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1871) * $signed(input_fmap_153[7:0]) +
	( 16'sd 19497) * $signed(input_fmap_154[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_155[7:0]) +
	( 15'sd 11816) * $signed(input_fmap_156[7:0]) +
	( 9'sd 232) * $signed(input_fmap_157[7:0]) +
	( 11'sd 599) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3687) * $signed(input_fmap_159[7:0]) +
	( 16'sd 23305) * $signed(input_fmap_160[7:0]) +
	( 16'sd 27089) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21120) * $signed(input_fmap_162[7:0]) +
	( 15'sd 14414) * $signed(input_fmap_163[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_164[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_165[7:0]) +
	( 16'sd 25307) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9742) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12441) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9621) * $signed(input_fmap_170[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12996) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1711) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32201) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29784) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2156) * $signed(input_fmap_177[7:0]) +
	( 16'sd 25032) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6790) * $signed(input_fmap_180[7:0]) +
	( 15'sd 13937) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26193) * $signed(input_fmap_182[7:0]) +
	( 16'sd 26782) * $signed(input_fmap_183[7:0]) +
	( 16'sd 20019) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22486) * $signed(input_fmap_185[7:0]) +
	( 12'sd 1423) * $signed(input_fmap_186[7:0]) +
	( 16'sd 23021) * $signed(input_fmap_187[7:0]) +
	( 16'sd 30141) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11820) * $signed(input_fmap_189[7:0]) +
	( 15'sd 11002) * $signed(input_fmap_190[7:0]) +
	( 16'sd 30877) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_192[7:0]) +
	( 11'sd 554) * $signed(input_fmap_193[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_194[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20930) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32548) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22383) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20476) * $signed(input_fmap_199[7:0]) +
	( 6'sd 25) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15064) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19458) * $signed(input_fmap_202[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32701) * $signed(input_fmap_204[7:0]) +
	( 15'sd 14552) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28453) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1932) * $signed(input_fmap_207[7:0]) +
	( 16'sd 23198) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26724) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3992) * $signed(input_fmap_210[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_211[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_212[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14880) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10626) * $signed(input_fmap_215[7:0]) +
	( 13'sd 4038) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_217[7:0]) +
	( 16'sd 19067) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14584) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4782) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25450) * $signed(input_fmap_221[7:0]) +
	( 16'sd 31295) * $signed(input_fmap_222[7:0]) +
	( 16'sd 20812) * $signed(input_fmap_223[7:0]) +
	( 16'sd 29266) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18774) * $signed(input_fmap_225[7:0]) +
	( 16'sd 21875) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3654) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_228[7:0]) +
	( 16'sd 18787) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15808) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17008) * $signed(input_fmap_231[7:0]) +
	( 16'sd 32385) * $signed(input_fmap_232[7:0]) +
	( 14'sd 6854) * $signed(input_fmap_233[7:0]) +
	( 16'sd 20228) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26803) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14878) * $signed(input_fmap_237[7:0]) +
	( 14'sd 6722) * $signed(input_fmap_238[7:0]) +
	( 13'sd 3292) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31221) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30064) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23381) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22328) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22050) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12473) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30458) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3188) * $signed(input_fmap_247[7:0]) +
	( 16'sd 23618) * $signed(input_fmap_248[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_250[7:0]) +
	( 16'sd 28314) * $signed(input_fmap_251[7:0]) +
	( 16'sd 31665) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13514) * $signed(input_fmap_253[7:0]) +
	( 11'sd 636) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_80;
assign conv_mac_80 = 
	( 14'sd 8134) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21229) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22217) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13346) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31180) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9512) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2645) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21191) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20269) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10101) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6251) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30088) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17695) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31519) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12967) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32575) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28632) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4697) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26662) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14825) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4512) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31465) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12073) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22425) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18577) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29566) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10289) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5411) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17016) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21903) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25582) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20547) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18220) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22491) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19476) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21704) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29415) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18967) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13522) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32682) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21700) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1301) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17885) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25841) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24590) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2634) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20440) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11516) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1669) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2289) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2451) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16433) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27971) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24001) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4324) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17092) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1856) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2199) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26818) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18538) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32087) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22874) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24016) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29358) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13333) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17199) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7791) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19003) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25395) * $signed(input_fmap_73[7:0]) +
	( 12'sd 1993) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32314) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18554) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7346) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13313) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14004) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1368) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8507) * $signed(input_fmap_84[7:0]) +
	( 10'sd 297) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17561) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14227) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8689) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12606) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4803) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21998) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19091) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15574) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11333) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6397) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15329) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31005) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22543) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24746) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6743) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4273) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20527) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31540) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19384) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7001) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28638) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1265) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9599) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7788) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15418) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29750) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22356) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13845) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5372) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19123) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15827) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19379) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28187) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13473) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1529) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24111) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19946) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5173) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_128[7:0]) +
	( 16'sd 30668) * $signed(input_fmap_129[7:0]) +
	( 14'sd 4445) * $signed(input_fmap_130[7:0]) +
	( 12'sd 1684) * $signed(input_fmap_131[7:0]) +
	( 16'sd 26529) * $signed(input_fmap_132[7:0]) +
	( 15'sd 16047) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24234) * $signed(input_fmap_134[7:0]) +
	( 14'sd 6137) * $signed(input_fmap_135[7:0]) +
	( 16'sd 28928) * $signed(input_fmap_136[7:0]) +
	( 16'sd 28566) * $signed(input_fmap_137[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31566) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30589) * $signed(input_fmap_140[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27227) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_143[7:0]) +
	( 16'sd 16710) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17845) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3724) * $signed(input_fmap_146[7:0]) +
	( 14'sd 4755) * $signed(input_fmap_147[7:0]) +
	( 16'sd 18159) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25571) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27076) * $signed(input_fmap_150[7:0]) +
	( 14'sd 7290) * $signed(input_fmap_151[7:0]) +
	( 15'sd 16130) * $signed(input_fmap_152[7:0]) +
	( 11'sd 569) * $signed(input_fmap_153[7:0]) +
	( 14'sd 5938) * $signed(input_fmap_154[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_156[7:0]) +
	( 16'sd 28502) * $signed(input_fmap_157[7:0]) +
	( 14'sd 5667) * $signed(input_fmap_158[7:0]) +
	( 16'sd 25235) * $signed(input_fmap_159[7:0]) +
	( 13'sd 2092) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1716) * $signed(input_fmap_161[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_162[7:0]) +
	( 16'sd 19820) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10562) * $signed(input_fmap_164[7:0]) +
	( 16'sd 31350) * $signed(input_fmap_165[7:0]) +
	( 15'sd 15745) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26655) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6884) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18992) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16687) * $signed(input_fmap_171[7:0]) +
	( 7'sd 38) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5830) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32190) * $signed(input_fmap_174[7:0]) +
	( 15'sd 12284) * $signed(input_fmap_175[7:0]) +
	( 12'sd 2003) * $signed(input_fmap_176[7:0]) +
	( 16'sd 25241) * $signed(input_fmap_177[7:0]) +
	( 16'sd 21957) * $signed(input_fmap_178[7:0]) +
	( 15'sd 14304) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_180[7:0]) +
	( 15'sd 12851) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26441) * $signed(input_fmap_182[7:0]) +
	( 15'sd 15099) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15494) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9272) * $signed(input_fmap_187[7:0]) +
	( 16'sd 28067) * $signed(input_fmap_188[7:0]) +
	( 16'sd 18779) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28135) * $signed(input_fmap_190[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19774) * $signed(input_fmap_192[7:0]) +
	( 13'sd 3430) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3640) * $signed(input_fmap_194[7:0]) +
	( 16'sd 28307) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22041) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19043) * $signed(input_fmap_197[7:0]) +
	( 14'sd 7851) * $signed(input_fmap_198[7:0]) +
	( 15'sd 11347) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25822) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22834) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18086) * $signed(input_fmap_202[7:0]) +
	( 15'sd 10833) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1080) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12947) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28138) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25844) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_210[7:0]) +
	( 14'sd 8149) * $signed(input_fmap_211[7:0]) +
	( 15'sd 9034) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2812) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17729) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11630) * $signed(input_fmap_215[7:0]) +
	( 16'sd 27695) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17639) * $signed(input_fmap_217[7:0]) +
	( 14'sd 4265) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21645) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1682) * $signed(input_fmap_220[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14889) * $signed(input_fmap_222[7:0]) +
	( 14'sd 4252) * $signed(input_fmap_223[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_224[7:0]) +
	( 15'sd 11163) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6898) * $signed(input_fmap_226[7:0]) +
	( 14'sd 4948) * $signed(input_fmap_227[7:0]) +
	( 14'sd 6916) * $signed(input_fmap_228[7:0]) +
	( 16'sd 21306) * $signed(input_fmap_229[7:0]) +
	( 15'sd 10152) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28043) * $signed(input_fmap_231[7:0]) +
	( 16'sd 19326) * $signed(input_fmap_232[7:0]) +
	( 16'sd 20144) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_234[7:0]) +
	( 15'sd 15226) * $signed(input_fmap_235[7:0]) +
	( 16'sd 16933) * $signed(input_fmap_236[7:0]) +
	( 15'sd 12068) * $signed(input_fmap_237[7:0]) +
	( 16'sd 30774) * $signed(input_fmap_238[7:0]) +
	( 16'sd 28699) * $signed(input_fmap_239[7:0]) +
	( 15'sd 15994) * $signed(input_fmap_240[7:0]) +
	( 15'sd 12578) * $signed(input_fmap_241[7:0]) +
	( 16'sd 24886) * $signed(input_fmap_242[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_243[7:0]) +
	( 16'sd 17100) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6857) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9627) * $signed(input_fmap_246[7:0]) +
	( 16'sd 31998) * $signed(input_fmap_247[7:0]) +
	( 15'sd 16325) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15048) * $signed(input_fmap_249[7:0]) +
	( 14'sd 4931) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21786) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12368) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25717) * $signed(input_fmap_253[7:0]) +
	( 16'sd 24872) * $signed(input_fmap_254[7:0]) +
	( 11'sd 973) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_81;
assign conv_mac_81 = 
	( 16'sd 21929) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13466) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1731) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27096) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18859) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25997) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28490) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2302) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7109) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26908) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18024) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12057) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16628) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17077) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22300) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21917) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24296) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17510) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20191) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19779) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22650) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27020) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3923) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26728) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16597) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31040) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19004) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29522) * $signed(input_fmap_30[7:0]) +
	( 11'sd 885) * $signed(input_fmap_31[7:0]) +
	( 6'sd 16) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30765) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17547) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14195) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19348) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8633) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28834) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1809) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12974) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2995) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25460) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28903) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7107) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27659) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5867) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10244) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14728) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3688) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25716) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8479) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24894) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4907) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15735) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31848) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4805) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23388) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13343) * $signed(input_fmap_61[7:0]) +
	( 11'sd 966) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5637) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9819) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23849) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15960) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14103) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11642) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15646) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17869) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18942) * $signed(input_fmap_71[7:0]) +
	( 15'sd 9397) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9762) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21660) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8206) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4298) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_78[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17392) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25899) * $signed(input_fmap_81[7:0]) +
	( 15'sd 16056) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16505) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10570) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11321) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24952) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22555) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8841) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9155) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12895) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28088) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29981) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23564) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1142) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8419) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31763) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29938) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12246) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26115) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18169) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6222) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22691) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19481) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27690) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13683) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26378) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6304) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26767) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31167) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28725) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12075) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26242) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25544) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30387) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25145) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20131) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21513) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31631) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28375) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27654) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16390) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21450) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30290) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12244) * $signed(input_fmap_126[7:0]) +
	( 11'sd 958) * $signed(input_fmap_127[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7892) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25014) * $signed(input_fmap_130[7:0]) +
	( 14'sd 4759) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14823) * $signed(input_fmap_132[7:0]) +
	( 11'sd 579) * $signed(input_fmap_133[7:0]) +
	( 16'sd 23398) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26936) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13735) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12628) * $signed(input_fmap_137[7:0]) +
	( 16'sd 26434) * $signed(input_fmap_138[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_140[7:0]) +
	( 10'sd 310) * $signed(input_fmap_141[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4705) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18734) * $signed(input_fmap_144[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_145[7:0]) +
	( 16'sd 31982) * $signed(input_fmap_146[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_148[7:0]) +
	( 16'sd 22099) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27530) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24848) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7856) * $signed(input_fmap_152[7:0]) +
	( 11'sd 762) * $signed(input_fmap_153[7:0]) +
	( 16'sd 20289) * $signed(input_fmap_154[7:0]) +
	( 14'sd 4348) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_156[7:0]) +
	( 15'sd 9165) * $signed(input_fmap_157[7:0]) +
	( 15'sd 12428) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26265) * $signed(input_fmap_159[7:0]) +
	( 7'sd 37) * $signed(input_fmap_160[7:0]) +
	( 15'sd 14639) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10490) * $signed(input_fmap_162[7:0]) +
	( 16'sd 17873) * $signed(input_fmap_163[7:0]) +
	( 16'sd 17328) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_165[7:0]) +
	( 14'sd 7354) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17984) * $signed(input_fmap_167[7:0]) +
	( 16'sd 23582) * $signed(input_fmap_168[7:0]) +
	( 12'sd 1637) * $signed(input_fmap_169[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20453) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4997) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27318) * $signed(input_fmap_173[7:0]) +
	( 12'sd 1393) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15014) * $signed(input_fmap_175[7:0]) +
	( 16'sd 30290) * $signed(input_fmap_176[7:0]) +
	( 16'sd 26313) * $signed(input_fmap_177[7:0]) +
	( 14'sd 6778) * $signed(input_fmap_178[7:0]) +
	( 16'sd 23341) * $signed(input_fmap_179[7:0]) +
	( 16'sd 20854) * $signed(input_fmap_180[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_181[7:0]) +
	( 16'sd 28957) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_184[7:0]) +
	( 14'sd 4281) * $signed(input_fmap_185[7:0]) +
	( 15'sd 10809) * $signed(input_fmap_186[7:0]) +
	( 15'sd 8921) * $signed(input_fmap_187[7:0]) +
	( 16'sd 27224) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17856) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32069) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12440) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6533) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21205) * $signed(input_fmap_194[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_195[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_197[7:0]) +
	( 13'sd 3842) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20805) * $signed(input_fmap_199[7:0]) +
	( 13'sd 2859) * $signed(input_fmap_200[7:0]) +
	( 16'sd 29798) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11388) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6999) * $signed(input_fmap_203[7:0]) +
	( 13'sd 3079) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28539) * $signed(input_fmap_205[7:0]) +
	( 10'sd 453) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7503) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11485) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26374) * $signed(input_fmap_209[7:0]) +
	( 16'sd 22573) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5326) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14617) * $signed(input_fmap_212[7:0]) +
	( 16'sd 31461) * $signed(input_fmap_213[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_214[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_216[7:0]) +
	( 12'sd 1300) * $signed(input_fmap_217[7:0]) +
	( 14'sd 4459) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10828) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22761) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12940) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25977) * $signed(input_fmap_222[7:0]) +
	( 16'sd 31208) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27029) * $signed(input_fmap_224[7:0]) +
	( 16'sd 24056) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18806) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6738) * $signed(input_fmap_227[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10128) * $signed(input_fmap_229[7:0]) +
	( 15'sd 12083) * $signed(input_fmap_230[7:0]) +
	( 14'sd 5612) * $signed(input_fmap_231[7:0]) +
	( 16'sd 31862) * $signed(input_fmap_232[7:0]) +
	( 10'sd 345) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5684) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12841) * $signed(input_fmap_236[7:0]) +
	( 16'sd 25893) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13971) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23707) * $signed(input_fmap_239[7:0]) +
	( 14'sd 5998) * $signed(input_fmap_240[7:0]) +
	( 15'sd 9074) * $signed(input_fmap_241[7:0]) +
	( 13'sd 4033) * $signed(input_fmap_242[7:0]) +
	( 16'sd 32748) * $signed(input_fmap_243[7:0]) +
	( 16'sd 27486) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3335) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31025) * $signed(input_fmap_246[7:0]) +
	( 16'sd 25502) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13293) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30697) * $signed(input_fmap_249[7:0]) +
	( 14'sd 6619) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28510) * $signed(input_fmap_252[7:0]) +
	( 16'sd 20833) * $signed(input_fmap_253[7:0]) +
	( 16'sd 24109) * $signed(input_fmap_254[7:0]) +
	( 16'sd 27828) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_82;
assign conv_mac_82 = 
	( 16'sd 16473) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31653) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24542) * $signed(input_fmap_2[7:0]) +
	( 10'sd 488) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19306) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11049) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17472) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16741) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17221) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2918) * $signed(input_fmap_9[7:0]) +
	( 15'sd 11461) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7639) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21815) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21073) * $signed(input_fmap_14[7:0]) +
	( 16'sd 19734) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27022) * $signed(input_fmap_16[7:0]) +
	( 12'sd 2017) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4469) * $signed(input_fmap_18[7:0]) +
	( 15'sd 16013) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32016) * $signed(input_fmap_20[7:0]) +
	( 10'sd 334) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21881) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23455) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2073) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10457) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2951) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21555) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17262) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11928) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28555) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27257) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10844) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9902) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9248) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4679) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7231) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7653) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11691) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29986) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10069) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3034) * $signed(input_fmap_44[7:0]) +
	( 7'sd 40) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32122) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31850) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4895) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27492) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15180) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28250) * $signed(input_fmap_52[7:0]) +
	( 14'sd 8132) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29474) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18986) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13077) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9683) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13481) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29512) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30800) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29108) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11113) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2125) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12871) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18315) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5069) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4608) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6627) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31887) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21153) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14808) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14844) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17016) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19245) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18806) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27936) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27117) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18377) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9389) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18539) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26677) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24120) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6242) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19464) * $signed(input_fmap_87[7:0]) +
	( 11'sd 989) * $signed(input_fmap_88[7:0]) +
	( 9'sd 128) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6532) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28103) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_94[7:0]) +
	( 10'sd 463) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21617) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13504) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7973) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31264) * $signed(input_fmap_101[7:0]) +
	( 12'sd 2036) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13392) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2601) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15686) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16668) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8501) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20818) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23457) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14657) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31938) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11617) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3832) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27573) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6259) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22444) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2580) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13799) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22390) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13698) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28068) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16843) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11547) * $signed(input_fmap_127[7:0]) +
	( 14'sd 6659) * $signed(input_fmap_128[7:0]) +
	( 15'sd 16223) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10531) * $signed(input_fmap_130[7:0]) +
	( 14'sd 6299) * $signed(input_fmap_131[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28801) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24576) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31888) * $signed(input_fmap_135[7:0]) +
	( 14'sd 8040) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_137[7:0]) +
	( 15'sd 12783) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_139[7:0]) +
	( 15'sd 14421) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12863) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22932) * $signed(input_fmap_142[7:0]) +
	( 16'sd 22991) * $signed(input_fmap_143[7:0]) +
	( 15'sd 15999) * $signed(input_fmap_144[7:0]) +
	( 15'sd 10365) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15374) * $signed(input_fmap_146[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_147[7:0]) +
	( 16'sd 27036) * $signed(input_fmap_148[7:0]) +
	( 16'sd 31502) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18279) * $signed(input_fmap_150[7:0]) +
	( 14'sd 5358) * $signed(input_fmap_151[7:0]) +
	( 12'sd 1204) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3041) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23837) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5326) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29806) * $signed(input_fmap_156[7:0]) +
	( 15'sd 12159) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18187) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6062) * $signed(input_fmap_159[7:0]) +
	( 12'sd 1799) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22564) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24776) * $signed(input_fmap_162[7:0]) +
	( 12'sd 1906) * $signed(input_fmap_163[7:0]) +
	( 8'sd 115) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4195) * $signed(input_fmap_165[7:0]) +
	( 15'sd 15909) * $signed(input_fmap_166[7:0]) +
	( 15'sd 10203) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29241) * $signed(input_fmap_168[7:0]) +
	( 15'sd 9419) * $signed(input_fmap_169[7:0]) +
	( 15'sd 16360) * $signed(input_fmap_170[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11571) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27004) * $signed(input_fmap_173[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_174[7:0]) +
	( 16'sd 29937) * $signed(input_fmap_175[7:0]) +
	( 16'sd 19047) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7854) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14583) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15259) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26385) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6234) * $signed(input_fmap_181[7:0]) +
	( 16'sd 25373) * $signed(input_fmap_182[7:0]) +
	( 16'sd 32358) * $signed(input_fmap_183[7:0]) +
	( 13'sd 2460) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17437) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2610) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1687) * $signed(input_fmap_187[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26438) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17415) * $signed(input_fmap_190[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_191[7:0]) +
	( 16'sd 21642) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9085) * $signed(input_fmap_193[7:0]) +
	( 15'sd 8821) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14775) * $signed(input_fmap_195[7:0]) +
	( 13'sd 2835) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5965) * $signed(input_fmap_197[7:0]) +
	( 16'sd 23531) * $signed(input_fmap_198[7:0]) +
	( 15'sd 8474) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8573) * $signed(input_fmap_200[7:0]) +
	( 14'sd 7745) * $signed(input_fmap_201[7:0]) +
	( 12'sd 1066) * $signed(input_fmap_202[7:0]) +
	( 16'sd 26280) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4865) * $signed(input_fmap_204[7:0]) +
	( 16'sd 20450) * $signed(input_fmap_205[7:0]) +
	( 16'sd 32363) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29448) * $signed(input_fmap_207[7:0]) +
	( 10'sd 281) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15360) * $signed(input_fmap_210[7:0]) +
	( 16'sd 21704) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14496) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3058) * $signed(input_fmap_213[7:0]) +
	( 15'sd 11550) * $signed(input_fmap_214[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_215[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_216[7:0]) +
	( 16'sd 23568) * $signed(input_fmap_217[7:0]) +
	( 16'sd 23933) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17566) * $signed(input_fmap_219[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25587) * $signed(input_fmap_221[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_222[7:0]) +
	( 16'sd 29297) * $signed(input_fmap_223[7:0]) +
	( 15'sd 16374) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1213) * $signed(input_fmap_225[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_226[7:0]) +
	( 16'sd 31290) * $signed(input_fmap_227[7:0]) +
	( 16'sd 17836) * $signed(input_fmap_228[7:0]) +
	( 16'sd 25169) * $signed(input_fmap_229[7:0]) +
	( 15'sd 11200) * $signed(input_fmap_230[7:0]) +
	( 14'sd 5459) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9617) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10315) * $signed(input_fmap_233[7:0]) +
	( 12'sd 1456) * $signed(input_fmap_234[7:0]) +
	( 15'sd 13252) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5557) * $signed(input_fmap_236[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_237[7:0]) +
	( 16'sd 18860) * $signed(input_fmap_238[7:0]) +
	( 14'sd 8188) * $signed(input_fmap_239[7:0]) +
	( 14'sd 8150) * $signed(input_fmap_240[7:0]) +
	( 13'sd 2114) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23208) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13151) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3248) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19300) * $signed(input_fmap_246[7:0]) +
	( 16'sd 23080) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13268) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3363) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30714) * $signed(input_fmap_250[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_251[7:0]) +
	( 16'sd 31723) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25418) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24391) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_83;
assign conv_mac_83 = 
	( 16'sd 32446) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6410) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28768) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19170) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3176) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9366) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18737) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22281) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24551) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6800) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6440) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17416) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17368) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11428) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14252) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4951) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24215) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12156) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18106) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13885) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31584) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25797) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17813) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7728) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15133) * $signed(input_fmap_25[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6627) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22463) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11015) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29352) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10324) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5160) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10562) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30795) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14699) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6690) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12150) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7861) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9520) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23945) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11018) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26449) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32623) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20739) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6874) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12776) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5585) * $signed(input_fmap_50[7:0]) +
	( 12'sd 2015) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12703) * $signed(input_fmap_52[7:0]) +
	( 9'sd 168) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7114) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5747) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28967) * $signed(input_fmap_58[7:0]) +
	( 11'sd 602) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25984) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15945) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31774) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10392) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17865) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13890) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19336) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14004) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15768) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10030) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12881) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18771) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16903) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14480) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25852) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19537) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23534) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21791) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19825) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15322) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20351) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30812) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5979) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27320) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18674) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17796) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9755) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23459) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8021) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13380) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32123) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26572) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22536) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13271) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30888) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8253) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13845) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16680) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20525) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6221) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12575) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20990) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30500) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32061) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14294) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13950) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9294) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20410) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21985) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1225) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29812) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17124) * $signed(input_fmap_119[7:0]) +
	( 11'sd 560) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11296) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1500) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2382) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27862) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1303) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18724) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2569) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27503) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25625) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19760) * $signed(input_fmap_131[7:0]) +
	( 13'sd 3150) * $signed(input_fmap_132[7:0]) +
	( 14'sd 7388) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5047) * $signed(input_fmap_134[7:0]) +
	( 14'sd 7031) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13391) * $signed(input_fmap_136[7:0]) +
	( 14'sd 5318) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9649) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28421) * $signed(input_fmap_140[7:0]) +
	( 16'sd 23872) * $signed(input_fmap_141[7:0]) +
	( 16'sd 23898) * $signed(input_fmap_142[7:0]) +
	( 16'sd 25493) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9548) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_145[7:0]) +
	( 16'sd 22783) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26135) * $signed(input_fmap_148[7:0]) +
	( 16'sd 32648) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27006) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14696) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25717) * $signed(input_fmap_153[7:0]) +
	( 16'sd 19052) * $signed(input_fmap_154[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_155[7:0]) +
	( 16'sd 31496) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15232) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4876) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21337) * $signed(input_fmap_159[7:0]) +
	( 13'sd 3772) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22459) * $signed(input_fmap_161[7:0]) +
	( 14'sd 5374) * $signed(input_fmap_162[7:0]) +
	( 15'sd 10170) * $signed(input_fmap_163[7:0]) +
	( 16'sd 18352) * $signed(input_fmap_164[7:0]) +
	( 16'sd 29560) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2310) * $signed(input_fmap_166[7:0]) +
	( 16'sd 21412) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14635) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25450) * $signed(input_fmap_169[7:0]) +
	( 12'sd 1740) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15628) * $signed(input_fmap_171[7:0]) +
	( 16'sd 27519) * $signed(input_fmap_172[7:0]) +
	( 16'sd 30148) * $signed(input_fmap_173[7:0]) +
	( 16'sd 28389) * $signed(input_fmap_174[7:0]) +
	( 16'sd 30074) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18175) * $signed(input_fmap_177[7:0]) +
	( 14'sd 7307) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28323) * $signed(input_fmap_179[7:0]) +
	( 16'sd 20018) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_181[7:0]) +
	( 13'sd 2682) * $signed(input_fmap_182[7:0]) +
	( 15'sd 11356) * $signed(input_fmap_183[7:0]) +
	( 14'sd 4461) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24939) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18425) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18391) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1506) * $signed(input_fmap_188[7:0]) +
	( 15'sd 15101) * $signed(input_fmap_189[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_190[7:0]) +
	( 15'sd 15018) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22903) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26582) * $signed(input_fmap_194[7:0]) +
	( 14'sd 7918) * $signed(input_fmap_195[7:0]) +
	( 15'sd 10970) * $signed(input_fmap_196[7:0]) +
	( 13'sd 3524) * $signed(input_fmap_197[7:0]) +
	( 16'sd 23372) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20297) * $signed(input_fmap_199[7:0]) +
	( 15'sd 9352) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9961) * $signed(input_fmap_201[7:0]) +
	( 16'sd 23340) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13852) * $signed(input_fmap_203[7:0]) +
	( 16'sd 28496) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28189) * $signed(input_fmap_205[7:0]) +
	( 16'sd 30148) * $signed(input_fmap_206[7:0]) +
	( 16'sd 32386) * $signed(input_fmap_207[7:0]) +
	( 14'sd 7172) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3302) * $signed(input_fmap_209[7:0]) +
	( 14'sd 7987) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5352) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24719) * $signed(input_fmap_212[7:0]) +
	( 16'sd 20325) * $signed(input_fmap_213[7:0]) +
	( 15'sd 8501) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7989) * $signed(input_fmap_215[7:0]) +
	( 16'sd 16549) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_217[7:0]) +
	( 13'sd 3966) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10835) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1182) * $signed(input_fmap_220[7:0]) +
	( 16'sd 16845) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2734) * $signed(input_fmap_222[7:0]) +
	( 11'sd 643) * $signed(input_fmap_223[7:0]) +
	( 15'sd 8258) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_225[7:0]) +
	( 15'sd 16282) * $signed(input_fmap_226[7:0]) +
	( 14'sd 7283) * $signed(input_fmap_227[7:0]) +
	( 11'sd 931) * $signed(input_fmap_228[7:0]) +
	( 16'sd 16985) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30985) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14062) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18602) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24283) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4570) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_235[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_236[7:0]) +
	( 15'sd 8698) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13833) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9830) * $signed(input_fmap_239[7:0]) +
	( 16'sd 16900) * $signed(input_fmap_240[7:0]) +
	( 12'sd 1078) * $signed(input_fmap_241[7:0]) +
	( 16'sd 20688) * $signed(input_fmap_242[7:0]) +
	( 16'sd 26773) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20821) * $signed(input_fmap_244[7:0]) +
	( 16'sd 21092) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9459) * $signed(input_fmap_246[7:0]) +
	( 14'sd 7297) * $signed(input_fmap_247[7:0]) +
	( 15'sd 8773) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9698) * $signed(input_fmap_249[7:0]) +
	( 15'sd 11034) * $signed(input_fmap_250[7:0]) +
	( 15'sd 11459) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2914) * $signed(input_fmap_252[7:0]) +
	( 15'sd 14707) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13818) * $signed(input_fmap_254[7:0]) +
	( 15'sd 12394) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_84;
assign conv_mac_84 = 
	( 14'sd 4293) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26086) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18443) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26599) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30409) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20327) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18509) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7048) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19188) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26744) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7034) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1448) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31215) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14890) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6953) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21120) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18483) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7171) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12413) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16542) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30038) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21557) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31646) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11178) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29299) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5813) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25167) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3759) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32487) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19448) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32067) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14935) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3218) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3183) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2785) * $signed(input_fmap_41[7:0]) +
	( 10'sd 506) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30931) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29391) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9936) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21641) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20880) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10600) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31472) * $signed(input_fmap_51[7:0]) +
	( 11'sd 908) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14567) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22063) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12002) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3703) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16957) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26617) * $signed(input_fmap_59[7:0]) +
	( 14'sd 8146) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30623) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12565) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1050) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24088) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23792) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5962) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5186) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31645) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20558) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20107) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6197) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5570) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2181) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7846) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21642) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7022) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7802) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16267) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5356) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6900) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28079) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4773) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4963) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29128) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7261) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20646) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2230) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20939) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20997) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16039) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22366) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15838) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1546) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3356) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24651) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21369) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8513) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11075) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24655) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8547) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13299) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16139) * $signed(input_fmap_108[7:0]) +
	( 10'sd 505) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5419) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28371) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20223) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15684) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23082) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23056) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16394) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1160) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10426) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22115) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12139) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29165) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23991) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4329) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17274) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8450) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19120) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18941) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10109) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_130[7:0]) +
	( 16'sd 17356) * $signed(input_fmap_131[7:0]) +
	( 13'sd 4091) * $signed(input_fmap_132[7:0]) +
	( 15'sd 8571) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1974) * $signed(input_fmap_134[7:0]) +
	( 14'sd 6284) * $signed(input_fmap_135[7:0]) +
	( 13'sd 3054) * $signed(input_fmap_136[7:0]) +
	( 16'sd 21800) * $signed(input_fmap_137[7:0]) +
	( 16'sd 24080) * $signed(input_fmap_138[7:0]) +
	( 16'sd 29395) * $signed(input_fmap_139[7:0]) +
	( 16'sd 23208) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19470) * $signed(input_fmap_141[7:0]) +
	( 14'sd 7569) * $signed(input_fmap_142[7:0]) +
	( 13'sd 3027) * $signed(input_fmap_143[7:0]) +
	( 15'sd 10772) * $signed(input_fmap_144[7:0]) +
	( 16'sd 31672) * $signed(input_fmap_145[7:0]) +
	( 16'sd 25945) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19204) * $signed(input_fmap_147[7:0]) +
	( 14'sd 7885) * $signed(input_fmap_148[7:0]) +
	( 15'sd 11411) * $signed(input_fmap_149[7:0]) +
	( 15'sd 11622) * $signed(input_fmap_150[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_151[7:0]) +
	( 15'sd 11866) * $signed(input_fmap_152[7:0]) +
	( 16'sd 19645) * $signed(input_fmap_153[7:0]) +
	( 13'sd 2263) * $signed(input_fmap_154[7:0]) +
	( 15'sd 14915) * $signed(input_fmap_155[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24747) * $signed(input_fmap_157[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_158[7:0]) +
	( 16'sd 23715) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22705) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20102) * $signed(input_fmap_161[7:0]) +
	( 16'sd 22383) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22834) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2107) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4341) * $signed(input_fmap_166[7:0]) +
	( 16'sd 18560) * $signed(input_fmap_167[7:0]) +
	( 15'sd 11906) * $signed(input_fmap_168[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_169[7:0]) +
	( 15'sd 12008) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24792) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3967) * $signed(input_fmap_172[7:0]) +
	( 13'sd 2931) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10268) * $signed(input_fmap_174[7:0]) +
	( 15'sd 11784) * $signed(input_fmap_175[7:0]) +
	( 14'sd 6924) * $signed(input_fmap_176[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15033) * $signed(input_fmap_178[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_179[7:0]) +
	( 13'sd 2561) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25530) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30307) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29874) * $signed(input_fmap_183[7:0]) +
	( 14'sd 8153) * $signed(input_fmap_184[7:0]) +
	( 15'sd 10986) * $signed(input_fmap_185[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_186[7:0]) +
	( 16'sd 16943) * $signed(input_fmap_187[7:0]) +
	( 16'sd 26780) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5297) * $signed(input_fmap_190[7:0]) +
	( 16'sd 18822) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15346) * $signed(input_fmap_192[7:0]) +
	( 16'sd 16757) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18244) * $signed(input_fmap_194[7:0]) +
	( 15'sd 9010) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11856) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31669) * $signed(input_fmap_197[7:0]) +
	( 16'sd 25625) * $signed(input_fmap_198[7:0]) +
	( 13'sd 2482) * $signed(input_fmap_199[7:0]) +
	( 16'sd 22025) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11458) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17344) * $signed(input_fmap_202[7:0]) +
	( 13'sd 4020) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15416) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1126) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21042) * $signed(input_fmap_206[7:0]) +
	( 16'sd 31546) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11979) * $signed(input_fmap_208[7:0]) +
	( 15'sd 8736) * $signed(input_fmap_209[7:0]) +
	( 15'sd 8343) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_211[7:0]) +
	( 16'sd 23874) * $signed(input_fmap_212[7:0]) +
	( 16'sd 17212) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4758) * $signed(input_fmap_216[7:0]) +
	( 16'sd 16601) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8622) * $signed(input_fmap_218[7:0]) +
	( 15'sd 8846) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1213) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23674) * $signed(input_fmap_221[7:0]) +
	( 14'sd 8117) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6851) * $signed(input_fmap_224[7:0]) +
	( 16'sd 28753) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_226[7:0]) +
	( 16'sd 17278) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31242) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6336) * $signed(input_fmap_229[7:0]) +
	( 16'sd 21224) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7179) * $signed(input_fmap_231[7:0]) +
	( 14'sd 5301) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_233[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11871) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11367) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6222) * $signed(input_fmap_237[7:0]) +
	( 15'sd 11274) * $signed(input_fmap_238[7:0]) +
	( 15'sd 14445) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_240[7:0]) +
	( 15'sd 10856) * $signed(input_fmap_241[7:0]) +
	( 14'sd 4550) * $signed(input_fmap_242[7:0]) +
	( 13'sd 3977) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24414) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10232) * $signed(input_fmap_245[7:0]) +
	( 15'sd 12324) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30713) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3669) * $signed(input_fmap_248[7:0]) +
	( 12'sd 1667) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21849) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27352) * $signed(input_fmap_252[7:0]) +
	( 16'sd 16661) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13531) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24981) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_85;
assign conv_mac_85 = 
	( 16'sd 31635) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6559) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4403) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17854) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16446) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7608) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11726) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17949) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18790) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17237) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23096) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1348) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8781) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6273) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14707) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13199) * $signed(input_fmap_17[7:0]) +
	( 15'sd 16313) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21414) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6683) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3011) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25090) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31078) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24138) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24969) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21476) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22545) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29733) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19925) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5774) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7422) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29742) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32362) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29705) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31137) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12380) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21659) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14573) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15495) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1457) * $signed(input_fmap_42[7:0]) +
	( 14'sd 4985) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17727) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13225) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19472) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24795) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6164) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16389) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26352) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6358) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_54[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23856) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18544) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24532) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15582) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4603) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21557) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12048) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12367) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32398) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31653) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27140) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27327) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21577) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9521) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7628) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3465) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19015) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11972) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16061) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32016) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7270) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10777) * $signed(input_fmap_79[7:0]) +
	( 15'sd 16067) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19674) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31169) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30924) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26990) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2483) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18173) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19239) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7002) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12827) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24141) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31347) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12080) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20931) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31535) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8543) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1504) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29268) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6007) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17089) * $signed(input_fmap_102[7:0]) +
	( 11'sd 568) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6642) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9459) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27905) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14391) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26104) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30321) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6896) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31308) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27275) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28436) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19790) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30324) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21678) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10307) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3538) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25085) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22106) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30667) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22908) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29242) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18030) * $signed(input_fmap_125[7:0]) +
	( 16'sd 22781) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11715) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17422) * $signed(input_fmap_128[7:0]) +
	( 9'sd 193) * $signed(input_fmap_129[7:0]) +
	( 15'sd 9099) * $signed(input_fmap_130[7:0]) +
	( 15'sd 9482) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14930) * $signed(input_fmap_132[7:0]) +
	( 13'sd 2451) * $signed(input_fmap_133[7:0]) +
	( 16'sd 17349) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18079) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2260) * $signed(input_fmap_136[7:0]) +
	( 16'sd 28518) * $signed(input_fmap_137[7:0]) +
	( 14'sd 5373) * $signed(input_fmap_138[7:0]) +
	( 16'sd 19480) * $signed(input_fmap_139[7:0]) +
	( 16'sd 32051) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22332) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_142[7:0]) +
	( 16'sd 21486) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22249) * $signed(input_fmap_144[7:0]) +
	( 16'sd 18173) * $signed(input_fmap_145[7:0]) +
	( 16'sd 31901) * $signed(input_fmap_146[7:0]) +
	( 16'sd 31937) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20782) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15886) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15244) * $signed(input_fmap_150[7:0]) +
	( 16'sd 20985) * $signed(input_fmap_151[7:0]) +
	( 15'sd 9188) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1504) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10906) * $signed(input_fmap_154[7:0]) +
	( 15'sd 9664) * $signed(input_fmap_155[7:0]) +
	( 11'sd 746) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11359) * $signed(input_fmap_157[7:0]) +
	( 16'sd 21262) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6292) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21470) * $signed(input_fmap_160[7:0]) +
	( 15'sd 11097) * $signed(input_fmap_161[7:0]) +
	( 16'sd 18001) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24108) * $signed(input_fmap_163[7:0]) +
	( 11'sd 689) * $signed(input_fmap_164[7:0]) +
	( 16'sd 25641) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9848) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30697) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4362) * $signed(input_fmap_168[7:0]) +
	( 16'sd 22244) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18896) * $signed(input_fmap_170[7:0]) +
	( 16'sd 17019) * $signed(input_fmap_171[7:0]) +
	( 15'sd 10735) * $signed(input_fmap_172[7:0]) +
	( 10'sd 324) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32434) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7678) * $signed(input_fmap_175[7:0]) +
	( 15'sd 8899) * $signed(input_fmap_176[7:0]) +
	( 16'sd 17456) * $signed(input_fmap_177[7:0]) +
	( 16'sd 25413) * $signed(input_fmap_178[7:0]) +
	( 15'sd 16133) * $signed(input_fmap_179[7:0]) +
	( 15'sd 13045) * $signed(input_fmap_180[7:0]) +
	( 14'sd 8013) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_182[7:0]) +
	( 16'sd 18433) * $signed(input_fmap_183[7:0]) +
	( 16'sd 21976) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15927) * $signed(input_fmap_185[7:0]) +
	( 6'sd 28) * $signed(input_fmap_186[7:0]) +
	( 16'sd 20222) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1152) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11918) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_190[7:0]) +
	( 15'sd 13643) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31971) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22545) * $signed(input_fmap_193[7:0]) +
	( 11'sd 784) * $signed(input_fmap_194[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_195[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_196[7:0]) +
	( 16'sd 27454) * $signed(input_fmap_197[7:0]) +
	( 16'sd 26832) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16350) * $signed(input_fmap_199[7:0]) +
	( 16'sd 27942) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13873) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2872) * $signed(input_fmap_202[7:0]) +
	( 16'sd 27508) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24402) * $signed(input_fmap_205[7:0]) +
	( 16'sd 22068) * $signed(input_fmap_206[7:0]) +
	( 16'sd 25758) * $signed(input_fmap_207[7:0]) +
	( 13'sd 2864) * $signed(input_fmap_208[7:0]) +
	( 16'sd 27370) * $signed(input_fmap_209[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_210[7:0]) +
	( 16'sd 21509) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19632) * $signed(input_fmap_212[7:0]) +
	( 14'sd 7546) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1268) * $signed(input_fmap_214[7:0]) +
	( 16'sd 26041) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28314) * $signed(input_fmap_216[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3685) * $signed(input_fmap_219[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6298) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12420) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9968) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19182) * $signed(input_fmap_224[7:0]) +
	( 15'sd 10461) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31985) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27306) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25782) * $signed(input_fmap_228[7:0]) +
	( 16'sd 25016) * $signed(input_fmap_229[7:0]) +
	( 16'sd 20197) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1354) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7338) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23946) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3770) * $signed(input_fmap_234[7:0]) +
	( 16'sd 18572) * $signed(input_fmap_235[7:0]) +
	( 16'sd 24029) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11281) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22235) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13215) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31858) * $signed(input_fmap_240[7:0]) +
	( 14'sd 6441) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28874) * $signed(input_fmap_242[7:0]) +
	( 16'sd 30090) * $signed(input_fmap_243[7:0]) +
	( 15'sd 8708) * $signed(input_fmap_244[7:0]) +
	( 16'sd 27002) * $signed(input_fmap_245[7:0]) +
	( 15'sd 12020) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18296) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13464) * $signed(input_fmap_248[7:0]) +
	( 15'sd 11474) * $signed(input_fmap_249[7:0]) +
	( 15'sd 14573) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12644) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28124) * $signed(input_fmap_252[7:0]) +
	( 16'sd 23472) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5844) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14296) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_86;
assign conv_mac_86 = 
	( 16'sd 21191) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16376) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30590) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3520) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2947) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9362) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31855) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12125) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9027) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7948) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21540) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18833) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9147) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20665) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28613) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11602) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17657) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31571) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14106) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13832) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7836) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21799) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28601) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15376) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28778) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6065) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19154) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5397) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20172) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25868) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27136) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18582) * $signed(input_fmap_36[7:0]) +
	( 14'sd 8181) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19982) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24482) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12071) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4576) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31975) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24371) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21075) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5172) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11611) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12874) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26013) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16461) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30984) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29855) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8235) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2552) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8293) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4695) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8695) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16911) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25355) * $signed(input_fmap_61[7:0]) +
	( 5'sd 15) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30619) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31939) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20248) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3086) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30080) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21212) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32641) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10451) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17559) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25665) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26948) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17008) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24771) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8558) * $signed(input_fmap_78[7:0]) +
	( 11'sd 583) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28413) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28194) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24363) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24284) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6024) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19435) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13391) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32508) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27333) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3618) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10158) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22006) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2594) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14083) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29356) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21170) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19507) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18519) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6332) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3884) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30608) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13082) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22959) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19060) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27704) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19000) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2683) * $signed(input_fmap_108[7:0]) +
	( 11'sd 871) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12267) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23869) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21322) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12850) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17380) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16549) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25580) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28600) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17960) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20412) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31127) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29811) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7141) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22923) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8325) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18398) * $signed(input_fmap_128[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_129[7:0]) +
	( 16'sd 32111) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24305) * $signed(input_fmap_131[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3694) * $signed(input_fmap_134[7:0]) +
	( 11'sd 780) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12122) * $signed(input_fmap_136[7:0]) +
	( 16'sd 17992) * $signed(input_fmap_137[7:0]) +
	( 16'sd 28813) * $signed(input_fmap_138[7:0]) +
	( 9'sd 241) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22628) * $signed(input_fmap_141[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17511) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6549) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2761) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14463) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17146) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_148[7:0]) +
	( 16'sd 28397) * $signed(input_fmap_149[7:0]) +
	( 16'sd 22033) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6328) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29183) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3070) * $signed(input_fmap_153[7:0]) +
	( 16'sd 26872) * $signed(input_fmap_154[7:0]) +
	( 14'sd 6115) * $signed(input_fmap_155[7:0]) +
	( 16'sd 16816) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11114) * $signed(input_fmap_157[7:0]) +
	( 16'sd 24489) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2430) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18739) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4795) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26929) * $signed(input_fmap_162[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_163[7:0]) +
	( 14'sd 5334) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23916) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18805) * $signed(input_fmap_166[7:0]) +
	( 13'sd 3776) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1371) * $signed(input_fmap_168[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23717) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12765) * $signed(input_fmap_171[7:0]) +
	( 16'sd 16571) * $signed(input_fmap_172[7:0]) +
	( 16'sd 24921) * $signed(input_fmap_173[7:0]) +
	( 16'sd 20701) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10030) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29473) * $signed(input_fmap_177[7:0]) +
	( 13'sd 3293) * $signed(input_fmap_178[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4134) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28691) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12776) * $signed(input_fmap_182[7:0]) +
	( 16'sd 22196) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24338) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1868) * $signed(input_fmap_185[7:0]) +
	( 16'sd 16832) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27692) * $signed(input_fmap_187[7:0]) +
	( 10'sd 416) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19512) * $signed(input_fmap_189[7:0]) +
	( 13'sd 2806) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3246) * $signed(input_fmap_191[7:0]) +
	( 16'sd 21957) * $signed(input_fmap_192[7:0]) +
	( 16'sd 21112) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26199) * $signed(input_fmap_194[7:0]) +
	( 14'sd 7987) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_196[7:0]) +
	( 16'sd 29926) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27786) * $signed(input_fmap_198[7:0]) +
	( 15'sd 8595) * $signed(input_fmap_199[7:0]) +
	( 14'sd 4655) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11541) * $signed(input_fmap_201[7:0]) +
	( 16'sd 32468) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24028) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12835) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2910) * $signed(input_fmap_205[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_206[7:0]) +
	( 15'sd 14762) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19141) * $signed(input_fmap_210[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_211[7:0]) +
	( 16'sd 23401) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28223) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18791) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11361) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11032) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30555) * $signed(input_fmap_218[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21064) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12413) * $signed(input_fmap_221[7:0]) +
	( 15'sd 16213) * $signed(input_fmap_222[7:0]) +
	( 16'sd 31093) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27825) * $signed(input_fmap_224[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_225[7:0]) +
	( 11'sd 756) * $signed(input_fmap_226[7:0]) +
	( 16'sd 32113) * $signed(input_fmap_227[7:0]) +
	( 15'sd 12333) * $signed(input_fmap_228[7:0]) +
	( 11'sd 897) * $signed(input_fmap_229[7:0]) +
	( 13'sd 3037) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18998) * $signed(input_fmap_231[7:0]) +
	( 16'sd 32612) * $signed(input_fmap_232[7:0]) +
	( 15'sd 12424) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_234[7:0]) +
	( 15'sd 8463) * $signed(input_fmap_235[7:0]) +
	( 16'sd 24280) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14562) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28696) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19462) * $signed(input_fmap_239[7:0]) +
	( 14'sd 7338) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7415) * $signed(input_fmap_241[7:0]) +
	( 16'sd 25962) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2828) * $signed(input_fmap_243[7:0]) +
	( 14'sd 5377) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7060) * $signed(input_fmap_245[7:0]) +
	( 16'sd 24339) * $signed(input_fmap_246[7:0]) +
	( 11'sd 775) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10159) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17050) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4515) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_252[7:0]) +
	( 16'sd 21538) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_254[7:0]) +
	( 12'sd 1292) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_87;
assign conv_mac_87 = 
	( 10'sd 466) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1368) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8533) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6756) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32414) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7185) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17926) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11504) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18613) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28697) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5166) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2067) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4777) * $signed(input_fmap_12[7:0]) +
	( 13'sd 4081) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28134) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9407) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16196) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18775) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15408) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23802) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2228) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18456) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23383) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11595) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28152) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8876) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29684) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27530) * $signed(input_fmap_32[7:0]) +
	( 16'sd 17106) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26743) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4172) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30380) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22621) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30133) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8567) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12583) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27232) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23901) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22532) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6839) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15979) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18228) * $signed(input_fmap_48[7:0]) +
	( 11'sd 585) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18126) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5539) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14930) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25014) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12680) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5475) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9956) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6402) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30486) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17236) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20689) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2686) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14530) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10984) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20677) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7055) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3014) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20471) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24539) * $signed(input_fmap_70[7:0]) +
	( 16'sd 22319) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20804) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16147) * $signed(input_fmap_73[7:0]) +
	( 8'sd 95) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11162) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15078) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19046) * $signed(input_fmap_79[7:0]) +
	( 10'sd 342) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30313) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21338) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9885) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23840) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2540) * $signed(input_fmap_86[7:0]) +
	( 10'sd 391) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24458) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10888) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19942) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14213) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21176) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14822) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2630) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25764) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20292) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22357) * $signed(input_fmap_98[7:0]) +
	( 11'sd 871) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6432) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24365) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31846) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20880) * $signed(input_fmap_103[7:0]) +
	( 11'sd 866) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13965) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12197) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3236) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30164) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12866) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16037) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29781) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27185) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23512) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26447) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18547) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13811) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16824) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2128) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24371) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26438) * $signed(input_fmap_123[7:0]) +
	( 11'sd 939) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25875) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16981) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22881) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15752) * $signed(input_fmap_128[7:0]) +
	( 13'sd 2728) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30556) * $signed(input_fmap_130[7:0]) +
	( 16'sd 29475) * $signed(input_fmap_131[7:0]) +
	( 15'sd 12395) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10144) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2220) * $signed(input_fmap_134[7:0]) +
	( 13'sd 3290) * $signed(input_fmap_135[7:0]) +
	( 14'sd 5871) * $signed(input_fmap_136[7:0]) +
	( 13'sd 3651) * $signed(input_fmap_137[7:0]) +
	( 13'sd 3053) * $signed(input_fmap_138[7:0]) +
	( 16'sd 29810) * $signed(input_fmap_139[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_140[7:0]) +
	( 16'sd 25243) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11732) * $signed(input_fmap_142[7:0]) +
	( 15'sd 13043) * $signed(input_fmap_143[7:0]) +
	( 12'sd 1305) * $signed(input_fmap_144[7:0]) +
	( 14'sd 4566) * $signed(input_fmap_145[7:0]) +
	( 14'sd 4315) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_148[7:0]) +
	( 15'sd 13004) * $signed(input_fmap_149[7:0]) +
	( 12'sd 1298) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3296) * $signed(input_fmap_151[7:0]) +
	( 14'sd 4300) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1893) * $signed(input_fmap_153[7:0]) +
	( 16'sd 28155) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_155[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5646) * $signed(input_fmap_157[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_158[7:0]) +
	( 16'sd 19106) * $signed(input_fmap_159[7:0]) +
	( 15'sd 8884) * $signed(input_fmap_160[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_161[7:0]) +
	( 16'sd 32096) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22787) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8831) * $signed(input_fmap_164[7:0]) +
	( 16'sd 21269) * $signed(input_fmap_165[7:0]) +
	( 14'sd 6665) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30072) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9242) * $signed(input_fmap_168[7:0]) +
	( 16'sd 31844) * $signed(input_fmap_169[7:0]) +
	( 16'sd 30665) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19394) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1571) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23613) * $signed(input_fmap_173[7:0]) +
	( 12'sd 1185) * $signed(input_fmap_174[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_175[7:0]) +
	( 16'sd 32133) * $signed(input_fmap_176[7:0]) +
	( 15'sd 13191) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2273) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15257) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26292) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23313) * $signed(input_fmap_181[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29142) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22221) * $signed(input_fmap_184[7:0]) +
	( 16'sd 21284) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13764) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11729) * $signed(input_fmap_187[7:0]) +
	( 16'sd 16781) * $signed(input_fmap_188[7:0]) +
	( 15'sd 10826) * $signed(input_fmap_189[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_190[7:0]) +
	( 16'sd 30322) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24080) * $signed(input_fmap_192[7:0]) +
	( 13'sd 2867) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9040) * $signed(input_fmap_194[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15955) * $signed(input_fmap_196[7:0]) +
	( 15'sd 13129) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5346) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10334) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13174) * $signed(input_fmap_200[7:0]) +
	( 16'sd 20038) * $signed(input_fmap_201[7:0]) +
	( 11'sd 776) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30992) * $signed(input_fmap_203[7:0]) +
	( 12'sd 1490) * $signed(input_fmap_204[7:0]) +
	( 15'sd 10129) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29330) * $signed(input_fmap_206[7:0]) +
	( 15'sd 8867) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30138) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7629) * $signed(input_fmap_209[7:0]) +
	( 14'sd 8187) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17312) * $signed(input_fmap_211[7:0]) +
	( 16'sd 25722) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9762) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18804) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17985) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_216[7:0]) +
	( 15'sd 15963) * $signed(input_fmap_217[7:0]) +
	( 16'sd 16714) * $signed(input_fmap_218[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24457) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13714) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_224[7:0]) +
	( 16'sd 17270) * $signed(input_fmap_225[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9382) * $signed(input_fmap_227[7:0]) +
	( 15'sd 16086) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23182) * $signed(input_fmap_229[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25949) * $signed(input_fmap_231[7:0]) +
	( 16'sd 21597) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15378) * $signed(input_fmap_233[7:0]) +
	( 16'sd 30244) * $signed(input_fmap_234[7:0]) +
	( 16'sd 18082) * $signed(input_fmap_235[7:0]) +
	( 15'sd 14772) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28442) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16789) * $signed(input_fmap_238[7:0]) +
	( 11'sd 723) * $signed(input_fmap_239[7:0]) +
	( 16'sd 21808) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15378) * $signed(input_fmap_241[7:0]) +
	( 10'sd 284) * $signed(input_fmap_242[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_244[7:0]) +
	( 15'sd 15049) * $signed(input_fmap_245[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13678) * $signed(input_fmap_247[7:0]) +
	( 15'sd 14922) * $signed(input_fmap_248[7:0]) +
	( 15'sd 8324) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3485) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_251[7:0]) +
	( 15'sd 11844) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6965) * $signed(input_fmap_253[7:0]) +
	( 16'sd 22402) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5941) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_88;
assign conv_mac_88 = 
	( 16'sd 26659) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21707) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4579) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28677) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7637) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5347) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28193) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25902) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14153) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25054) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21079) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19330) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13098) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6084) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9291) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12001) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5561) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3196) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21305) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10014) * $signed(input_fmap_22[7:0]) +
	( 11'sd 677) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3297) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15173) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23402) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24079) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19313) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24824) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13260) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2273) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19761) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17520) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26132) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6268) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9422) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10719) * $signed(input_fmap_38[7:0]) +
	( 11'sd 870) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25881) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20399) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3694) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11382) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20709) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23821) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13461) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23105) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4761) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21003) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18648) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14602) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19153) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24835) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31834) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7614) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30234) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16271) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6921) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3127) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15134) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6872) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25678) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25002) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19841) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25895) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6529) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10121) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15119) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7447) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6271) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2535) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11386) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4334) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_80[7:0]) +
	( 14'sd 8021) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10650) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10874) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10334) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6828) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17249) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18189) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17445) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11270) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15571) * $signed(input_fmap_90[7:0]) +
	( 10'sd 347) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7127) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26775) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29407) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12459) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24207) * $signed(input_fmap_98[7:0]) +
	( 11'sd 643) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11978) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1438) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21438) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1940) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24709) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7322) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7634) * $signed(input_fmap_107[7:0]) +
	( 14'sd 8168) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16409) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18167) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3096) * $signed(input_fmap_112[7:0]) +
	( 10'sd 265) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15763) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16699) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27847) * $signed(input_fmap_116[7:0]) +
	( 11'sd 802) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31558) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22207) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7539) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21948) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6927) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2539) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4332) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3377) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4931) * $signed(input_fmap_127[7:0]) +
	( 16'sd 24907) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1522) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10604) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8463) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31423) * $signed(input_fmap_133[7:0]) +
	( 16'sd 28698) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26949) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7016) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9543) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10950) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28562) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9408) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13479) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31308) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23212) * $signed(input_fmap_143[7:0]) +
	( 16'sd 23260) * $signed(input_fmap_144[7:0]) +
	( 14'sd 6871) * $signed(input_fmap_145[7:0]) +
	( 16'sd 23930) * $signed(input_fmap_146[7:0]) +
	( 16'sd 20734) * $signed(input_fmap_147[7:0]) +
	( 16'sd 31023) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15273) * $signed(input_fmap_149[7:0]) +
	( 16'sd 22640) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18033) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31197) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12884) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30117) * $signed(input_fmap_154[7:0]) +
	( 16'sd 26733) * $signed(input_fmap_155[7:0]) +
	( 16'sd 27126) * $signed(input_fmap_156[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_157[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_158[7:0]) +
	( 14'sd 8094) * $signed(input_fmap_159[7:0]) +
	( 16'sd 23918) * $signed(input_fmap_160[7:0]) +
	( 13'sd 2529) * $signed(input_fmap_161[7:0]) +
	( 14'sd 6602) * $signed(input_fmap_162[7:0]) +
	( 11'sd 762) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25213) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2305) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30736) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31476) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17227) * $signed(input_fmap_168[7:0]) +
	( 14'sd 5211) * $signed(input_fmap_169[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3621) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31711) * $signed(input_fmap_172[7:0]) +
	( 16'sd 31316) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7742) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_175[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10605) * $signed(input_fmap_178[7:0]) +
	( 12'sd 1108) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3236) * $signed(input_fmap_180[7:0]) +
	( 15'sd 12426) * $signed(input_fmap_181[7:0]) +
	( 13'sd 3811) * $signed(input_fmap_182[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22802) * $signed(input_fmap_184[7:0]) +
	( 16'sd 29179) * $signed(input_fmap_185[7:0]) +
	( 10'sd 387) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5796) * $signed(input_fmap_187[7:0]) +
	( 14'sd 6907) * $signed(input_fmap_188[7:0]) +
	( 16'sd 21235) * $signed(input_fmap_189[7:0]) +
	( 13'sd 3817) * $signed(input_fmap_190[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14952) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6682) * $signed(input_fmap_193[7:0]) +
	( 16'sd 31218) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13060) * $signed(input_fmap_195[7:0]) +
	( 16'sd 32604) * $signed(input_fmap_196[7:0]) +
	( 16'sd 17703) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10766) * $signed(input_fmap_198[7:0]) +
	( 13'sd 3668) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_200[7:0]) +
	( 16'sd 23681) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19818) * $signed(input_fmap_202[7:0]) +
	( 16'sd 20153) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17893) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31131) * $signed(input_fmap_205[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1654) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30615) * $signed(input_fmap_208[7:0]) +
	( 9'sd 158) * $signed(input_fmap_209[7:0]) +
	( 15'sd 13886) * $signed(input_fmap_210[7:0]) +
	( 14'sd 7248) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19896) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11095) * $signed(input_fmap_213[7:0]) +
	( 15'sd 8195) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17205) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4718) * $signed(input_fmap_216[7:0]) +
	( 12'sd 1683) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7807) * $signed(input_fmap_218[7:0]) +
	( 11'sd 756) * $signed(input_fmap_219[7:0]) +
	( 16'sd 32487) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12247) * $signed(input_fmap_222[7:0]) +
	( 15'sd 11096) * $signed(input_fmap_223[7:0]) +
	( 16'sd 28402) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3401) * $signed(input_fmap_225[7:0]) +
	( 12'sd 2022) * $signed(input_fmap_226[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8962) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3061) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18171) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_231[7:0]) +
	( 11'sd 926) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23811) * $signed(input_fmap_233[7:0]) +
	( 15'sd 11307) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31372) * $signed(input_fmap_236[7:0]) +
	( 16'sd 16470) * $signed(input_fmap_237[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20148) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9780) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26673) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29310) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2928) * $signed(input_fmap_243[7:0]) +
	( 13'sd 3739) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22259) * $signed(input_fmap_245[7:0]) +
	( 16'sd 21651) * $signed(input_fmap_246[7:0]) +
	( 15'sd 14127) * $signed(input_fmap_247[7:0]) +
	( 11'sd 575) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30902) * $signed(input_fmap_249[7:0]) +
	( 12'sd 1566) * $signed(input_fmap_250[7:0]) +
	( 15'sd 9888) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20641) * $signed(input_fmap_252[7:0]) +
	( 14'sd 7137) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10285) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5102) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_89;
assign conv_mac_89 = 
	( 16'sd 18258) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17380) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5193) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7708) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4824) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12771) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30545) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17515) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20517) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31228) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14039) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29486) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3799) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15711) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14922) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25791) * $signed(input_fmap_17[7:0]) +
	( 11'sd 841) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15912) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18769) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18367) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29201) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5309) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19090) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24134) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14990) * $signed(input_fmap_27[7:0]) +
	( 8'sd 81) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10098) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10442) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1413) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27140) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12787) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16048) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18233) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19408) * $signed(input_fmap_37[7:0]) +
	( 15'sd 12976) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31141) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7747) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12650) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16983) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28618) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12332) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6975) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9974) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21165) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21545) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4705) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3063) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21886) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18637) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13666) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23519) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20029) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23673) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15893) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1065) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21878) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28040) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25170) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32099) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15426) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20172) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24911) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26303) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14436) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10120) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9945) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22411) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2201) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12284) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5801) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18583) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14163) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3966) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1552) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27952) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32331) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25813) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8661) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14998) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22664) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32696) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26721) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15072) * $signed(input_fmap_92[7:0]) +
	( 9'sd 209) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14525) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23652) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32703) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21139) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9599) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21118) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24368) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20974) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26685) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7793) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29608) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12955) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30258) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24273) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16022) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25372) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13140) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16455) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32624) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6146) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27876) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20243) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12091) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18990) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16257) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6727) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30467) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4461) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10002) * $signed(input_fmap_127[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_128[7:0]) +
	( 11'sd 557) * $signed(input_fmap_129[7:0]) +
	( 16'sd 32372) * $signed(input_fmap_130[7:0]) +
	( 13'sd 2056) * $signed(input_fmap_131[7:0]) +
	( 16'sd 27756) * $signed(input_fmap_132[7:0]) +
	( 16'sd 24521) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5555) * $signed(input_fmap_134[7:0]) +
	( 13'sd 3962) * $signed(input_fmap_135[7:0]) +
	( 13'sd 3348) * $signed(input_fmap_136[7:0]) +
	( 16'sd 30245) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19548) * $signed(input_fmap_138[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3653) * $signed(input_fmap_140[7:0]) +
	( 14'sd 8096) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21321) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_143[7:0]) +
	( 9'sd 180) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25197) * $signed(input_fmap_145[7:0]) +
	( 16'sd 17626) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29404) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17871) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_149[7:0]) +
	( 16'sd 19859) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23401) * $signed(input_fmap_151[7:0]) +
	( 16'sd 27217) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17285) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31230) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7008) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29774) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29549) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8819) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4764) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_160[7:0]) +
	( 14'sd 7373) * $signed(input_fmap_161[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_162[7:0]) +
	( 15'sd 14892) * $signed(input_fmap_163[7:0]) +
	( 16'sd 23447) * $signed(input_fmap_164[7:0]) +
	( 11'sd 980) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8625) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13591) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5206) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18672) * $signed(input_fmap_169[7:0]) +
	( 16'sd 21675) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24369) * $signed(input_fmap_171[7:0]) +
	( 10'sd 457) * $signed(input_fmap_172[7:0]) +
	( 14'sd 7888) * $signed(input_fmap_173[7:0]) +
	( 14'sd 8170) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5297) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_176[7:0]) +
	( 13'sd 3417) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17458) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15838) * $signed(input_fmap_179[7:0]) +
	( 12'sd 1087) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23985) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19414) * $signed(input_fmap_182[7:0]) +
	( 16'sd 28199) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22976) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24406) * $signed(input_fmap_185[7:0]) +
	( 16'sd 28306) * $signed(input_fmap_186[7:0]) +
	( 16'sd 20380) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29466) * $signed(input_fmap_188[7:0]) +
	( 14'sd 6812) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5304) * $signed(input_fmap_191[7:0]) +
	( 16'sd 23454) * $signed(input_fmap_192[7:0]) +
	( 16'sd 16565) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30557) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27333) * $signed(input_fmap_195[7:0]) +
	( 14'sd 4916) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31445) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19300) * $signed(input_fmap_198[7:0]) +
	( 16'sd 31931) * $signed(input_fmap_199[7:0]) +
	( 16'sd 22963) * $signed(input_fmap_200[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_201[7:0]) +
	( 16'sd 24324) * $signed(input_fmap_202[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_204[7:0]) +
	( 14'sd 7497) * $signed(input_fmap_205[7:0]) +
	( 16'sd 26141) * $signed(input_fmap_206[7:0]) +
	( 15'sd 10473) * $signed(input_fmap_207[7:0]) +
	( 16'sd 24554) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30038) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30871) * $signed(input_fmap_211[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23815) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31817) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_215[7:0]) +
	( 15'sd 15301) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17656) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7076) * $signed(input_fmap_218[7:0]) +
	( 15'sd 11662) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30094) * $signed(input_fmap_220[7:0]) +
	( 16'sd 32542) * $signed(input_fmap_221[7:0]) +
	( 16'sd 27722) * $signed(input_fmap_222[7:0]) +
	( 16'sd 31058) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13968) * $signed(input_fmap_224[7:0]) +
	( 16'sd 23217) * $signed(input_fmap_225[7:0]) +
	( 16'sd 23202) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20144) * $signed(input_fmap_227[7:0]) +
	( 15'sd 13178) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26012) * $signed(input_fmap_229[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14868) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9956) * $signed(input_fmap_232[7:0]) +
	( 15'sd 9590) * $signed(input_fmap_233[7:0]) +
	( 14'sd 7045) * $signed(input_fmap_234[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_235[7:0]) +
	( 16'sd 21925) * $signed(input_fmap_236[7:0]) +
	( 14'sd 5068) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27754) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_239[7:0]) +
	( 15'sd 12637) * $signed(input_fmap_240[7:0]) +
	( 16'sd 27777) * $signed(input_fmap_241[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7978) * $signed(input_fmap_243[7:0]) +
	( 14'sd 7222) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22211) * $signed(input_fmap_245[7:0]) +
	( 16'sd 25329) * $signed(input_fmap_246[7:0]) +
	( 15'sd 10020) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18804) * $signed(input_fmap_248[7:0]) +
	( 16'sd 26472) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25464) * $signed(input_fmap_250[7:0]) +
	( 13'sd 3853) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6175) * $signed(input_fmap_252[7:0]) +
	( 16'sd 18906) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26381) * $signed(input_fmap_254[7:0]) +
	( 16'sd 25810) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_90;
assign conv_mac_90 = 
	( 15'sd 12186) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26231) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21387) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32217) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10181) * $signed(input_fmap_5[7:0]) +
	( 8'sd 92) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2908) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26689) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4446) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3960) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15556) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27080) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2731) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1854) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19201) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14756) * $signed(input_fmap_17[7:0]) +
	( 11'sd 967) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16787) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21771) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16999) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25860) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20830) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12313) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8059) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28263) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1235) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3909) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14954) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23003) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11063) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7731) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23791) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31809) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25154) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30721) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18842) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26890) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7717) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22820) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15423) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9569) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31449) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27658) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24710) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15365) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9431) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11175) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19006) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15286) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17234) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21119) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29025) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14500) * $signed(input_fmap_58[7:0]) +
	( 12'sd 2026) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11908) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5882) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30108) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31702) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16209) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14364) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16078) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28617) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9159) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28703) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17523) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28249) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1277) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3391) * $signed(input_fmap_76[7:0]) +
	( 11'sd 677) * $signed(input_fmap_77[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4718) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26375) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2093) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5677) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25381) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4808) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24452) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32323) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32497) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23537) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22032) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28943) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18536) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23647) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30254) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22385) * $signed(input_fmap_99[7:0]) +
	( 11'sd 1007) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3185) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10444) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16026) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26663) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21592) * $signed(input_fmap_106[7:0]) +
	( 13'sd 4044) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19311) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20477) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19380) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4837) * $signed(input_fmap_112[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12550) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28562) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31712) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24045) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22139) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15304) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20436) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6530) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23233) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31000) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27415) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8388) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11876) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_127[7:0]) +
	( 14'sd 6905) * $signed(input_fmap_128[7:0]) +
	( 15'sd 12247) * $signed(input_fmap_129[7:0]) +
	( 15'sd 16243) * $signed(input_fmap_130[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1340) * $signed(input_fmap_132[7:0]) +
	( 16'sd 19952) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_134[7:0]) +
	( 15'sd 11518) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23895) * $signed(input_fmap_136[7:0]) +
	( 16'sd 29865) * $signed(input_fmap_137[7:0]) +
	( 14'sd 5988) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11229) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26041) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5568) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7065) * $signed(input_fmap_143[7:0]) +
	( 15'sd 14656) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21882) * $signed(input_fmap_145[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_146[7:0]) +
	( 16'sd 25710) * $signed(input_fmap_147[7:0]) +
	( 16'sd 24199) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18553) * $signed(input_fmap_149[7:0]) +
	( 14'sd 8068) * $signed(input_fmap_150[7:0]) +
	( 14'sd 7972) * $signed(input_fmap_151[7:0]) +
	( 16'sd 18478) * $signed(input_fmap_152[7:0]) +
	( 11'sd 836) * $signed(input_fmap_153[7:0]) +
	( 16'sd 29889) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7330) * $signed(input_fmap_155[7:0]) +
	( 15'sd 9123) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11295) * $signed(input_fmap_157[7:0]) +
	( 14'sd 7724) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21866) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17117) * $signed(input_fmap_160[7:0]) +
	( 16'sd 27831) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4424) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_163[7:0]) +
	( 16'sd 31354) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4566) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8730) * $signed(input_fmap_166[7:0]) +
	( 9'sd 165) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20528) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6280) * $signed(input_fmap_169[7:0]) +
	( 16'sd 21600) * $signed(input_fmap_170[7:0]) +
	( 16'sd 17601) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11995) * $signed(input_fmap_172[7:0]) +
	( 16'sd 20212) * $signed(input_fmap_173[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1511) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18994) * $signed(input_fmap_177[7:0]) +
	( 16'sd 24089) * $signed(input_fmap_178[7:0]) +
	( 16'sd 19113) * $signed(input_fmap_179[7:0]) +
	( 15'sd 11531) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23607) * $signed(input_fmap_181[7:0]) +
	( 15'sd 13914) * $signed(input_fmap_182[7:0]) +
	( 16'sd 28394) * $signed(input_fmap_183[7:0]) +
	( 6'sd 25) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24023) * $signed(input_fmap_185[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18957) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31593) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17269) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13152) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31859) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27695) * $signed(input_fmap_192[7:0]) +
	( 16'sd 32737) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29569) * $signed(input_fmap_194[7:0]) +
	( 10'sd 496) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11695) * $signed(input_fmap_196[7:0]) +
	( 15'sd 13176) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2249) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24179) * $signed(input_fmap_199[7:0]) +
	( 16'sd 19732) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3183) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7942) * $signed(input_fmap_202[7:0]) +
	( 16'sd 28187) * $signed(input_fmap_203[7:0]) +
	( 16'sd 27177) * $signed(input_fmap_204[7:0]) +
	( 15'sd 9082) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_206[7:0]) +
	( 16'sd 16753) * $signed(input_fmap_207[7:0]) +
	( 15'sd 9491) * $signed(input_fmap_208[7:0]) +
	( 16'sd 28030) * $signed(input_fmap_209[7:0]) +
	( 15'sd 13674) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6483) * $signed(input_fmap_211[7:0]) +
	( 14'sd 6950) * $signed(input_fmap_212[7:0]) +
	( 15'sd 13273) * $signed(input_fmap_213[7:0]) +
	( 14'sd 6615) * $signed(input_fmap_214[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_215[7:0]) +
	( 14'sd 6448) * $signed(input_fmap_216[7:0]) +
	( 13'sd 4092) * $signed(input_fmap_217[7:0]) +
	( 16'sd 19308) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14969) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19081) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12957) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2223) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6316) * $signed(input_fmap_224[7:0]) +
	( 15'sd 16367) * $signed(input_fmap_225[7:0]) +
	( 13'sd 2844) * $signed(input_fmap_226[7:0]) +
	( 16'sd 28293) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10249) * $signed(input_fmap_228[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_229[7:0]) +
	( 11'sd 583) * $signed(input_fmap_230[7:0]) +
	( 14'sd 5963) * $signed(input_fmap_231[7:0]) +
	( 16'sd 31001) * $signed(input_fmap_232[7:0]) +
	( 16'sd 25559) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_234[7:0]) +
	( 16'sd 18741) * $signed(input_fmap_235[7:0]) +
	( 15'sd 15854) * $signed(input_fmap_236[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_237[7:0]) +
	( 16'sd 32075) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12444) * $signed(input_fmap_239[7:0]) +
	( 16'sd 30747) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25391) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5731) * $signed(input_fmap_242[7:0]) +
	( 15'sd 15314) * $signed(input_fmap_243[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7715) * $signed(input_fmap_245[7:0]) +
	( 9'sd 141) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17976) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1740) * $signed(input_fmap_248[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9379) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26704) * $signed(input_fmap_251[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_252[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10287) * $signed(input_fmap_254[7:0]) +
	( 16'sd 16539) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_91;
assign conv_mac_91 = 
	( 14'sd 6901) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8304) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31359) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7676) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32602) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11214) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17138) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2629) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29323) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17057) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18045) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26546) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4780) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25168) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24003) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13717) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20693) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29646) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23660) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15369) * $signed(input_fmap_20[7:0]) +
	( 11'sd 584) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28848) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20079) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26481) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1987) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26997) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21366) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9755) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3627) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32640) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16501) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30060) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13313) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7909) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4680) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23501) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13283) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_41[7:0]) +
	( 11'sd 893) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8961) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2367) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2424) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24119) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27945) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28753) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8746) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30991) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2721) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26106) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18803) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12983) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11715) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16553) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24651) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14368) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30983) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15077) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11824) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12936) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26698) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26311) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29259) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3602) * $signed(input_fmap_70[7:0]) +
	( 12'sd 2026) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3083) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18971) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6225) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9127) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20448) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12333) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31858) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9883) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2710) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1834) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15101) * $signed(input_fmap_83[7:0]) +
	( 16'sd 24615) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27178) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14592) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14607) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25361) * $signed(input_fmap_88[7:0]) +
	( 14'sd 6306) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18612) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23529) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18907) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28894) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29274) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29016) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12479) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12148) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4388) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28127) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2414) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9350) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26934) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24367) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14292) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19466) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_109[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15998) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1541) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22799) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30455) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12776) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12736) * $signed(input_fmap_117[7:0]) +
	( 15'sd 16016) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26815) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21534) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32457) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1302) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6920) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6434) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16444) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1242) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26659) * $signed(input_fmap_127[7:0]) +
	( 16'sd 26813) * $signed(input_fmap_128[7:0]) +
	( 16'sd 21922) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31188) * $signed(input_fmap_130[7:0]) +
	( 16'sd 16575) * $signed(input_fmap_131[7:0]) +
	( 16'sd 26948) * $signed(input_fmap_132[7:0]) +
	( 8'sd 75) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11850) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28792) * $signed(input_fmap_135[7:0]) +
	( 16'sd 29039) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27737) * $signed(input_fmap_137[7:0]) +
	( 13'sd 3604) * $signed(input_fmap_138[7:0]) +
	( 16'sd 22574) * $signed(input_fmap_139[7:0]) +
	( 15'sd 11693) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22147) * $signed(input_fmap_141[7:0]) +
	( 15'sd 13847) * $signed(input_fmap_142[7:0]) +
	( 11'sd 630) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18320) * $signed(input_fmap_144[7:0]) +
	( 13'sd 3114) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17158) * $signed(input_fmap_147[7:0]) +
	( 16'sd 24003) * $signed(input_fmap_148[7:0]) +
	( 8'sd 89) * $signed(input_fmap_149[7:0]) +
	( 10'sd 500) * $signed(input_fmap_150[7:0]) +
	( 15'sd 13404) * $signed(input_fmap_151[7:0]) +
	( 15'sd 12982) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2835) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30961) * $signed(input_fmap_154[7:0]) +
	( 15'sd 16314) * $signed(input_fmap_155[7:0]) +
	( 11'sd 918) * $signed(input_fmap_156[7:0]) +
	( 16'sd 19006) * $signed(input_fmap_157[7:0]) +
	( 16'sd 19714) * $signed(input_fmap_158[7:0]) +
	( 16'sd 25981) * $signed(input_fmap_159[7:0]) +
	( 16'sd 25960) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14497) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2196) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19670) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19737) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4830) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9399) * $signed(input_fmap_167[7:0]) +
	( 15'sd 12300) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30566) * $signed(input_fmap_169[7:0]) +
	( 15'sd 10761) * $signed(input_fmap_170[7:0]) +
	( 15'sd 9940) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9200) * $signed(input_fmap_172[7:0]) +
	( 16'sd 32252) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_174[7:0]) +
	( 16'sd 19694) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1438) * $signed(input_fmap_176[7:0]) +
	( 14'sd 4652) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27836) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28497) * $signed(input_fmap_179[7:0]) +
	( 15'sd 10936) * $signed(input_fmap_180[7:0]) +
	( 13'sd 2450) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_183[7:0]) +
	( 12'sd 1506) * $signed(input_fmap_184[7:0]) +
	( 15'sd 12796) * $signed(input_fmap_185[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_186[7:0]) +
	( 13'sd 3266) * $signed(input_fmap_187[7:0]) +
	( 15'sd 15650) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17151) * $signed(input_fmap_190[7:0]) +
	( 10'sd 366) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28318) * $signed(input_fmap_192[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_193[7:0]) +
	( 15'sd 8428) * $signed(input_fmap_194[7:0]) +
	( 16'sd 20020) * $signed(input_fmap_195[7:0]) +
	( 15'sd 13089) * $signed(input_fmap_196[7:0]) +
	( 16'sd 17940) * $signed(input_fmap_197[7:0]) +
	( 15'sd 8239) * $signed(input_fmap_198[7:0]) +
	( 13'sd 2799) * $signed(input_fmap_199[7:0]) +
	( 16'sd 32254) * $signed(input_fmap_200[7:0]) +
	( 16'sd 17371) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18034) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25073) * $signed(input_fmap_203[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_204[7:0]) +
	( 16'sd 22452) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6899) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17064) * $signed(input_fmap_207[7:0]) +
	( 16'sd 31773) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14378) * $signed(input_fmap_209[7:0]) +
	( 16'sd 22653) * $signed(input_fmap_210[7:0]) +
	( 15'sd 8926) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19769) * $signed(input_fmap_212[7:0]) +
	( 15'sd 15880) * $signed(input_fmap_213[7:0]) +
	( 11'sd 981) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25717) * $signed(input_fmap_215[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_216[7:0]) +
	( 13'sd 3540) * $signed(input_fmap_217[7:0]) +
	( 13'sd 3810) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5452) * $signed(input_fmap_219[7:0]) +
	( 13'sd 3647) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12931) * $signed(input_fmap_221[7:0]) +
	( 16'sd 26300) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15174) * $signed(input_fmap_223[7:0]) +
	( 15'sd 15003) * $signed(input_fmap_224[7:0]) +
	( 7'sd 54) * $signed(input_fmap_225[7:0]) +
	( 16'sd 23977) * $signed(input_fmap_226[7:0]) +
	( 12'sd 1851) * $signed(input_fmap_227[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29254) * $signed(input_fmap_229[7:0]) +
	( 14'sd 4616) * $signed(input_fmap_230[7:0]) +
	( 16'sd 21314) * $signed(input_fmap_231[7:0]) +
	( 16'sd 23355) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_233[7:0]) +
	( 9'sd 205) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22213) * $signed(input_fmap_235[7:0]) +
	( 16'sd 32435) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14225) * $signed(input_fmap_237[7:0]) +
	( 14'sd 4923) * $signed(input_fmap_238[7:0]) +
	( 15'sd 15447) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23286) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23747) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15163) * $signed(input_fmap_242[7:0]) +
	( 15'sd 9120) * $signed(input_fmap_243[7:0]) +
	( 16'sd 17246) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22943) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19121) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12468) * $signed(input_fmap_247[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_248[7:0]) +
	( 10'sd 480) * $signed(input_fmap_249[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_250[7:0]) +
	( 15'sd 8980) * $signed(input_fmap_251[7:0]) +
	( 16'sd 21987) * $signed(input_fmap_252[7:0]) +
	( 11'sd 851) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23216) * $signed(input_fmap_254[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_92;
assign conv_mac_92 = 
	( 16'sd 23848) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7896) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26580) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12832) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20955) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7643) * $signed(input_fmap_5[7:0]) +
	( 10'sd 295) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7813) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12949) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7194) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14453) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11951) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15596) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5103) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24719) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29388) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6964) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18532) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30239) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7361) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24763) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23561) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21115) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26791) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28154) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22877) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32120) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19632) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20318) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24345) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13864) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12677) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22906) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12544) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20404) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9426) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19630) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11375) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6777) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31336) * $signed(input_fmap_43[7:0]) +
	( 11'sd 587) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11030) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24564) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12043) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25445) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22951) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18552) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19831) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28788) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22657) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17695) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15354) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6914) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32682) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14691) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14325) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11687) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17982) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11807) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25249) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30461) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5950) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10241) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12930) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19168) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5614) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32299) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29700) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19872) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28828) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12074) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18459) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25196) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8891) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31809) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30562) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14712) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6757) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29195) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16965) * $signed(input_fmap_89[7:0]) +
	( 11'sd 844) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16940) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2696) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8095) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1760) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5557) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2197) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28954) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9905) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23620) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27492) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19666) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3447) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22425) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28995) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15846) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13331) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25039) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17517) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20994) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7621) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22989) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25303) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10279) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26629) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17894) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10274) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21722) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21438) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16458) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7961) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32125) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10385) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20860) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19356) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10051) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19597) * $signed(input_fmap_127[7:0]) +
	( 14'sd 6880) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19199) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6004) * $signed(input_fmap_130[7:0]) +
	( 15'sd 9336) * $signed(input_fmap_131[7:0]) +
	( 16'sd 27517) * $signed(input_fmap_132[7:0]) +
	( 4'sd 5) * $signed(input_fmap_133[7:0]) +
	( 16'sd 16444) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27610) * $signed(input_fmap_135[7:0]) +
	( 13'sd 3205) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11783) * $signed(input_fmap_137[7:0]) +
	( 16'sd 26684) * $signed(input_fmap_138[7:0]) +
	( 14'sd 5423) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15962) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19091) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31093) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31106) * $signed(input_fmap_144[7:0]) +
	( 15'sd 15098) * $signed(input_fmap_145[7:0]) +
	( 14'sd 4328) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13687) * $signed(input_fmap_147[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23134) * $signed(input_fmap_149[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_150[7:0]) +
	( 15'sd 9976) * $signed(input_fmap_151[7:0]) +
	( 16'sd 18826) * $signed(input_fmap_152[7:0]) +
	( 16'sd 21589) * $signed(input_fmap_153[7:0]) +
	( 13'sd 2842) * $signed(input_fmap_154[7:0]) +
	( 15'sd 8603) * $signed(input_fmap_155[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15921) * $signed(input_fmap_157[7:0]) +
	( 15'sd 12622) * $signed(input_fmap_158[7:0]) +
	( 16'sd 25557) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22952) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22552) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10371) * $signed(input_fmap_162[7:0]) +
	( 15'sd 11943) * $signed(input_fmap_163[7:0]) +
	( 16'sd 27763) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14708) * $signed(input_fmap_165[7:0]) +
	( 16'sd 24864) * $signed(input_fmap_166[7:0]) +
	( 16'sd 19526) * $signed(input_fmap_167[7:0]) +
	( 16'sd 27668) * $signed(input_fmap_168[7:0]) +
	( 13'sd 2446) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7835) * $signed(input_fmap_170[7:0]) +
	( 15'sd 8196) * $signed(input_fmap_171[7:0]) +
	( 14'sd 8154) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29684) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26451) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3948) * $signed(input_fmap_175[7:0]) +
	( 14'sd 5523) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6427) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17886) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15970) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23468) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19032) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12038) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31928) * $signed(input_fmap_184[7:0]) +
	( 15'sd 13244) * $signed(input_fmap_185[7:0]) +
	( 16'sd 32210) * $signed(input_fmap_186[7:0]) +
	( 11'sd 631) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13807) * $signed(input_fmap_188[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_189[7:0]) +
	( 16'sd 25961) * $signed(input_fmap_190[7:0]) +
	( 12'sd 1931) * $signed(input_fmap_191[7:0]) +
	( 14'sd 5726) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_193[7:0]) +
	( 16'sd 16804) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1100) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12148) * $signed(input_fmap_196[7:0]) +
	( 14'sd 4885) * $signed(input_fmap_197[7:0]) +
	( 16'sd 20182) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14120) * $signed(input_fmap_199[7:0]) +
	( 16'sd 27899) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27038) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31202) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19596) * $signed(input_fmap_204[7:0]) +
	( 16'sd 19734) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31861) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17792) * $signed(input_fmap_207[7:0]) +
	( 16'sd 21241) * $signed(input_fmap_208[7:0]) +
	( 14'sd 6904) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15489) * $signed(input_fmap_210[7:0]) +
	( 16'sd 21113) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14576) * $signed(input_fmap_212[7:0]) +
	( 11'sd 900) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30811) * $signed(input_fmap_214[7:0]) +
	( 15'sd 15853) * $signed(input_fmap_215[7:0]) +
	( 16'sd 31431) * $signed(input_fmap_216[7:0]) +
	( 11'sd 922) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8229) * $signed(input_fmap_218[7:0]) +
	( 14'sd 8047) * $signed(input_fmap_219[7:0]) +
	( 16'sd 23476) * $signed(input_fmap_220[7:0]) +
	( 13'sd 2978) * $signed(input_fmap_221[7:0]) +
	( 16'sd 27342) * $signed(input_fmap_222[7:0]) +
	( 15'sd 11227) * $signed(input_fmap_223[7:0]) +
	( 16'sd 26325) * $signed(input_fmap_224[7:0]) +
	( 16'sd 28839) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29346) * $signed(input_fmap_226[7:0]) +
	( 16'sd 21821) * $signed(input_fmap_227[7:0]) +
	( 15'sd 11870) * $signed(input_fmap_228[7:0]) +
	( 16'sd 19604) * $signed(input_fmap_229[7:0]) +
	( 16'sd 32643) * $signed(input_fmap_230[7:0]) +
	( 14'sd 4915) * $signed(input_fmap_231[7:0]) +
	( 14'sd 6083) * $signed(input_fmap_232[7:0]) +
	( 10'sd 387) * $signed(input_fmap_233[7:0]) +
	( 12'sd 1641) * $signed(input_fmap_234[7:0]) +
	( 16'sd 31182) * $signed(input_fmap_235[7:0]) +
	( 16'sd 29591) * $signed(input_fmap_236[7:0]) +
	( 15'sd 13736) * $signed(input_fmap_237[7:0]) +
	( 15'sd 9476) * $signed(input_fmap_238[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_239[7:0]) +
	( 14'sd 5165) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20934) * $signed(input_fmap_241[7:0]) +
	( 16'sd 22948) * $signed(input_fmap_242[7:0]) +
	( 15'sd 11539) * $signed(input_fmap_243[7:0]) +
	( 10'sd 488) * $signed(input_fmap_244[7:0]) +
	( 16'sd 25595) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9124) * $signed(input_fmap_246[7:0]) +
	( 16'sd 23174) * $signed(input_fmap_247[7:0]) +
	( 16'sd 28125) * $signed(input_fmap_248[7:0]) +
	( 15'sd 8680) * $signed(input_fmap_249[7:0]) +
	( 13'sd 2405) * $signed(input_fmap_250[7:0]) +
	( 16'sd 20318) * $signed(input_fmap_251[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_252[7:0]) +
	( 16'sd 31011) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5015) * $signed(input_fmap_254[7:0]) +
	( 15'sd 9592) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_93;
assign conv_mac_93 = 
	( 16'sd 27120) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11056) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17327) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8398) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28423) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4852) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5409) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18775) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25733) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5480) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6393) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25011) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8730) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17686) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5652) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6495) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5220) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23466) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6451) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13735) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31549) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9539) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25828) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24449) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6737) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28959) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18088) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29385) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32008) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10094) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31745) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14774) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6838) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16923) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25618) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29844) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3400) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26701) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29965) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4584) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9753) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24337) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27760) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26991) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24480) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31604) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17340) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1130) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13773) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15396) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7720) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25639) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12702) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25316) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14530) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3987) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3804) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28145) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30908) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18594) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31496) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32132) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10990) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15343) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17086) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15161) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30467) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16997) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21178) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31762) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5235) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10874) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30419) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11558) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23666) * $signed(input_fmap_82[7:0]) +
	( 11'sd 977) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19929) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1647) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17751) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3618) * $signed(input_fmap_88[7:0]) +
	( 11'sd 741) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21809) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30878) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9701) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25297) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4262) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1167) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19519) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13218) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12421) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2968) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9238) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13505) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22353) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8322) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3081) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21154) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24352) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7065) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15480) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6763) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32369) * $signed(input_fmap_112[7:0]) +
	( 15'sd 9494) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3924) * $signed(input_fmap_115[7:0]) +
	( 11'sd 514) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19483) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9362) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27093) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20071) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29681) * $signed(input_fmap_121[7:0]) +
	( 11'sd 863) * $signed(input_fmap_122[7:0]) +
	( 10'sd 388) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22738) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21892) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6386) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12621) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9287) * $signed(input_fmap_128[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_129[7:0]) +
	( 15'sd 8786) * $signed(input_fmap_130[7:0]) +
	( 15'sd 10658) * $signed(input_fmap_131[7:0]) +
	( 16'sd 17334) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11159) * $signed(input_fmap_133[7:0]) +
	( 16'sd 20322) * $signed(input_fmap_134[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_135[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11551) * $signed(input_fmap_137[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20286) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29004) * $signed(input_fmap_140[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_141[7:0]) +
	( 12'sd 2016) * $signed(input_fmap_142[7:0]) +
	( 14'sd 6709) * $signed(input_fmap_143[7:0]) +
	( 15'sd 16316) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23499) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19792) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27149) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6289) * $signed(input_fmap_148[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27159) * $signed(input_fmap_150[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_151[7:0]) +
	( 10'sd 444) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27719) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7219) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13357) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14162) * $signed(input_fmap_156[7:0]) +
	( 15'sd 10748) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4922) * $signed(input_fmap_158[7:0]) +
	( 15'sd 15662) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11880) * $signed(input_fmap_160[7:0]) +
	( 13'sd 2699) * $signed(input_fmap_161[7:0]) +
	( 15'sd 12085) * $signed(input_fmap_162[7:0]) +
	( 15'sd 10226) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19854) * $signed(input_fmap_164[7:0]) +
	( 11'sd 896) * $signed(input_fmap_165[7:0]) +
	( 12'sd 1613) * $signed(input_fmap_166[7:0]) +
	( 16'sd 28750) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17498) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6388) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14353) * $signed(input_fmap_170[7:0]) +
	( 16'sd 28355) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12747) * $signed(input_fmap_172[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_173[7:0]) +
	( 12'sd 1098) * $signed(input_fmap_174[7:0]) +
	( 16'sd 26348) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3768) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30399) * $signed(input_fmap_177[7:0]) +
	( 9'sd 227) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20258) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23429) * $signed(input_fmap_180[7:0]) +
	( 15'sd 10871) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19186) * $signed(input_fmap_182[7:0]) +
	( 15'sd 9806) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14413) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24122) * $signed(input_fmap_185[7:0]) +
	( 16'sd 20906) * $signed(input_fmap_186[7:0]) +
	( 16'sd 19473) * $signed(input_fmap_187[7:0]) +
	( 16'sd 18990) * $signed(input_fmap_188[7:0]) +
	( 15'sd 14183) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31789) * $signed(input_fmap_190[7:0]) +
	( 16'sd 22605) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19438) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15207) * $signed(input_fmap_193[7:0]) +
	( 16'sd 16384) * $signed(input_fmap_194[7:0]) +
	( 15'sd 8255) * $signed(input_fmap_195[7:0]) +
	( 16'sd 23684) * $signed(input_fmap_196[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_197[7:0]) +
	( 16'sd 20912) * $signed(input_fmap_198[7:0]) +
	( 15'sd 9909) * $signed(input_fmap_199[7:0]) +
	( 15'sd 9910) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16701) * $signed(input_fmap_201[7:0]) +
	( 14'sd 4836) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13560) * $signed(input_fmap_203[7:0]) +
	( 15'sd 9963) * $signed(input_fmap_204[7:0]) +
	( 14'sd 7717) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30328) * $signed(input_fmap_207[7:0]) +
	( 12'sd 1193) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7524) * $signed(input_fmap_209[7:0]) +
	( 16'sd 22611) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30700) * $signed(input_fmap_211[7:0]) +
	( 16'sd 20215) * $signed(input_fmap_212[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17002) * $signed(input_fmap_214[7:0]) +
	( 16'sd 27649) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20810) * $signed(input_fmap_216[7:0]) +
	( 16'sd 31160) * $signed(input_fmap_217[7:0]) +
	( 15'sd 12704) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21687) * $signed(input_fmap_219[7:0]) +
	( 11'sd 564) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_221[7:0]) +
	( 16'sd 31393) * $signed(input_fmap_222[7:0]) +
	( 15'sd 10797) * $signed(input_fmap_223[7:0]) +
	( 11'sd 976) * $signed(input_fmap_224[7:0]) +
	( 16'sd 16719) * $signed(input_fmap_225[7:0]) +
	( 16'sd 24376) * $signed(input_fmap_226[7:0]) +
	( 12'sd 1617) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25623) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3067) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29168) * $signed(input_fmap_230[7:0]) +
	( 16'sd 19274) * $signed(input_fmap_231[7:0]) +
	( 16'sd 21958) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14094) * $signed(input_fmap_233[7:0]) +
	( 16'sd 30388) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3491) * $signed(input_fmap_235[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20947) * $signed(input_fmap_237[7:0]) +
	( 7'sd 60) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12056) * $signed(input_fmap_239[7:0]) +
	( 11'sd 743) * $signed(input_fmap_240[7:0]) +
	( 16'sd 31803) * $signed(input_fmap_241[7:0]) +
	( 16'sd 20950) * $signed(input_fmap_242[7:0]) +
	( 16'sd 17196) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7933) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20668) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20563) * $signed(input_fmap_247[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_249[7:0]) +
	( 16'sd 28874) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_251[7:0]) +
	( 15'sd 14578) * $signed(input_fmap_252[7:0]) +
	( 14'sd 4967) * $signed(input_fmap_253[7:0]) +
	( 14'sd 6156) * $signed(input_fmap_254[7:0]) +
	( 16'sd 27998) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_94;
assign conv_mac_94 = 
	( 16'sd 16766) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15274) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16541) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21709) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14042) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10304) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25255) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12497) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2177) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23579) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23304) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25603) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7332) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4870) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17072) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18020) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_18[7:0]) +
	( 8'sd 79) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20753) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13885) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5787) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2300) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23356) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30186) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27203) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10098) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31216) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11873) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14977) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18670) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20845) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12325) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10073) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25664) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10627) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26863) * $signed(input_fmap_39[7:0]) +
	( 15'sd 16317) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30697) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7890) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6050) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13756) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29619) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13101) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21407) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10749) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4757) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3214) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23201) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9715) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8401) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10515) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4141) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26480) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9126) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23651) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6656) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7448) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20713) * $signed(input_fmap_65[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29891) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7799) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16826) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18569) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7436) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31359) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19518) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20312) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30766) * $signed(input_fmap_75[7:0]) +
	( 9'sd 185) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3452) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24791) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31713) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22647) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26933) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21925) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30097) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30757) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23086) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6378) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26032) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16182) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7535) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31533) * $signed(input_fmap_90[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17422) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26692) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27018) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12947) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17306) * $signed(input_fmap_96[7:0]) +
	( 7'sd 55) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15979) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22029) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7500) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13980) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27107) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1323) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28227) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15161) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24893) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15957) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25502) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16233) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23204) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7137) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5525) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7386) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6903) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28186) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30845) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24536) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20999) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11170) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7041) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3501) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9181) * $signed(input_fmap_125[7:0]) +
	( 13'sd 4062) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23509) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31774) * $signed(input_fmap_129[7:0]) +
	( 14'sd 7608) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18663) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10433) * $signed(input_fmap_133[7:0]) +
	( 11'sd 898) * $signed(input_fmap_134[7:0]) +
	( 15'sd 12831) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31586) * $signed(input_fmap_136[7:0]) +
	( 13'sd 2614) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27603) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11130) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17013) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13241) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28420) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20770) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4808) * $signed(input_fmap_144[7:0]) +
	( 15'sd 13255) * $signed(input_fmap_145[7:0]) +
	( 15'sd 10129) * $signed(input_fmap_146[7:0]) +
	( 16'sd 23799) * $signed(input_fmap_147[7:0]) +
	( 15'sd 14462) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27736) * $signed(input_fmap_149[7:0]) +
	( 13'sd 2334) * $signed(input_fmap_150[7:0]) +
	( 15'sd 9190) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22103) * $signed(input_fmap_152[7:0]) +
	( 16'sd 22659) * $signed(input_fmap_153[7:0]) +
	( 15'sd 15523) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25257) * $signed(input_fmap_156[7:0]) +
	( 14'sd 7263) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8813) * $signed(input_fmap_158[7:0]) +
	( 16'sd 30451) * $signed(input_fmap_159[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_160[7:0]) +
	( 15'sd 13636) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26780) * $signed(input_fmap_162[7:0]) +
	( 16'sd 21523) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13222) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12442) * $signed(input_fmap_165[7:0]) +
	( 15'sd 16350) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7364) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6737) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28059) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12044) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31907) * $signed(input_fmap_172[7:0]) +
	( 16'sd 32747) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15241) * $signed(input_fmap_175[7:0]) +
	( 15'sd 16151) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1627) * $signed(input_fmap_177[7:0]) +
	( 16'sd 30484) * $signed(input_fmap_178[7:0]) +
	( 15'sd 10861) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23267) * $signed(input_fmap_180[7:0]) +
	( 14'sd 5463) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12313) * $signed(input_fmap_182[7:0]) +
	( 16'sd 16783) * $signed(input_fmap_183[7:0]) +
	( 15'sd 15421) * $signed(input_fmap_184[7:0]) +
	( 15'sd 16151) * $signed(input_fmap_185[7:0]) +
	( 16'sd 32462) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11967) * $signed(input_fmap_187[7:0]) +
	( 15'sd 11288) * $signed(input_fmap_188[7:0]) +
	( 16'sd 21720) * $signed(input_fmap_189[7:0]) +
	( 16'sd 26994) * $signed(input_fmap_190[7:0]) +
	( 15'sd 9619) * $signed(input_fmap_191[7:0]) +
	( 16'sd 25637) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6725) * $signed(input_fmap_193[7:0]) +
	( 15'sd 15890) * $signed(input_fmap_194[7:0]) +
	( 13'sd 3513) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7548) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24075) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_198[7:0]) +
	( 16'sd 19028) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26147) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1309) * $signed(input_fmap_201[7:0]) +
	( 16'sd 16723) * $signed(input_fmap_202[7:0]) +
	( 16'sd 18134) * $signed(input_fmap_203[7:0]) +
	( 16'sd 24567) * $signed(input_fmap_204[7:0]) +
	( 14'sd 7548) * $signed(input_fmap_205[7:0]) +
	( 16'sd 26797) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28232) * $signed(input_fmap_207[7:0]) +
	( 11'sd 625) * $signed(input_fmap_208[7:0]) +
	( 15'sd 9427) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4243) * $signed(input_fmap_210[7:0]) +
	( 13'sd 2082) * $signed(input_fmap_211[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18083) * $signed(input_fmap_214[7:0]) +
	( 15'sd 15738) * $signed(input_fmap_215[7:0]) +
	( 13'sd 4066) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24369) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22130) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12796) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24030) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19322) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9986) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19932) * $signed(input_fmap_224[7:0]) +
	( 15'sd 10734) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31360) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3756) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25815) * $signed(input_fmap_228[7:0]) +
	( 14'sd 7745) * $signed(input_fmap_229[7:0]) +
	( 11'sd 696) * $signed(input_fmap_230[7:0]) +
	( 16'sd 21469) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_232[7:0]) +
	( 14'sd 7700) * $signed(input_fmap_233[7:0]) +
	( 16'sd 17889) * $signed(input_fmap_234[7:0]) +
	( 14'sd 6347) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25749) * $signed(input_fmap_236[7:0]) +
	( 12'sd 1082) * $signed(input_fmap_237[7:0]) +
	( 11'sd 545) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9775) * $signed(input_fmap_239[7:0]) +
	( 16'sd 30973) * $signed(input_fmap_240[7:0]) +
	( 16'sd 28997) * $signed(input_fmap_241[7:0]) +
	( 16'sd 18728) * $signed(input_fmap_242[7:0]) +
	( 11'sd 745) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2121) * $signed(input_fmap_244[7:0]) +
	( 14'sd 4698) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17269) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_247[7:0]) +
	( 16'sd 28655) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14993) * $signed(input_fmap_249[7:0]) +
	( 16'sd 27013) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19306) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20179) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24864) * $signed(input_fmap_253[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_254[7:0]) +
	( 16'sd 28609) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_95;
assign conv_mac_95 = 
	( 16'sd 24462) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9784) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20957) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29578) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11277) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6494) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27189) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25294) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4767) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11726) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26461) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29152) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20569) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24118) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6745) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13195) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16641) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5860) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25845) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27836) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10636) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13693) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12814) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19761) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7838) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16961) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23460) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32529) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16514) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13447) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28079) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11311) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18248) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15777) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17208) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4701) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24229) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18523) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31774) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7600) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19089) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6344) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28060) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18798) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12628) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27221) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24401) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12461) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29829) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13459) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22343) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32426) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22743) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32367) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30180) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23993) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6028) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17648) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1228) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19864) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7961) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12099) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3275) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27552) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16323) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6319) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31906) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16815) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25765) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9633) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7678) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22550) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19235) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13356) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3896) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1527) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_85[7:0]) +
	( 16'sd 27644) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3552) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11334) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14063) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11533) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1419) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4147) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16641) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1298) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10176) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19970) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2224) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24242) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2711) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3133) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5541) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31592) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17121) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1025) * $signed(input_fmap_106[7:0]) +
	( 3'sd 2) * $signed(input_fmap_107[7:0]) +
	( 16'sd 21083) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16084) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30392) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7921) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15199) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10830) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6113) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13100) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27722) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6028) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3287) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10789) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10692) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3029) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1126) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1602) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2592) * $signed(input_fmap_127[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7752) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19479) * $signed(input_fmap_130[7:0]) +
	( 16'sd 22573) * $signed(input_fmap_131[7:0]) +
	( 16'sd 19343) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29250) * $signed(input_fmap_133[7:0]) +
	( 16'sd 17685) * $signed(input_fmap_134[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_135[7:0]) +
	( 15'sd 11458) * $signed(input_fmap_136[7:0]) +
	( 16'sd 31006) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10574) * $signed(input_fmap_138[7:0]) +
	( 16'sd 25129) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1451) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20649) * $signed(input_fmap_141[7:0]) +
	( 16'sd 17327) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23531) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13715) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25309) * $signed(input_fmap_145[7:0]) +
	( 13'sd 2802) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21486) * $signed(input_fmap_147[7:0]) +
	( 13'sd 2569) * $signed(input_fmap_148[7:0]) +
	( 16'sd 20366) * $signed(input_fmap_149[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_150[7:0]) +
	( 16'sd 26465) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29106) * $signed(input_fmap_152[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7037) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19683) * $signed(input_fmap_155[7:0]) +
	( 14'sd 6052) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6913) * $signed(input_fmap_157[7:0]) +
	( 16'sd 26386) * $signed(input_fmap_158[7:0]) +
	( 15'sd 13049) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_160[7:0]) +
	( 15'sd 12943) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4965) * $signed(input_fmap_162[7:0]) +
	( 15'sd 12953) * $signed(input_fmap_163[7:0]) +
	( 16'sd 32035) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19095) * $signed(input_fmap_165[7:0]) +
	( 15'sd 16147) * $signed(input_fmap_166[7:0]) +
	( 15'sd 14891) * $signed(input_fmap_167[7:0]) +
	( 16'sd 24244) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11575) * $signed(input_fmap_170[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_171[7:0]) +
	( 16'sd 20598) * $signed(input_fmap_172[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_173[7:0]) +
	( 12'sd 1212) * $signed(input_fmap_174[7:0]) +
	( 16'sd 19337) * $signed(input_fmap_175[7:0]) +
	( 16'sd 24852) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31025) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31610) * $signed(input_fmap_178[7:0]) +
	( 16'sd 16599) * $signed(input_fmap_179[7:0]) +
	( 16'sd 20590) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18726) * $signed(input_fmap_181[7:0]) +
	( 16'sd 20784) * $signed(input_fmap_182[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13659) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13994) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18513) * $signed(input_fmap_187[7:0]) +
	( 16'sd 20753) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17847) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9511) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26665) * $signed(input_fmap_191[7:0]) +
	( 15'sd 10121) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19527) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18662) * $signed(input_fmap_194[7:0]) +
	( 16'sd 16634) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19416) * $signed(input_fmap_196[7:0]) +
	( 14'sd 7120) * $signed(input_fmap_197[7:0]) +
	( 16'sd 25229) * $signed(input_fmap_198[7:0]) +
	( 15'sd 8853) * $signed(input_fmap_199[7:0]) +
	( 12'sd 1348) * $signed(input_fmap_200[7:0]) +
	( 16'sd 25422) * $signed(input_fmap_201[7:0]) +
	( 15'sd 16179) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5885) * $signed(input_fmap_203[7:0]) +
	( 16'sd 27813) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30522) * $signed(input_fmap_205[7:0]) +
	( 16'sd 17947) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29798) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30996) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13196) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18562) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6920) * $signed(input_fmap_211[7:0]) +
	( 14'sd 5000) * $signed(input_fmap_212[7:0]) +
	( 14'sd 7268) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20592) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5224) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25613) * $signed(input_fmap_217[7:0]) +
	( 12'sd 1923) * $signed(input_fmap_218[7:0]) +
	( 14'sd 6092) * $signed(input_fmap_219[7:0]) +
	( 14'sd 5146) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19481) * $signed(input_fmap_221[7:0]) +
	( 16'sd 23503) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15934) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2179) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27313) * $signed(input_fmap_226[7:0]) +
	( 16'sd 21534) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2360) * $signed(input_fmap_228[7:0]) +
	( 15'sd 15233) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27863) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28422) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8327) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5749) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23547) * $signed(input_fmap_234[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_235[7:0]) +
	( 16'sd 16455) * $signed(input_fmap_236[7:0]) +
	( 16'sd 25886) * $signed(input_fmap_237[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18307) * $signed(input_fmap_240[7:0]) +
	( 15'sd 16088) * $signed(input_fmap_241[7:0]) +
	( 13'sd 3719) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31765) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6420) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22741) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30607) * $signed(input_fmap_247[7:0]) +
	( 16'sd 22601) * $signed(input_fmap_248[7:0]) +
	( 16'sd 19345) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7286) * $signed(input_fmap_250[7:0]) +
	( 15'sd 9373) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5635) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6992) * $signed(input_fmap_253[7:0]) +
	( 16'sd 28327) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14553) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_96;
assign conv_mac_96 = 
	( 15'sd 12711) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21616) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10900) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3520) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11466) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5339) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7087) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21193) * $signed(input_fmap_9[7:0]) +
	( 15'sd 13883) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25617) * $signed(input_fmap_11[7:0]) +
	( 12'sd 2037) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20850) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16784) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4866) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1153) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19068) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16853) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29573) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26123) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15109) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6795) * $signed(input_fmap_24[7:0]) +
	( 8'sd 95) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30633) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28992) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18354) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9172) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12928) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21758) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1862) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8996) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16247) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25213) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20224) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24926) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6360) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30603) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7183) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7869) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24748) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21912) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17563) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11954) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10047) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8574) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6049) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1262) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16623) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21270) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28892) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32034) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22346) * $signed(input_fmap_60[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22984) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15641) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11504) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2973) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20469) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7386) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16743) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21091) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25644) * $signed(input_fmap_71[7:0]) +
	( 13'sd 4090) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2257) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6107) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23954) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3649) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23214) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32554) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21377) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27302) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31175) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8392) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7399) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19970) * $signed(input_fmap_85[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3852) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14983) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25628) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23254) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12441) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21235) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2297) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4321) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22384) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10458) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7227) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18281) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4570) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10498) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30558) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14354) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14636) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27623) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23092) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15123) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30007) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21328) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30792) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24454) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2651) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12373) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17263) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7357) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27699) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12686) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15307) * $signed(input_fmap_121[7:0]) +
	( 11'sd 589) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7074) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3654) * $signed(input_fmap_124[7:0]) +
	( 14'sd 6392) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18758) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21755) * $signed(input_fmap_127[7:0]) +
	( 16'sd 26270) * $signed(input_fmap_128[7:0]) +
	( 14'sd 6542) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12736) * $signed(input_fmap_130[7:0]) +
	( 16'sd 28726) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25059) * $signed(input_fmap_132[7:0]) +
	( 14'sd 6254) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_134[7:0]) +
	( 15'sd 15979) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15751) * $signed(input_fmap_136[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_137[7:0]) +
	( 16'sd 18489) * $signed(input_fmap_138[7:0]) +
	( 16'sd 32395) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1164) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_141[7:0]) +
	( 16'sd 29508) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4527) * $signed(input_fmap_143[7:0]) +
	( 15'sd 10029) * $signed(input_fmap_144[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7172) * $signed(input_fmap_146[7:0]) +
	( 16'sd 31633) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28164) * $signed(input_fmap_148[7:0]) +
	( 16'sd 19648) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5855) * $signed(input_fmap_150[7:0]) +
	( 15'sd 11901) * $signed(input_fmap_151[7:0]) +
	( 16'sd 27156) * $signed(input_fmap_152[7:0]) +
	( 14'sd 5783) * $signed(input_fmap_153[7:0]) +
	( 16'sd 26660) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7318) * $signed(input_fmap_155[7:0]) +
	( 16'sd 19197) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_157[7:0]) +
	( 15'sd 13625) * $signed(input_fmap_158[7:0]) +
	( 16'sd 23831) * $signed(input_fmap_159[7:0]) +
	( 12'sd 1517) * $signed(input_fmap_160[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10471) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28519) * $signed(input_fmap_163[7:0]) +
	( 16'sd 27649) * $signed(input_fmap_164[7:0]) +
	( 16'sd 17972) * $signed(input_fmap_165[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_166[7:0]) +
	( 16'sd 16564) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4732) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6552) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5088) * $signed(input_fmap_170[7:0]) +
	( 15'sd 10852) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31441) * $signed(input_fmap_172[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11269) * $signed(input_fmap_174[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7839) * $signed(input_fmap_176[7:0]) +
	( 15'sd 13989) * $signed(input_fmap_177[7:0]) +
	( 14'sd 4388) * $signed(input_fmap_178[7:0]) +
	( 12'sd 1458) * $signed(input_fmap_179[7:0]) +
	( 16'sd 20587) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15992) * $signed(input_fmap_181[7:0]) +
	( 8'sd 80) * $signed(input_fmap_182[7:0]) +
	( 15'sd 10336) * $signed(input_fmap_183[7:0]) +
	( 15'sd 12753) * $signed(input_fmap_184[7:0]) +
	( 16'sd 23665) * $signed(input_fmap_185[7:0]) +
	( 16'sd 30845) * $signed(input_fmap_186[7:0]) +
	( 14'sd 7438) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12302) * $signed(input_fmap_188[7:0]) +
	( 16'sd 29403) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27680) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5225) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12343) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19696) * $signed(input_fmap_193[7:0]) +
	( 14'sd 5771) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29040) * $signed(input_fmap_195[7:0]) +
	( 16'sd 28226) * $signed(input_fmap_196[7:0]) +
	( 15'sd 12283) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5565) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12352) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15672) * $signed(input_fmap_200[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19481) * $signed(input_fmap_202[7:0]) +
	( 16'sd 17495) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11638) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11321) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20537) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_208[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_209[7:0]) +
	( 16'sd 32307) * $signed(input_fmap_210[7:0]) +
	( 16'sd 32616) * $signed(input_fmap_211[7:0]) +
	( 15'sd 8454) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9156) * $signed(input_fmap_213[7:0]) +
	( 16'sd 21261) * $signed(input_fmap_214[7:0]) +
	( 16'sd 18388) * $signed(input_fmap_215[7:0]) +
	( 13'sd 3917) * $signed(input_fmap_216[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10052) * $signed(input_fmap_218[7:0]) +
	( 16'sd 32056) * $signed(input_fmap_219[7:0]) +
	( 16'sd 27509) * $signed(input_fmap_220[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_221[7:0]) +
	( 14'sd 4982) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12546) * $signed(input_fmap_223[7:0]) +
	( 15'sd 9412) * $signed(input_fmap_224[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32657) * $signed(input_fmap_226[7:0]) +
	( 15'sd 12811) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8614) * $signed(input_fmap_228[7:0]) +
	( 16'sd 32039) * $signed(input_fmap_229[7:0]) +
	( 16'sd 22634) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10629) * $signed(input_fmap_231[7:0]) +
	( 14'sd 6382) * $signed(input_fmap_232[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15845) * $signed(input_fmap_234[7:0]) +
	( 15'sd 8890) * $signed(input_fmap_235[7:0]) +
	( 15'sd 16104) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2426) * $signed(input_fmap_237[7:0]) +
	( 12'sd 1889) * $signed(input_fmap_238[7:0]) +
	( 14'sd 7077) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9708) * $signed(input_fmap_240[7:0]) +
	( 13'sd 2836) * $signed(input_fmap_241[7:0]) +
	( 16'sd 32419) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13113) * $signed(input_fmap_243[7:0]) +
	( 16'sd 25559) * $signed(input_fmap_244[7:0]) +
	( 16'sd 27283) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20013) * $signed(input_fmap_247[7:0]) +
	( 15'sd 8816) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9732) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9578) * $signed(input_fmap_250[7:0]) +
	( 12'sd 1898) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2158) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2431) * $signed(input_fmap_253[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_254[7:0]) +
	( 14'sd 4567) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_97;
assign conv_mac_97 = 
	( 14'sd 4462) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23778) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24886) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14439) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25833) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14455) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12373) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4149) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17009) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6810) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25309) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13844) * $signed(input_fmap_12[7:0]) +
	( 10'sd 318) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13387) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27473) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16181) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13860) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4424) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18715) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15466) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15721) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9140) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26370) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19928) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16503) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6319) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4314) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17836) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19773) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20377) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1269) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23161) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21870) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21640) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6638) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11448) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3329) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21519) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12193) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8907) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4139) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12528) * $signed(input_fmap_45[7:0]) +
	( 16'sd 32674) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22824) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20383) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26952) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5876) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1231) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20856) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4155) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21252) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3704) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6875) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29828) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29123) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32373) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9723) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27016) * $signed(input_fmap_62[7:0]) +
	( 11'sd 898) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9594) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29075) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22798) * $signed(input_fmap_66[7:0]) +
	( 11'sd 711) * $signed(input_fmap_67[7:0]) +
	( 11'sd 982) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13854) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6592) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16272) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7397) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31736) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6479) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23687) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2136) * $signed(input_fmap_78[7:0]) +
	( 15'sd 15744) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32124) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32123) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32023) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21521) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25591) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1635) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20415) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13820) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13074) * $signed(input_fmap_90[7:0]) +
	( 13'sd 2515) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16481) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28147) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31584) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15382) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14292) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14840) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16661) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12467) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21511) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2601) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22526) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28536) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8515) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32569) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11674) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8719) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11861) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25886) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20249) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14916) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25102) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2676) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2116) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12024) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27673) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2328) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18738) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9238) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23708) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11003) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1397) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27133) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1553) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29784) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29531) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8480) * $signed(input_fmap_128[7:0]) +
	( 15'sd 11135) * $signed(input_fmap_129[7:0]) +
	( 16'sd 28031) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31117) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14281) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12888) * $signed(input_fmap_133[7:0]) +
	( 13'sd 4037) * $signed(input_fmap_134[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15290) * $signed(input_fmap_136[7:0]) +
	( 16'sd 16558) * $signed(input_fmap_137[7:0]) +
	( 16'sd 23512) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8611) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28053) * $signed(input_fmap_140[7:0]) +
	( 16'sd 21803) * $signed(input_fmap_141[7:0]) +
	( 13'sd 2245) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_143[7:0]) +
	( 16'sd 24755) * $signed(input_fmap_144[7:0]) +
	( 15'sd 10871) * $signed(input_fmap_145[7:0]) +
	( 13'sd 2916) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21245) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11265) * $signed(input_fmap_148[7:0]) +
	( 16'sd 26587) * $signed(input_fmap_149[7:0]) +
	( 16'sd 17724) * $signed(input_fmap_150[7:0]) +
	( 15'sd 10250) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6545) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2177) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5907) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13546) * $signed(input_fmap_156[7:0]) +
	( 13'sd 2065) * $signed(input_fmap_157[7:0]) +
	( 11'sd 581) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21848) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5853) * $signed(input_fmap_160[7:0]) +
	( 16'sd 29848) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27502) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15666) * $signed(input_fmap_163[7:0]) +
	( 15'sd 16219) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11910) * $signed(input_fmap_165[7:0]) +
	( 10'sd 492) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26346) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5395) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20619) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9198) * $signed(input_fmap_170[7:0]) +
	( 16'sd 23068) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19694) * $signed(input_fmap_172[7:0]) +
	( 14'sd 7357) * $signed(input_fmap_173[7:0]) +
	( 14'sd 5818) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15139) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3236) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2364) * $signed(input_fmap_177[7:0]) +
	( 14'sd 4553) * $signed(input_fmap_178[7:0]) +
	( 14'sd 4113) * $signed(input_fmap_179[7:0]) +
	( 16'sd 19741) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3842) * $signed(input_fmap_181[7:0]) +
	( 16'sd 32605) * $signed(input_fmap_182[7:0]) +
	( 16'sd 22974) * $signed(input_fmap_183[7:0]) +
	( 15'sd 16036) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13557) * $signed(input_fmap_186[7:0]) +
	( 16'sd 17281) * $signed(input_fmap_187[7:0]) +
	( 15'sd 10391) * $signed(input_fmap_188[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_189[7:0]) +
	( 16'sd 23382) * $signed(input_fmap_190[7:0]) +
	( 16'sd 21595) * $signed(input_fmap_191[7:0]) +
	( 16'sd 32355) * $signed(input_fmap_192[7:0]) +
	( 14'sd 7128) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14466) * $signed(input_fmap_194[7:0]) +
	( 15'sd 9161) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11298) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31606) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29174) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16014) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26206) * $signed(input_fmap_200[7:0]) +
	( 16'sd 24659) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21011) * $signed(input_fmap_202[7:0]) +
	( 16'sd 27035) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15789) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29323) * $signed(input_fmap_205[7:0]) +
	( 12'sd 2001) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18780) * $signed(input_fmap_207[7:0]) +
	( 15'sd 14713) * $signed(input_fmap_208[7:0]) +
	( 15'sd 8371) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30122) * $signed(input_fmap_210[7:0]) +
	( 13'sd 2622) * $signed(input_fmap_211[7:0]) +
	( 16'sd 31760) * $signed(input_fmap_212[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_213[7:0]) +
	( 16'sd 27722) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23025) * $signed(input_fmap_215[7:0]) +
	( 16'sd 25953) * $signed(input_fmap_216[7:0]) +
	( 13'sd 2789) * $signed(input_fmap_217[7:0]) +
	( 16'sd 27311) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28107) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13700) * $signed(input_fmap_221[7:0]) +
	( 15'sd 11819) * $signed(input_fmap_222[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27631) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10056) * $signed(input_fmap_226[7:0]) +
	( 16'sd 32670) * $signed(input_fmap_227[7:0]) +
	( 14'sd 7191) * $signed(input_fmap_228[7:0]) +
	( 16'sd 28306) * $signed(input_fmap_229[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_230[7:0]) +
	( 15'sd 11027) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3898) * $signed(input_fmap_233[7:0]) +
	( 16'sd 24217) * $signed(input_fmap_234[7:0]) +
	( 14'sd 8182) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25234) * $signed(input_fmap_236[7:0]) +
	( 16'sd 17024) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23937) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21070) * $signed(input_fmap_239[7:0]) +
	( 16'sd 32367) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15409) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29922) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13310) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12802) * $signed(input_fmap_245[7:0]) +
	( 16'sd 26875) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8945) * $signed(input_fmap_247[7:0]) +
	( 14'sd 5381) * $signed(input_fmap_248[7:0]) +
	( 14'sd 6916) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25677) * $signed(input_fmap_250[7:0]) +
	( 15'sd 9942) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12767) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25188) * $signed(input_fmap_253[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_254[7:0]) +
	( 16'sd 21466) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_98;
assign conv_mac_98 = 
	( 15'sd 15014) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17148) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27079) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8325) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12020) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20318) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23036) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9293) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26049) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8414) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4359) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4526) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23225) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30442) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12431) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31302) * $signed(input_fmap_16[7:0]) +
	( 16'sd 24636) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27814) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1821) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26990) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32230) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19106) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24977) * $signed(input_fmap_23[7:0]) +
	( 14'sd 6764) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4978) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8879) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21030) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4247) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3187) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1923) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5387) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10143) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14262) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15473) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25511) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1690) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26340) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12274) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18237) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12706) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31846) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5056) * $signed(input_fmap_46[7:0]) +
	( 6'sd 29) * $signed(input_fmap_47[7:0]) +
	( 16'sd 16555) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10049) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7518) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25831) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8445) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17639) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16316) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27663) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19669) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23232) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6187) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14894) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30207) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9089) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2295) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30248) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15009) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12086) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7255) * $signed(input_fmap_67[7:0]) +
	( 12'sd 2040) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21387) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11213) * $signed(input_fmap_70[7:0]) +
	( 15'sd 13552) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30809) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9561) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3741) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25832) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8142) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10090) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2964) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32736) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23329) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20580) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27610) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6517) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21984) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28952) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29826) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24235) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29748) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13686) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14769) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1418) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29021) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11716) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6720) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14059) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25075) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11579) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8786) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4828) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27993) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30014) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7385) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30877) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18394) * $signed(input_fmap_110[7:0]) +
	( 9'sd 166) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2515) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19339) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19677) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5953) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25291) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5165) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15900) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25851) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2881) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23053) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29089) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19545) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23374) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11039) * $signed(input_fmap_126[7:0]) +
	( 15'sd 14914) * $signed(input_fmap_127[7:0]) +
	( 16'sd 20218) * $signed(input_fmap_128[7:0]) +
	( 14'sd 4189) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18786) * $signed(input_fmap_130[7:0]) +
	( 16'sd 21357) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25995) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21171) * $signed(input_fmap_133[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10312) * $signed(input_fmap_135[7:0]) +
	( 16'sd 29477) * $signed(input_fmap_136[7:0]) +
	( 12'sd 1476) * $signed(input_fmap_137[7:0]) +
	( 15'sd 8628) * $signed(input_fmap_138[7:0]) +
	( 16'sd 23005) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29919) * $signed(input_fmap_140[7:0]) +
	( 13'sd 4058) * $signed(input_fmap_141[7:0]) +
	( 15'sd 12133) * $signed(input_fmap_142[7:0]) +
	( 16'sd 24472) * $signed(input_fmap_143[7:0]) +
	( 16'sd 27867) * $signed(input_fmap_144[7:0]) +
	( 15'sd 12680) * $signed(input_fmap_145[7:0]) +
	( 16'sd 23721) * $signed(input_fmap_146[7:0]) +
	( 16'sd 20279) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17774) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25835) * $signed(input_fmap_149[7:0]) +
	( 16'sd 26670) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28560) * $signed(input_fmap_151[7:0]) +
	( 14'sd 5094) * $signed(input_fmap_152[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_153[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_154[7:0]) +
	( 15'sd 9907) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13703) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11040) * $signed(input_fmap_157[7:0]) +
	( 16'sd 19436) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20038) * $signed(input_fmap_159[7:0]) +
	( 16'sd 20945) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4487) * $signed(input_fmap_161[7:0]) +
	( 15'sd 12779) * $signed(input_fmap_162[7:0]) +
	( 15'sd 9478) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9751) * $signed(input_fmap_164[7:0]) +
	( 16'sd 20619) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19356) * $signed(input_fmap_166[7:0]) +
	( 16'sd 32053) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26703) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21904) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31289) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15545) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_172[7:0]) +
	( 16'sd 20837) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_174[7:0]) +
	( 16'sd 18481) * $signed(input_fmap_175[7:0]) +
	( 16'sd 26526) * $signed(input_fmap_176[7:0]) +
	( 15'sd 10243) * $signed(input_fmap_177[7:0]) +
	( 13'sd 3995) * $signed(input_fmap_178[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23594) * $signed(input_fmap_180[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29406) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12383) * $signed(input_fmap_183[7:0]) +
	( 14'sd 7375) * $signed(input_fmap_184[7:0]) +
	( 16'sd 16888) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12405) * $signed(input_fmap_186[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13479) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17692) * $signed(input_fmap_189[7:0]) +
	( 12'sd 1097) * $signed(input_fmap_190[7:0]) +
	( 16'sd 22897) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14136) * $signed(input_fmap_192[7:0]) +
	( 14'sd 7149) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_194[7:0]) +
	( 15'sd 10454) * $signed(input_fmap_195[7:0]) +
	( 15'sd 10025) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14875) * $signed(input_fmap_197[7:0]) +
	( 16'sd 17431) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1380) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18668) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12033) * $signed(input_fmap_201[7:0]) +
	( 16'sd 22820) * $signed(input_fmap_202[7:0]) +
	( 15'sd 15832) * $signed(input_fmap_203[7:0]) +
	( 16'sd 25616) * $signed(input_fmap_204[7:0]) +
	( 16'sd 21360) * $signed(input_fmap_205[7:0]) +
	( 16'sd 32090) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29129) * $signed(input_fmap_207[7:0]) +
	( 15'sd 14888) * $signed(input_fmap_208[7:0]) +
	( 13'sd 2537) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23362) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10318) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24130) * $signed(input_fmap_212[7:0]) +
	( 16'sd 25026) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14554) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6952) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11519) * $signed(input_fmap_216[7:0]) +
	( 15'sd 12320) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31519) * $signed(input_fmap_218[7:0]) +
	( 14'sd 7686) * $signed(input_fmap_219[7:0]) +
	( 14'sd 6871) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13764) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18578) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28505) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7459) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26555) * $signed(input_fmap_225[7:0]) +
	( 11'sd 718) * $signed(input_fmap_226[7:0]) +
	( 16'sd 21723) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1146) * $signed(input_fmap_228[7:0]) +
	( 16'sd 31533) * $signed(input_fmap_229[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15224) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24961) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12641) * $signed(input_fmap_235[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_236[7:0]) +
	( 13'sd 3196) * $signed(input_fmap_237[7:0]) +
	( 11'sd 774) * $signed(input_fmap_238[7:0]) +
	( 16'sd 29599) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9726) * $signed(input_fmap_240[7:0]) +
	( 16'sd 19566) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11046) * $signed(input_fmap_242[7:0]) +
	( 16'sd 16463) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_244[7:0]) +
	( 16'sd 23341) * $signed(input_fmap_245[7:0]) +
	( 16'sd 21418) * $signed(input_fmap_246[7:0]) +
	( 13'sd 2607) * $signed(input_fmap_247[7:0]) +
	( 16'sd 28921) * $signed(input_fmap_248[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_249[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18338) * $signed(input_fmap_251[7:0]) +
	( 15'sd 9989) * $signed(input_fmap_252[7:0]) +
	( 16'sd 18373) * $signed(input_fmap_253[7:0]) +
	( 16'sd 28965) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10893) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_99;
assign conv_mac_99 = 
	( 14'sd 4111) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4749) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2868) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5059) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14773) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29802) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9434) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17861) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27361) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26829) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11320) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6779) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27868) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5451) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25880) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31563) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2441) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2786) * $signed(input_fmap_22[7:0]) +
	( 11'sd 578) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21571) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16767) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11662) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26638) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13459) * $signed(input_fmap_28[7:0]) +
	( 10'sd 361) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27720) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_33[7:0]) +
	( 7'sd 50) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26969) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12784) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19429) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7471) * $signed(input_fmap_38[7:0]) +
	( 10'sd 340) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5447) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9581) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9545) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12036) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2974) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26931) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17773) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26982) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10509) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21225) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4811) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6433) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3520) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25006) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16367) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17707) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19500) * $signed(input_fmap_63[7:0]) +
	( 9'sd 209) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1240) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21163) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19740) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18095) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26078) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16499) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17825) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20238) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24910) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29680) * $signed(input_fmap_74[7:0]) +
	( 13'sd 4071) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21746) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23486) * $signed(input_fmap_77[7:0]) +
	( 10'sd 481) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11864) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24635) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24563) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3137) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30045) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10549) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1270) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10447) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5498) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7874) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24262) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32494) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21819) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10064) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5777) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13302) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18595) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4844) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3073) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17634) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29880) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25105) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30902) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23824) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19458) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23323) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4567) * $signed(input_fmap_109[7:0]) +
	( 11'sd 582) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25967) * $signed(input_fmap_111[7:0]) +
	( 8'sd 87) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28467) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23931) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10640) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2753) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8874) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7071) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19639) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26855) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19715) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8793) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16462) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17122) * $signed(input_fmap_128[7:0]) +
	( 16'sd 20753) * $signed(input_fmap_129[7:0]) +
	( 16'sd 29039) * $signed(input_fmap_130[7:0]) +
	( 13'sd 2640) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1354) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10529) * $signed(input_fmap_133[7:0]) +
	( 14'sd 7362) * $signed(input_fmap_134[7:0]) +
	( 15'sd 12292) * $signed(input_fmap_135[7:0]) +
	( 14'sd 6078) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24944) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11926) * $signed(input_fmap_138[7:0]) +
	( 14'sd 5226) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26185) * $signed(input_fmap_140[7:0]) +
	( 15'sd 14561) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31042) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18317) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17227) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1603) * $signed(input_fmap_146[7:0]) +
	( 16'sd 16946) * $signed(input_fmap_147[7:0]) +
	( 15'sd 13360) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31598) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6063) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16493) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14343) * $signed(input_fmap_153[7:0]) +
	( 15'sd 14436) * $signed(input_fmap_154[7:0]) +
	( 15'sd 14224) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10835) * $signed(input_fmap_156[7:0]) +
	( 16'sd 32405) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8665) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3145) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_160[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4518) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28995) * $signed(input_fmap_163[7:0]) +
	( 14'sd 5534) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10943) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12840) * $signed(input_fmap_166[7:0]) +
	( 15'sd 11491) * $signed(input_fmap_167[7:0]) +
	( 15'sd 11403) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17677) * $signed(input_fmap_169[7:0]) +
	( 15'sd 10523) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24907) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4189) * $signed(input_fmap_172[7:0]) +
	( 15'sd 8746) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32553) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21050) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18986) * $signed(input_fmap_176[7:0]) +
	( 15'sd 9372) * $signed(input_fmap_177[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_178[7:0]) +
	( 16'sd 32081) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_180[7:0]) +
	( 15'sd 9079) * $signed(input_fmap_181[7:0]) +
	( 14'sd 7575) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29000) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22549) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11312) * $signed(input_fmap_185[7:0]) +
	( 16'sd 31009) * $signed(input_fmap_186[7:0]) +
	( 15'sd 8492) * $signed(input_fmap_187[7:0]) +
	( 16'sd 30066) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17905) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30857) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14928) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20108) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29820) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1823) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5972) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31807) * $signed(input_fmap_197[7:0]) +
	( 14'sd 8174) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10905) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29568) * $signed(input_fmap_200[7:0]) +
	( 14'sd 4229) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17460) * $signed(input_fmap_202[7:0]) +
	( 15'sd 11461) * $signed(input_fmap_203[7:0]) +
	( 15'sd 9546) * $signed(input_fmap_204[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_205[7:0]) +
	( 16'sd 17341) * $signed(input_fmap_206[7:0]) +
	( 15'sd 16217) * $signed(input_fmap_207[7:0]) +
	( 10'sd 392) * $signed(input_fmap_208[7:0]) +
	( 16'sd 25514) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3642) * $signed(input_fmap_210[7:0]) +
	( 15'sd 14525) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24114) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23458) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29897) * $signed(input_fmap_215[7:0]) +
	( 14'sd 7893) * $signed(input_fmap_216[7:0]) +
	( 16'sd 16994) * $signed(input_fmap_217[7:0]) +
	( 14'sd 4539) * $signed(input_fmap_218[7:0]) +
	( 15'sd 16265) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28930) * $signed(input_fmap_220[7:0]) +
	( 16'sd 21356) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5996) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22859) * $signed(input_fmap_223[7:0]) +
	( 13'sd 3479) * $signed(input_fmap_224[7:0]) +
	( 15'sd 8762) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32362) * $signed(input_fmap_226[7:0]) +
	( 16'sd 30288) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25666) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17191) * $signed(input_fmap_229[7:0]) +
	( 15'sd 8874) * $signed(input_fmap_230[7:0]) +
	( 14'sd 5073) * $signed(input_fmap_231[7:0]) +
	( 15'sd 16061) * $signed(input_fmap_232[7:0]) +
	( 16'sd 31548) * $signed(input_fmap_233[7:0]) +
	( 11'sd 855) * $signed(input_fmap_234[7:0]) +
	( 13'sd 4034) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10161) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27249) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19004) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23314) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5648) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17696) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31472) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24267) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17851) * $signed(input_fmap_247[7:0]) +
	( 16'sd 30031) * $signed(input_fmap_248[7:0]) +
	( 16'sd 26472) * $signed(input_fmap_249[7:0]) +
	( 16'sd 21098) * $signed(input_fmap_250[7:0]) +
	( 12'sd 1969) * $signed(input_fmap_251[7:0]) +
	( 16'sd 23742) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13810) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14914) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_100;
assign conv_mac_100 = 
	( 15'sd 10411) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21449) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31528) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20997) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7430) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4993) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17289) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4636) * $signed(input_fmap_9[7:0]) +
	( 11'sd 721) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26152) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1830) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15156) * $signed(input_fmap_13[7:0]) +
	( 16'sd 30208) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10510) * $signed(input_fmap_15[7:0]) +
	( 11'sd 659) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32582) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18934) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16624) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20587) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1324) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4773) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20095) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23801) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30894) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20070) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32518) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15069) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1897) * $signed(input_fmap_33[7:0]) +
	( 14'sd 8155) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20954) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7301) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18566) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26773) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22330) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32569) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16057) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27138) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29876) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16133) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28651) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22644) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28687) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14428) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18761) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1232) * $signed(input_fmap_52[7:0]) +
	( 9'sd 250) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22138) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11346) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20155) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15129) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9822) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21227) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19602) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12929) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5430) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6125) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11352) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11617) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22920) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11911) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29120) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21659) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2072) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21569) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8812) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13757) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2799) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17513) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2509) * $signed(input_fmap_79[7:0]) +
	( 10'sd 313) * $signed(input_fmap_80[7:0]) +
	( 15'sd 15496) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23320) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9375) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28658) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5116) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21044) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30209) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16444) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8943) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23824) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20473) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17275) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13935) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9841) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10654) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_101[7:0]) +
	( 11'sd 651) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22722) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13295) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31562) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2383) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27485) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6594) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17361) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16450) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7078) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21236) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29344) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3837) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1638) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24065) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24880) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_119[7:0]) +
	( 9'sd 229) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23360) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19936) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7701) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6986) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12864) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26425) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32212) * $signed(input_fmap_127[7:0]) +
	( 16'sd 28051) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1729) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27228) * $signed(input_fmap_130[7:0]) +
	( 16'sd 21194) * $signed(input_fmap_131[7:0]) +
	( 13'sd 3899) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11758) * $signed(input_fmap_133[7:0]) +
	( 14'sd 7072) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27559) * $signed(input_fmap_135[7:0]) +
	( 16'sd 24051) * $signed(input_fmap_136[7:0]) +
	( 16'sd 19666) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32190) * $signed(input_fmap_138[7:0]) +
	( 16'sd 30858) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26823) * $signed(input_fmap_140[7:0]) +
	( 13'sd 2548) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30601) * $signed(input_fmap_142[7:0]) +
	( 15'sd 9440) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2608) * $signed(input_fmap_144[7:0]) +
	( 16'sd 24007) * $signed(input_fmap_145[7:0]) +
	( 13'sd 2292) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27782) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20427) * $signed(input_fmap_148[7:0]) +
	( 16'sd 26592) * $signed(input_fmap_149[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_151[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_152[7:0]) +
	( 16'sd 18978) * $signed(input_fmap_153[7:0]) +
	( 16'sd 16913) * $signed(input_fmap_154[7:0]) +
	( 16'sd 16784) * $signed(input_fmap_155[7:0]) +
	( 15'sd 12832) * $signed(input_fmap_156[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_157[7:0]) +
	( 13'sd 3667) * $signed(input_fmap_158[7:0]) +
	( 16'sd 17588) * $signed(input_fmap_159[7:0]) +
	( 16'sd 19843) * $signed(input_fmap_160[7:0]) +
	( 10'sd 408) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24986) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24579) * $signed(input_fmap_164[7:0]) +
	( 16'sd 20972) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13847) * $signed(input_fmap_166[7:0]) +
	( 15'sd 10897) * $signed(input_fmap_167[7:0]) +
	( 16'sd 31632) * $signed(input_fmap_168[7:0]) +
	( 11'sd 967) * $signed(input_fmap_169[7:0]) +
	( 16'sd 16475) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18644) * $signed(input_fmap_171[7:0]) +
	( 16'sd 32445) * $signed(input_fmap_172[7:0]) +
	( 16'sd 17386) * $signed(input_fmap_173[7:0]) +
	( 15'sd 13598) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_175[7:0]) +
	( 16'sd 23967) * $signed(input_fmap_176[7:0]) +
	( 15'sd 14438) * $signed(input_fmap_177[7:0]) +
	( 15'sd 8702) * $signed(input_fmap_178[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29006) * $signed(input_fmap_180[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4741) * $signed(input_fmap_182[7:0]) +
	( 11'sd 617) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_184[7:0]) +
	( 16'sd 30398) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17856) * $signed(input_fmap_186[7:0]) +
	( 15'sd 10781) * $signed(input_fmap_187[7:0]) +
	( 16'sd 19111) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26236) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17263) * $signed(input_fmap_190[7:0]) +
	( 16'sd 28324) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24432) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5858) * $signed(input_fmap_193[7:0]) +
	( 15'sd 11097) * $signed(input_fmap_194[7:0]) +
	( 16'sd 31293) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17968) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1206) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19926) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14437) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16413) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11994) * $signed(input_fmap_202[7:0]) +
	( 16'sd 29435) * $signed(input_fmap_203[7:0]) +
	( 16'sd 25745) * $signed(input_fmap_204[7:0]) +
	( 16'sd 19956) * $signed(input_fmap_205[7:0]) +
	( 14'sd 8042) * $signed(input_fmap_206[7:0]) +
	( 16'sd 26618) * $signed(input_fmap_207[7:0]) +
	( 15'sd 9758) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3652) * $signed(input_fmap_209[7:0]) +
	( 14'sd 7670) * $signed(input_fmap_210[7:0]) +
	( 12'sd 1856) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1774) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11046) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18197) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2853) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20556) * $signed(input_fmap_216[7:0]) +
	( 15'sd 14055) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22651) * $signed(input_fmap_218[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21810) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12128) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25577) * $signed(input_fmap_222[7:0]) +
	( 16'sd 21613) * $signed(input_fmap_223[7:0]) +
	( 15'sd 10488) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20594) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_226[7:0]) +
	( 15'sd 11652) * $signed(input_fmap_227[7:0]) +
	( 13'sd 3068) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20234) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30081) * $signed(input_fmap_230[7:0]) +
	( 14'sd 4756) * $signed(input_fmap_231[7:0]) +
	( 16'sd 30635) * $signed(input_fmap_232[7:0]) +
	( 15'sd 8712) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23718) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11059) * $signed(input_fmap_235[7:0]) +
	( 16'sd 20644) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11654) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13851) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26288) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1490) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30091) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28109) * $signed(input_fmap_242[7:0]) +
	( 16'sd 29911) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19957) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2393) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20040) * $signed(input_fmap_246[7:0]) +
	( 16'sd 24158) * $signed(input_fmap_247[7:0]) +
	( 15'sd 15468) * $signed(input_fmap_248[7:0]) +
	( 16'sd 20742) * $signed(input_fmap_249[7:0]) +
	( 16'sd 23882) * $signed(input_fmap_250[7:0]) +
	( 16'sd 17027) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30651) * $signed(input_fmap_252[7:0]) +
	( 16'sd 19906) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19835) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20790) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_101;
assign conv_mac_101 = 
	( 12'sd 1434) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13476) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15492) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30570) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6508) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16472) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11366) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16932) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20951) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29152) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25866) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31669) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21369) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32759) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20353) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17917) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32388) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6026) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28799) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29713) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14712) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2567) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17902) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17893) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27680) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12884) * $signed(input_fmap_27[7:0]) +
	( 14'sd 5737) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27725) * $signed(input_fmap_29[7:0]) +
	( 11'sd 959) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12729) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30059) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19152) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3699) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29499) * $signed(input_fmap_35[7:0]) +
	( 15'sd 16098) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32037) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5602) * $signed(input_fmap_38[7:0]) +
	( 8'sd 112) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28281) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23452) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5737) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25688) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6628) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6916) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23472) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23249) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14273) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6570) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20448) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4848) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9249) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14327) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9326) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14595) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30575) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31606) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14813) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19972) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19342) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2106) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15193) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14320) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32105) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20377) * $signed(input_fmap_68[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29812) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3016) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10711) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7341) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18272) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3533) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8687) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29454) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11045) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8562) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24402) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26555) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1932) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13247) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11024) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31239) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13147) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9347) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14852) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28479) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4785) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27875) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15880) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22973) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13016) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18814) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8279) * $signed(input_fmap_98[7:0]) +
	( 11'sd 996) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31699) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25517) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26364) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10738) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15951) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31404) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28760) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21263) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8872) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23602) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20541) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3271) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13515) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15515) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22517) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8370) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32709) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5615) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21172) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17904) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21944) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28137) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7435) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17883) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23468) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5630) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30913) * $signed(input_fmap_130[7:0]) +
	( 14'sd 4410) * $signed(input_fmap_131[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_132[7:0]) +
	( 14'sd 7655) * $signed(input_fmap_133[7:0]) +
	( 14'sd 6910) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2840) * $signed(input_fmap_136[7:0]) +
	( 15'sd 10558) * $signed(input_fmap_137[7:0]) +
	( 12'sd 1421) * $signed(input_fmap_138[7:0]) +
	( 15'sd 13134) * $signed(input_fmap_139[7:0]) +
	( 15'sd 11181) * $signed(input_fmap_140[7:0]) +
	( 14'sd 4202) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26823) * $signed(input_fmap_143[7:0]) +
	( 16'sd 23485) * $signed(input_fmap_144[7:0]) +
	( 16'sd 32540) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7746) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14035) * $signed(input_fmap_147[7:0]) +
	( 14'sd 7077) * $signed(input_fmap_148[7:0]) +
	( 16'sd 16493) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27644) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18808) * $signed(input_fmap_151[7:0]) +
	( 13'sd 4057) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27656) * $signed(input_fmap_153[7:0]) +
	( 16'sd 17681) * $signed(input_fmap_154[7:0]) +
	( 16'sd 31191) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30898) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17225) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26012) * $signed(input_fmap_159[7:0]) +
	( 16'sd 28062) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1087) * $signed(input_fmap_161[7:0]) +
	( 15'sd 12841) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27973) * $signed(input_fmap_163[7:0]) +
	( 15'sd 14135) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14874) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_166[7:0]) +
	( 15'sd 14362) * $signed(input_fmap_167[7:0]) +
	( 15'sd 12557) * $signed(input_fmap_168[7:0]) +
	( 14'sd 5114) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20533) * $signed(input_fmap_170[7:0]) +
	( 16'sd 25766) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_172[7:0]) +
	( 14'sd 6915) * $signed(input_fmap_173[7:0]) +
	( 14'sd 5482) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15240) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7548) * $signed(input_fmap_177[7:0]) +
	( 15'sd 11099) * $signed(input_fmap_178[7:0]) +
	( 16'sd 32080) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27054) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28625) * $signed(input_fmap_181[7:0]) +
	( 16'sd 27670) * $signed(input_fmap_182[7:0]) +
	( 11'sd 540) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31528) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_185[7:0]) +
	( 16'sd 27662) * $signed(input_fmap_186[7:0]) +
	( 16'sd 20264) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1194) * $signed(input_fmap_188[7:0]) +
	( 15'sd 8799) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17276) * $signed(input_fmap_190[7:0]) +
	( 16'sd 28593) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20729) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22062) * $signed(input_fmap_193[7:0]) +
	( 16'sd 20089) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29728) * $signed(input_fmap_195[7:0]) +
	( 16'sd 29290) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14545) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2624) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_199[7:0]) +
	( 15'sd 12038) * $signed(input_fmap_200[7:0]) +
	( 16'sd 31754) * $signed(input_fmap_201[7:0]) +
	( 15'sd 9614) * $signed(input_fmap_202[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19378) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6121) * $signed(input_fmap_205[7:0]) +
	( 16'sd 22312) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21378) * $signed(input_fmap_207[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_208[7:0]) +
	( 14'sd 5626) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19149) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15322) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18691) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12075) * $signed(input_fmap_213[7:0]) +
	( 15'sd 16042) * $signed(input_fmap_214[7:0]) +
	( 16'sd 26095) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4425) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5522) * $signed(input_fmap_218[7:0]) +
	( 16'sd 25325) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19097) * $signed(input_fmap_221[7:0]) +
	( 15'sd 13674) * $signed(input_fmap_222[7:0]) +
	( 15'sd 10574) * $signed(input_fmap_223[7:0]) +
	( 16'sd 31651) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15441) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11996) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9928) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18635) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6404) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7972) * $signed(input_fmap_230[7:0]) +
	( 15'sd 11213) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15630) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24318) * $signed(input_fmap_233[7:0]) +
	( 15'sd 16357) * $signed(input_fmap_234[7:0]) +
	( 16'sd 30329) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12539) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6883) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13835) * $signed(input_fmap_238[7:0]) +
	( 16'sd 17275) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6748) * $signed(input_fmap_240[7:0]) +
	( 16'sd 16476) * $signed(input_fmap_241[7:0]) +
	( 16'sd 30082) * $signed(input_fmap_242[7:0]) +
	( 16'sd 21533) * $signed(input_fmap_243[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2788) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28856) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15170) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15467) * $signed(input_fmap_249[7:0]) +
	( 12'sd 1802) * $signed(input_fmap_250[7:0]) +
	( 13'sd 4073) * $signed(input_fmap_251[7:0]) +
	( 16'sd 32444) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28931) * $signed(input_fmap_253[7:0]) +
	( 15'sd 15527) * $signed(input_fmap_254[7:0]) +
	( 15'sd 15785) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_102;
assign conv_mac_102 = 
	( 16'sd 24030) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30787) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10058) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27714) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25991) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11461) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23404) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29526) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17088) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25851) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17283) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14673) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21129) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6006) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21087) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1911) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14964) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10833) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26292) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13834) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28804) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13019) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30293) * $signed(input_fmap_26[7:0]) +
	( 11'sd 561) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4756) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10990) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23194) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27685) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7363) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19501) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3943) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23113) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15288) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30542) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15080) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6794) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14695) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5838) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23562) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13586) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2205) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18342) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26682) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10039) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18887) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10219) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21873) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32112) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29157) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22440) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2072) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18538) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25282) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2327) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14206) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8593) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13331) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25203) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19554) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28555) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32557) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13174) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25098) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18281) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29324) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31269) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_74[7:0]) +
	( 10'sd 494) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18001) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21819) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19470) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17217) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2481) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11867) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22273) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5137) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14218) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10080) * $signed(input_fmap_88[7:0]) +
	( 13'sd 4054) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20559) * $signed(input_fmap_90[7:0]) +
	( 14'sd 8191) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30840) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1229) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14694) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28376) * $signed(input_fmap_95[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27063) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31453) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15123) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6465) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5089) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17476) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25582) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18936) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18989) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30680) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10045) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25552) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16463) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20485) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6212) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25280) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14776) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32238) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32559) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30241) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30784) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16620) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10685) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6078) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18460) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11947) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30324) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23173) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3449) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32489) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8245) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28646) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25933) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15656) * $signed(input_fmap_131[7:0]) +
	( 16'sd 19042) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22592) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4771) * $signed(input_fmap_134[7:0]) +
	( 16'sd 30199) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_136[7:0]) +
	( 16'sd 16686) * $signed(input_fmap_137[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_138[7:0]) +
	( 14'sd 7418) * $signed(input_fmap_139[7:0]) +
	( 16'sd 31417) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3739) * $signed(input_fmap_141[7:0]) +
	( 16'sd 32648) * $signed(input_fmap_142[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_143[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_144[7:0]) +
	( 15'sd 9035) * $signed(input_fmap_145[7:0]) +
	( 14'sd 4890) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3097) * $signed(input_fmap_148[7:0]) +
	( 16'sd 29921) * $signed(input_fmap_149[7:0]) +
	( 16'sd 20530) * $signed(input_fmap_150[7:0]) +
	( 15'sd 11193) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22929) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23615) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27085) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20579) * $signed(input_fmap_156[7:0]) +
	( 16'sd 16748) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12170) * $signed(input_fmap_159[7:0]) +
	( 13'sd 3871) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31770) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13388) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2398) * $signed(input_fmap_163[7:0]) +
	( 16'sd 27612) * $signed(input_fmap_164[7:0]) +
	( 16'sd 21136) * $signed(input_fmap_165[7:0]) +
	( 14'sd 5249) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24331) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4262) * $signed(input_fmap_168[7:0]) +
	( 15'sd 15711) * $signed(input_fmap_169[7:0]) +
	( 14'sd 4700) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15076) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15904) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1025) * $signed(input_fmap_173[7:0]) +
	( 16'sd 21374) * $signed(input_fmap_174[7:0]) +
	( 15'sd 9387) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21697) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27147) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32608) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15857) * $signed(input_fmap_179[7:0]) +
	( 15'sd 11650) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3476) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26189) * $signed(input_fmap_182[7:0]) +
	( 16'sd 28681) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24355) * $signed(input_fmap_184[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6745) * $signed(input_fmap_186[7:0]) +
	( 11'sd 872) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2853) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7574) * $signed(input_fmap_189[7:0]) +
	( 16'sd 18728) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3777) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20558) * $signed(input_fmap_192[7:0]) +
	( 14'sd 7620) * $signed(input_fmap_193[7:0]) +
	( 14'sd 4540) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29044) * $signed(input_fmap_195[7:0]) +
	( 15'sd 9480) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19761) * $signed(input_fmap_197[7:0]) +
	( 16'sd 16550) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16041) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18870) * $signed(input_fmap_200[7:0]) +
	( 14'sd 4476) * $signed(input_fmap_201[7:0]) +
	( 16'sd 28041) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21115) * $signed(input_fmap_203[7:0]) +
	( 16'sd 29849) * $signed(input_fmap_204[7:0]) +
	( 11'sd 713) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28581) * $signed(input_fmap_206[7:0]) +
	( 14'sd 4277) * $signed(input_fmap_207[7:0]) +
	( 16'sd 21021) * $signed(input_fmap_208[7:0]) +
	( 15'sd 16231) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11637) * $signed(input_fmap_210[7:0]) +
	( 16'sd 27111) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_213[7:0]) +
	( 15'sd 16139) * $signed(input_fmap_214[7:0]) +
	( 15'sd 12828) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_216[7:0]) +
	( 11'sd 714) * $signed(input_fmap_217[7:0]) +
	( 15'sd 11062) * $signed(input_fmap_218[7:0]) +
	( 16'sd 26359) * $signed(input_fmap_219[7:0]) +
	( 14'sd 7561) * $signed(input_fmap_220[7:0]) +
	( 16'sd 24757) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28825) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25066) * $signed(input_fmap_223[7:0]) +
	( 11'sd 770) * $signed(input_fmap_224[7:0]) +
	( 16'sd 29229) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10724) * $signed(input_fmap_226[7:0]) +
	( 16'sd 25250) * $signed(input_fmap_227[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17325) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28090) * $signed(input_fmap_230[7:0]) +
	( 16'sd 22694) * $signed(input_fmap_231[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_232[7:0]) +
	( 16'sd 29509) * $signed(input_fmap_233[7:0]) +
	( 16'sd 22209) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29296) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23632) * $signed(input_fmap_236[7:0]) +
	( 16'sd 16678) * $signed(input_fmap_237[7:0]) +
	( 16'sd 26619) * $signed(input_fmap_238[7:0]) +
	( 13'sd 3902) * $signed(input_fmap_239[7:0]) +
	( 15'sd 16227) * $signed(input_fmap_240[7:0]) +
	( 15'sd 8844) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28658) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13334) * $signed(input_fmap_244[7:0]) +
	( 16'sd 23014) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17321) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27444) * $signed(input_fmap_247[7:0]) +
	( 15'sd 8398) * $signed(input_fmap_248[7:0]) +
	( 14'sd 7303) * $signed(input_fmap_249[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7125) * $signed(input_fmap_251[7:0]) +
	( 16'sd 21963) * $signed(input_fmap_252[7:0]) +
	( 15'sd 9107) * $signed(input_fmap_253[7:0]) +
	( 16'sd 25472) * $signed(input_fmap_254[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_103;
assign conv_mac_103 = 
	( 16'sd 22920) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17838) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19561) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1531) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2218) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25554) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11490) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30714) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11027) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31584) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8845) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19952) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20003) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20902) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4585) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4261) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11348) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15742) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17804) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25410) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24010) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_21[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21913) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13203) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27001) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12116) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29175) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14864) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3272) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11606) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30417) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14580) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26317) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11883) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2547) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26944) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18278) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16789) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11928) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7048) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19508) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11000) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13215) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12555) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22106) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27473) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2875) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6690) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27804) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15974) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29572) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32733) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10354) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5335) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29223) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32622) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27442) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8333) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27691) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7283) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22903) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30183) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9245) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32686) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13619) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19930) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10491) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31525) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15950) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4603) * $signed(input_fmap_77[7:0]) +
	( 13'sd 4014) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5234) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11509) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12565) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28664) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4205) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16702) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6628) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26568) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8237) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7578) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3409) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11085) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5562) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2630) * $signed(input_fmap_94[7:0]) +
	( 11'sd 689) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10868) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26037) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20014) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19833) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3913) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22622) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11436) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30717) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3975) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4247) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27843) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4974) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31621) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15818) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14842) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12719) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2051) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11740) * $signed(input_fmap_114[7:0]) +
	( 10'sd 456) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28921) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24252) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11533) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3670) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12605) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22401) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11525) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12550) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24649) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8817) * $signed(input_fmap_128[7:0]) +
	( 11'sd 583) * $signed(input_fmap_129[7:0]) +
	( 15'sd 11598) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5912) * $signed(input_fmap_131[7:0]) +
	( 13'sd 3088) * $signed(input_fmap_132[7:0]) +
	( 16'sd 23848) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25220) * $signed(input_fmap_134[7:0]) +
	( 16'sd 25750) * $signed(input_fmap_135[7:0]) +
	( 16'sd 19564) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11434) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28737) * $signed(input_fmap_139[7:0]) +
	( 14'sd 5148) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19487) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21832) * $signed(input_fmap_142[7:0]) +
	( 13'sd 2881) * $signed(input_fmap_143[7:0]) +
	( 15'sd 12553) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28397) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19983) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_147[7:0]) +
	( 16'sd 30721) * $signed(input_fmap_148[7:0]) +
	( 11'sd 664) * $signed(input_fmap_149[7:0]) +
	( 16'sd 20472) * $signed(input_fmap_150[7:0]) +
	( 16'sd 31241) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23455) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12889) * $signed(input_fmap_153[7:0]) +
	( 10'sd 438) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20476) * $signed(input_fmap_155[7:0]) +
	( 16'sd 21509) * $signed(input_fmap_156[7:0]) +
	( 15'sd 9698) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8426) * $signed(input_fmap_158[7:0]) +
	( 16'sd 22302) * $signed(input_fmap_159[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28973) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_162[7:0]) +
	( 14'sd 6812) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9336) * $signed(input_fmap_164[7:0]) +
	( 16'sd 26649) * $signed(input_fmap_165[7:0]) +
	( 16'sd 17890) * $signed(input_fmap_166[7:0]) +
	( 16'sd 18681) * $signed(input_fmap_167[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_168[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_169[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30470) * $signed(input_fmap_171[7:0]) +
	( 15'sd 10850) * $signed(input_fmap_172[7:0]) +
	( 13'sd 2199) * $signed(input_fmap_173[7:0]) +
	( 16'sd 22655) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28653) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13252) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22345) * $signed(input_fmap_177[7:0]) +
	( 16'sd 21559) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25332) * $signed(input_fmap_179[7:0]) +
	( 16'sd 19982) * $signed(input_fmap_180[7:0]) +
	( 15'sd 16140) * $signed(input_fmap_181[7:0]) +
	( 15'sd 14745) * $signed(input_fmap_182[7:0]) +
	( 16'sd 20226) * $signed(input_fmap_183[7:0]) +
	( 11'sd 872) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12248) * $signed(input_fmap_186[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_187[7:0]) +
	( 16'sd 25140) * $signed(input_fmap_188[7:0]) +
	( 15'sd 8957) * $signed(input_fmap_189[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14348) * $signed(input_fmap_191[7:0]) +
	( 13'sd 3733) * $signed(input_fmap_192[7:0]) +
	( 16'sd 23869) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27809) * $signed(input_fmap_195[7:0]) +
	( 15'sd 9644) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15458) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10445) * $signed(input_fmap_198[7:0]) +
	( 9'sd 141) * $signed(input_fmap_199[7:0]) +
	( 16'sd 30034) * $signed(input_fmap_200[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6774) * $signed(input_fmap_203[7:0]) +
	( 16'sd 28859) * $signed(input_fmap_204[7:0]) +
	( 16'sd 16635) * $signed(input_fmap_205[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_207[7:0]) +
	( 12'sd 1938) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20545) * $signed(input_fmap_209[7:0]) +
	( 16'sd 20908) * $signed(input_fmap_210[7:0]) +
	( 16'sd 19437) * $signed(input_fmap_211[7:0]) +
	( 11'sd 581) * $signed(input_fmap_212[7:0]) +
	( 16'sd 19414) * $signed(input_fmap_213[7:0]) +
	( 10'sd 276) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7860) * $signed(input_fmap_215[7:0]) +
	( 16'sd 26675) * $signed(input_fmap_216[7:0]) +
	( 14'sd 5078) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31798) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14289) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4840) * $signed(input_fmap_220[7:0]) +
	( 15'sd 14601) * $signed(input_fmap_221[7:0]) +
	( 16'sd 26106) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24016) * $signed(input_fmap_223[7:0]) +
	( 16'sd 20389) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20633) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18584) * $signed(input_fmap_226[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8720) * $signed(input_fmap_228[7:0]) +
	( 16'sd 19646) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_230[7:0]) +
	( 15'sd 12945) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18995) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14395) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13879) * $signed(input_fmap_234[7:0]) +
	( 16'sd 27014) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27105) * $signed(input_fmap_236[7:0]) +
	( 12'sd 1448) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5999) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22309) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6734) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25904) * $signed(input_fmap_241[7:0]) +
	( 16'sd 25509) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10199) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_244[7:0]) +
	( 16'sd 18550) * $signed(input_fmap_245[7:0]) +
	( 13'sd 3484) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18306) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13248) * $signed(input_fmap_248[7:0]) +
	( 16'sd 27432) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25212) * $signed(input_fmap_250[7:0]) +
	( 16'sd 31459) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28832) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1064) * $signed(input_fmap_254[7:0]) +
	( 15'sd 13404) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_104;
assign conv_mac_104 = 
	( 15'sd 9056) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4927) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3696) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8284) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24975) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11383) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31131) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30919) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30309) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15331) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17347) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2971) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14350) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23591) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10478) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4218) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7938) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3569) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18241) * $signed(input_fmap_18[7:0]) +
	( 15'sd 12387) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25137) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7744) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1300) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24944) * $signed(input_fmap_23[7:0]) +
	( 16'sd 23333) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8085) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11460) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14398) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30828) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13695) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28473) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12994) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32419) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3545) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24718) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10893) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26449) * $signed(input_fmap_37[7:0]) +
	( 15'sd 16075) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26087) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10304) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4461) * $signed(input_fmap_41[7:0]) +
	( 11'sd 549) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18448) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19807) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16806) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26180) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7767) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21401) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32300) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28909) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10675) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27780) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17318) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29596) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12021) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29730) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20226) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22678) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29104) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26026) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29321) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17689) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18319) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14270) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5950) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4128) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6388) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19125) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22403) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1320) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31081) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25914) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31985) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11075) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10788) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11474) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7867) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19344) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21898) * $signed(input_fmap_83[7:0]) +
	( 10'sd 465) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26658) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28923) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25943) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24016) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27877) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3725) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15774) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12283) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26850) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4983) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2653) * $signed(input_fmap_96[7:0]) +
	( 12'sd 2044) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23845) * $signed(input_fmap_98[7:0]) +
	( 11'sd 553) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25011) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6533) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5802) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10403) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13434) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8243) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30913) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26883) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9158) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11510) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24196) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2889) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19107) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29102) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1852) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10109) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26817) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13383) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5817) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21000) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26604) * $signed(input_fmap_122[7:0]) +
	( 13'sd 4004) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18712) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31169) * $signed(input_fmap_125[7:0]) +
	( 10'sd 329) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_127[7:0]) +
	( 16'sd 20326) * $signed(input_fmap_128[7:0]) +
	( 16'sd 20598) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1862) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14618) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10180) * $signed(input_fmap_132[7:0]) +
	( 16'sd 18471) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5141) * $signed(input_fmap_134[7:0]) +
	( 15'sd 8667) * $signed(input_fmap_135[7:0]) +
	( 16'sd 29441) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12796) * $signed(input_fmap_137[7:0]) +
	( 14'sd 4565) * $signed(input_fmap_138[7:0]) +
	( 16'sd 29085) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30435) * $signed(input_fmap_140[7:0]) +
	( 14'sd 4941) * $signed(input_fmap_141[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_142[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31808) * $signed(input_fmap_144[7:0]) +
	( 16'sd 18864) * $signed(input_fmap_145[7:0]) +
	( 16'sd 22227) * $signed(input_fmap_146[7:0]) +
	( 16'sd 31540) * $signed(input_fmap_147[7:0]) +
	( 16'sd 30370) * $signed(input_fmap_148[7:0]) +
	( 16'sd 32413) * $signed(input_fmap_149[7:0]) +
	( 15'sd 10952) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4298) * $signed(input_fmap_151[7:0]) +
	( 15'sd 9034) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17593) * $signed(input_fmap_153[7:0]) +
	( 16'sd 29745) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12619) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13055) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_157[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4775) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6396) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_161[7:0]) +
	( 16'sd 28486) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2336) * $signed(input_fmap_163[7:0]) +
	( 16'sd 29531) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23909) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12445) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20729) * $signed(input_fmap_167[7:0]) +
	( 11'sd 655) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25065) * $signed(input_fmap_169[7:0]) +
	( 16'sd 16846) * $signed(input_fmap_170[7:0]) +
	( 15'sd 8690) * $signed(input_fmap_171[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_172[7:0]) +
	( 11'sd 1005) * $signed(input_fmap_173[7:0]) +
	( 16'sd 23501) * $signed(input_fmap_174[7:0]) +
	( 16'sd 30776) * $signed(input_fmap_175[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_176[7:0]) +
	( 14'sd 4927) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10874) * $signed(input_fmap_178[7:0]) +
	( 13'sd 4035) * $signed(input_fmap_179[7:0]) +
	( 15'sd 9421) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18060) * $signed(input_fmap_181[7:0]) +
	( 15'sd 11763) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27230) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30991) * $signed(input_fmap_184[7:0]) +
	( 16'sd 20477) * $signed(input_fmap_185[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1709) * $signed(input_fmap_187[7:0]) +
	( 16'sd 20194) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7062) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17792) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31118) * $signed(input_fmap_191[7:0]) +
	( 14'sd 7653) * $signed(input_fmap_192[7:0]) +
	( 16'sd 25160) * $signed(input_fmap_193[7:0]) +
	( 13'sd 2176) * $signed(input_fmap_194[7:0]) +
	( 14'sd 6953) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15830) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26929) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27715) * $signed(input_fmap_198[7:0]) +
	( 11'sd 656) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29811) * $signed(input_fmap_200[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_201[7:0]) +
	( 15'sd 13753) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12581) * $signed(input_fmap_203[7:0]) +
	( 16'sd 21851) * $signed(input_fmap_204[7:0]) +
	( 15'sd 13785) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31363) * $signed(input_fmap_206[7:0]) +
	( 15'sd 14681) * $signed(input_fmap_207[7:0]) +
	( 15'sd 10738) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19795) * $signed(input_fmap_209[7:0]) +
	( 15'sd 13912) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23977) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19712) * $signed(input_fmap_212[7:0]) +
	( 16'sd 26849) * $signed(input_fmap_213[7:0]) +
	( 14'sd 4720) * $signed(input_fmap_214[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_215[7:0]) +
	( 11'sd 598) * $signed(input_fmap_216[7:0]) +
	( 15'sd 12206) * $signed(input_fmap_217[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10548) * $signed(input_fmap_219[7:0]) +
	( 15'sd 12137) * $signed(input_fmap_220[7:0]) +
	( 16'sd 24774) * $signed(input_fmap_221[7:0]) +
	( 16'sd 23466) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19750) * $signed(input_fmap_223[7:0]) +
	( 15'sd 9605) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5709) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24318) * $signed(input_fmap_227[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3248) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30186) * $signed(input_fmap_230[7:0]) +
	( 14'sd 4793) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9969) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18313) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19440) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5172) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30092) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_237[7:0]) +
	( 16'sd 29564) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31853) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22836) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29914) * $signed(input_fmap_241[7:0]) +
	( 15'sd 8443) * $signed(input_fmap_242[7:0]) +
	( 16'sd 29721) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6474) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5748) * $signed(input_fmap_245[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_246[7:0]) +
	( 16'sd 32753) * $signed(input_fmap_247[7:0]) +
	( 15'sd 12802) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14831) * $signed(input_fmap_249[7:0]) +
	( 16'sd 28275) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26003) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6595) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5832) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1755) * $signed(input_fmap_254[7:0]) +
	( 14'sd 6889) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_105;
assign conv_mac_105 = 
	( 15'sd 16163) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25507) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19677) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5391) * $signed(input_fmap_3[7:0]) +
	( 13'sd 4040) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17479) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11772) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5333) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5661) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6946) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32075) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30233) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18682) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23535) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30444) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31580) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18686) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18393) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19793) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31053) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1135) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29909) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32186) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8310) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30291) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29199) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22180) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2105) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24018) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30978) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12802) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23593) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9223) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8840) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23909) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28795) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10382) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18926) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10752) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7164) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1032) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2623) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4654) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16898) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8333) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15884) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32609) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21846) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31624) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29475) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2197) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24141) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22434) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9617) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13766) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26753) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5856) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17689) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18462) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25688) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20078) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27261) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5424) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27436) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19679) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15507) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29181) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17745) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29081) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25880) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8561) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16646) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5971) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13499) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21010) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24038) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25113) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9420) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1303) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22288) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11621) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15389) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10119) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26596) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30620) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14976) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22383) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4489) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16019) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32350) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20776) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21294) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10003) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18188) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7454) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15149) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13048) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24489) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26139) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31614) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28626) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24087) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6767) * $signed(input_fmap_116[7:0]) +
	( 14'sd 8074) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28454) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14626) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8353) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8965) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27560) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32191) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27042) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3596) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23683) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29325) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2576) * $signed(input_fmap_128[7:0]) +
	( 16'sd 32432) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10524) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5083) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14226) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12803) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32604) * $signed(input_fmap_134[7:0]) +
	( 13'sd 3539) * $signed(input_fmap_135[7:0]) +
	( 15'sd 14974) * $signed(input_fmap_136[7:0]) +
	( 13'sd 2180) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32414) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14499) * $signed(input_fmap_139[7:0]) +
	( 11'sd 572) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13860) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28996) * $signed(input_fmap_142[7:0]) +
	( 16'sd 24416) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2515) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29163) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21086) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23422) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12335) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21772) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23694) * $signed(input_fmap_151[7:0]) +
	( 12'sd 1502) * $signed(input_fmap_152[7:0]) +
	( 15'sd 13079) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23453) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20511) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25427) * $signed(input_fmap_157[7:0]) +
	( 16'sd 29472) * $signed(input_fmap_158[7:0]) +
	( 15'sd 15991) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17855) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1108) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21230) * $signed(input_fmap_162[7:0]) +
	( 15'sd 12937) * $signed(input_fmap_163[7:0]) +
	( 15'sd 12677) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11771) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13175) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17419) * $signed(input_fmap_168[7:0]) +
	( 16'sd 22344) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11545) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19145) * $signed(input_fmap_171[7:0]) +
	( 16'sd 28569) * $signed(input_fmap_172[7:0]) +
	( 16'sd 28165) * $signed(input_fmap_173[7:0]) +
	( 16'sd 24578) * $signed(input_fmap_174[7:0]) +
	( 15'sd 13804) * $signed(input_fmap_175[7:0]) +
	( 16'sd 23683) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2992) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31912) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22661) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6205) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_181[7:0]) +
	( 16'sd 32143) * $signed(input_fmap_182[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_184[7:0]) +
	( 15'sd 16021) * $signed(input_fmap_185[7:0]) +
	( 16'sd 31514) * $signed(input_fmap_186[7:0]) +
	( 16'sd 23349) * $signed(input_fmap_187[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_188[7:0]) +
	( 16'sd 32021) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27697) * $signed(input_fmap_190[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_192[7:0]) +
	( 16'sd 23617) * $signed(input_fmap_193[7:0]) +
	( 12'sd 1060) * $signed(input_fmap_194[7:0]) +
	( 15'sd 15708) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12561) * $signed(input_fmap_196[7:0]) +
	( 14'sd 7754) * $signed(input_fmap_197[7:0]) +
	( 16'sd 16824) * $signed(input_fmap_198[7:0]) +
	( 16'sd 32394) * $signed(input_fmap_199[7:0]) +
	( 16'sd 28916) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_201[7:0]) +
	( 16'sd 20853) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14490) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31768) * $signed(input_fmap_205[7:0]) +
	( 16'sd 22191) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17144) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15270) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22053) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30492) * $signed(input_fmap_210[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12970) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1403) * $signed(input_fmap_213[7:0]) +
	( 10'sd 494) * $signed(input_fmap_214[7:0]) +
	( 16'sd 32495) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19016) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25278) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13213) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_219[7:0]) +
	( 14'sd 5210) * $signed(input_fmap_220[7:0]) +
	( 14'sd 4453) * $signed(input_fmap_221[7:0]) +
	( 14'sd 7581) * $signed(input_fmap_222[7:0]) +
	( 14'sd 5915) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25532) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15386) * $signed(input_fmap_225[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_226[7:0]) +
	( 14'sd 8053) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25526) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8672) * $signed(input_fmap_229[7:0]) +
	( 15'sd 13342) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20467) * $signed(input_fmap_231[7:0]) +
	( 14'sd 5723) * $signed(input_fmap_232[7:0]) +
	( 14'sd 6943) * $signed(input_fmap_233[7:0]) +
	( 16'sd 31747) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11905) * $signed(input_fmap_235[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_236[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_237[7:0]) +
	( 15'sd 8311) * $signed(input_fmap_238[7:0]) +
	( 14'sd 4699) * $signed(input_fmap_239[7:0]) +
	( 16'sd 20464) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3588) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17933) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22180) * $signed(input_fmap_243[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_244[7:0]) +
	( 16'sd 18144) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31380) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11298) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26126) * $signed(input_fmap_248[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17514) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22220) * $signed(input_fmap_251[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28398) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20316) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26349) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_106;
assign conv_mac_106 = 
	( 16'sd 22635) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13548) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2871) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31641) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32746) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18181) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13905) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8643) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9302) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21097) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32490) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20663) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4358) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28581) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31315) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26742) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_16[7:0]) +
	( 14'sd 8001) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5971) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9120) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20429) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22716) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20912) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13153) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18672) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30393) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30587) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27653) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5416) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20167) * $signed(input_fmap_31[7:0]) +
	( 9'sd 199) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21865) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13638) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16361) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23926) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19583) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15876) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23002) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4789) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20088) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5678) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23031) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5381) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26795) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17497) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24911) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26387) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12690) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21536) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17526) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5154) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22519) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4362) * $signed(input_fmap_56[7:0]) +
	( 7'sd 40) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19266) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26988) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14601) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24483) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28062) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28696) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19073) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9254) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20683) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24933) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23779) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10811) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7314) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3264) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21971) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22018) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7399) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11519) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23512) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26824) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21516) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22476) * $signed(input_fmap_82[7:0]) +
	( 11'sd 791) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6021) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19634) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27433) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25556) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23383) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21943) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6907) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27395) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14844) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17568) * $signed(input_fmap_96[7:0]) +
	( 8'sd 83) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21465) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2872) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1117) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14987) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2375) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22869) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24454) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7308) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2112) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28970) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6760) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10242) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25428) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4837) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30932) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26138) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18176) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15279) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32091) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13112) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13559) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1996) * $signed(input_fmap_123[7:0]) +
	( 16'sd 19465) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26742) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20137) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1089) * $signed(input_fmap_127[7:0]) +
	( 14'sd 5019) * $signed(input_fmap_128[7:0]) +
	( 16'sd 25232) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30530) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24803) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1218) * $signed(input_fmap_132[7:0]) +
	( 15'sd 13835) * $signed(input_fmap_133[7:0]) +
	( 14'sd 6286) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23222) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21304) * $signed(input_fmap_136[7:0]) +
	( 16'sd 16903) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29440) * $signed(input_fmap_138[7:0]) +
	( 14'sd 5745) * $signed(input_fmap_139[7:0]) +
	( 15'sd 14921) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24507) * $signed(input_fmap_141[7:0]) +
	( 16'sd 23328) * $signed(input_fmap_142[7:0]) +
	( 16'sd 21865) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19437) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22147) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13983) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_148[7:0]) +
	( 16'sd 16818) * $signed(input_fmap_149[7:0]) +
	( 15'sd 10467) * $signed(input_fmap_150[7:0]) +
	( 15'sd 13023) * $signed(input_fmap_151[7:0]) +
	( 16'sd 27097) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25554) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31386) * $signed(input_fmap_154[7:0]) +
	( 16'sd 32477) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29915) * $signed(input_fmap_156[7:0]) +
	( 12'sd 1791) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18012) * $signed(input_fmap_158[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_159[7:0]) +
	( 12'sd 1275) * $signed(input_fmap_160[7:0]) +
	( 15'sd 11848) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_162[7:0]) +
	( 16'sd 19905) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9621) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_165[7:0]) +
	( 16'sd 29881) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9993) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9226) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12778) * $signed(input_fmap_169[7:0]) +
	( 15'sd 15121) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12279) * $signed(input_fmap_171[7:0]) +
	( 16'sd 32093) * $signed(input_fmap_172[7:0]) +
	( 11'sd 691) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27031) * $signed(input_fmap_174[7:0]) +
	( 15'sd 9463) * $signed(input_fmap_175[7:0]) +
	( 16'sd 25867) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19952) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17376) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6713) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15659) * $signed(input_fmap_180[7:0]) +
	( 15'sd 14884) * $signed(input_fmap_181[7:0]) +
	( 15'sd 9624) * $signed(input_fmap_182[7:0]) +
	( 13'sd 3131) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11535) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_185[7:0]) +
	( 16'sd 21605) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18201) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23124) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17011) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30863) * $signed(input_fmap_190[7:0]) +
	( 14'sd 6485) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_192[7:0]) +
	( 15'sd 16019) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14869) * $signed(input_fmap_194[7:0]) +
	( 16'sd 23028) * $signed(input_fmap_195[7:0]) +
	( 16'sd 27007) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5042) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5520) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29435) * $signed(input_fmap_199[7:0]) +
	( 15'sd 12266) * $signed(input_fmap_200[7:0]) +
	( 16'sd 20286) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14558) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12490) * $signed(input_fmap_203[7:0]) +
	( 16'sd 21889) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2955) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_206[7:0]) +
	( 15'sd 14526) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_208[7:0]) +
	( 14'sd 5794) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15529) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12738) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14992) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12874) * $signed(input_fmap_213[7:0]) +
	( 13'sd 4070) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17643) * $signed(input_fmap_215[7:0]) +
	( 15'sd 16157) * $signed(input_fmap_216[7:0]) +
	( 16'sd 20947) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21131) * $signed(input_fmap_218[7:0]) +
	( 15'sd 8363) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31883) * $signed(input_fmap_220[7:0]) +
	( 16'sd 26617) * $signed(input_fmap_221[7:0]) +
	( 14'sd 7879) * $signed(input_fmap_222[7:0]) +
	( 14'sd 6193) * $signed(input_fmap_223[7:0]) +
	( 11'sd 653) * $signed(input_fmap_224[7:0]) +
	( 16'sd 22064) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22386) * $signed(input_fmap_226[7:0]) +
	( 15'sd 16203) * $signed(input_fmap_227[7:0]) +
	( 15'sd 9079) * $signed(input_fmap_228[7:0]) +
	( 7'sd 36) * $signed(input_fmap_229[7:0]) +
	( 15'sd 8692) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_231[7:0]) +
	( 10'sd 457) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23168) * $signed(input_fmap_233[7:0]) +
	( 16'sd 25483) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14322) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28631) * $signed(input_fmap_236[7:0]) +
	( 16'sd 32252) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5391) * $signed(input_fmap_238[7:0]) +
	( 11'sd 999) * $signed(input_fmap_239[7:0]) +
	( 15'sd 11082) * $signed(input_fmap_240[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1809) * $signed(input_fmap_242[7:0]) +
	( 14'sd 4973) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18728) * $signed(input_fmap_244[7:0]) +
	( 12'sd 2045) * $signed(input_fmap_245[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_246[7:0]) +
	( 14'sd 4163) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1502) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4574) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7850) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_251[7:0]) +
	( 16'sd 25198) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29055) * $signed(input_fmap_253[7:0]) +
	( 10'sd 396) * $signed(input_fmap_254[7:0]) +
	( 15'sd 15347) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_107;
assign conv_mac_107 = 
	( 15'sd 10758) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8836) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18240) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7860) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30246) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19169) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4968) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29936) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7822) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22752) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1850) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24748) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12426) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19755) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15039) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22811) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7407) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30046) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11533) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2288) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2075) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32468) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28394) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22479) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22357) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20197) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1420) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11665) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6499) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23461) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25560) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27130) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25174) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4829) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4690) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21851) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18362) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24610) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30537) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19662) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25066) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14621) * $signed(input_fmap_45[7:0]) +
	( 13'sd 4041) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22691) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20615) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25653) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1916) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14425) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21197) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14406) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17532) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13874) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17955) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13707) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31361) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9658) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6118) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5057) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11405) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18715) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22986) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25726) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22823) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12671) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1572) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27443) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12001) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21550) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27903) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15005) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27557) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27857) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17474) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11326) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20465) * $signed(input_fmap_82[7:0]) +
	( 15'sd 13130) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30083) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5818) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18118) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4618) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20128) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17481) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18112) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12069) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23593) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24159) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26761) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29591) * $signed(input_fmap_96[7:0]) +
	( 11'sd 696) * $signed(input_fmap_97[7:0]) +
	( 12'sd 2028) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28428) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16682) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26704) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5518) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17965) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12491) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18785) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19844) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8497) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27884) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29530) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12861) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23376) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28028) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28081) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3335) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7418) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31752) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21481) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25981) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15643) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30471) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14170) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31612) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3136) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19341) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27237) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15914) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31412) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_129[7:0]) +
	( 14'sd 4644) * $signed(input_fmap_130[7:0]) +
	( 14'sd 4890) * $signed(input_fmap_131[7:0]) +
	( 14'sd 4585) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11154) * $signed(input_fmap_133[7:0]) +
	( 14'sd 7999) * $signed(input_fmap_134[7:0]) +
	( 16'sd 17052) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9330) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_138[7:0]) +
	( 14'sd 5487) * $signed(input_fmap_139[7:0]) +
	( 15'sd 13179) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19234) * $signed(input_fmap_141[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_142[7:0]) +
	( 16'sd 30924) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28518) * $signed(input_fmap_144[7:0]) +
	( 16'sd 16605) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27980) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13830) * $signed(input_fmap_147[7:0]) +
	( 15'sd 8689) * $signed(input_fmap_148[7:0]) +
	( 16'sd 24352) * $signed(input_fmap_149[7:0]) +
	( 16'sd 28577) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20463) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11633) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7264) * $signed(input_fmap_154[7:0]) +
	( 12'sd 1690) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29025) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9729) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5835) * $signed(input_fmap_159[7:0]) +
	( 10'sd 349) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20070) * $signed(input_fmap_161[7:0]) +
	( 14'sd 6146) * $signed(input_fmap_162[7:0]) +
	( 15'sd 12143) * $signed(input_fmap_163[7:0]) +
	( 15'sd 16358) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14761) * $signed(input_fmap_165[7:0]) +
	( 16'sd 26473) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17752) * $signed(input_fmap_167[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_168[7:0]) +
	( 16'sd 24000) * $signed(input_fmap_169[7:0]) +
	( 13'sd 3113) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19453) * $signed(input_fmap_171[7:0]) +
	( 10'sd 264) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12533) * $signed(input_fmap_173[7:0]) +
	( 15'sd 16232) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7835) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9857) * $signed(input_fmap_178[7:0]) +
	( 15'sd 13897) * $signed(input_fmap_179[7:0]) +
	( 14'sd 8044) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10417) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30989) * $signed(input_fmap_183[7:0]) +
	( 10'sd 455) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11272) * $signed(input_fmap_185[7:0]) +
	( 16'sd 22232) * $signed(input_fmap_186[7:0]) +
	( 15'sd 16381) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17611) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_189[7:0]) +
	( 15'sd 8380) * $signed(input_fmap_190[7:0]) +
	( 16'sd 30696) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28414) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12830) * $signed(input_fmap_193[7:0]) +
	( 16'sd 16446) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10391) * $signed(input_fmap_197[7:0]) +
	( 10'sd 386) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29356) * $signed(input_fmap_199[7:0]) +
	( 16'sd 22411) * $signed(input_fmap_200[7:0]) +
	( 16'sd 25171) * $signed(input_fmap_201[7:0]) +
	( 16'sd 27192) * $signed(input_fmap_202[7:0]) +
	( 15'sd 14443) * $signed(input_fmap_203[7:0]) +
	( 16'sd 23070) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28240) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27030) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11900) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7407) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9288) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17219) * $signed(input_fmap_211[7:0]) +
	( 16'sd 25700) * $signed(input_fmap_212[7:0]) +
	( 14'sd 4811) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23996) * $signed(input_fmap_214[7:0]) +
	( 11'sd 840) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11714) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_218[7:0]) +
	( 16'sd 24267) * $signed(input_fmap_219[7:0]) +
	( 16'sd 16564) * $signed(input_fmap_220[7:0]) +
	( 14'sd 4710) * $signed(input_fmap_221[7:0]) +
	( 10'sd 325) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15248) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19061) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15278) * $signed(input_fmap_225[7:0]) +
	( 16'sd 16716) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14477) * $signed(input_fmap_227[7:0]) +
	( 10'sd 334) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29808) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14382) * $signed(input_fmap_230[7:0]) +
	( 13'sd 2461) * $signed(input_fmap_231[7:0]) +
	( 15'sd 13935) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28823) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5292) * $signed(input_fmap_234[7:0]) +
	( 14'sd 4282) * $signed(input_fmap_235[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14272) * $signed(input_fmap_238[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9312) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20554) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5953) * $signed(input_fmap_242[7:0]) +
	( 16'sd 27899) * $signed(input_fmap_243[7:0]) +
	( 16'sd 21002) * $signed(input_fmap_244[7:0]) +
	( 14'sd 4362) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10094) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12222) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9907) * $signed(input_fmap_249[7:0]) +
	( 15'sd 10919) * $signed(input_fmap_250[7:0]) +
	( 13'sd 3940) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12041) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2679) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5442) * $signed(input_fmap_254[7:0]) +
	( 15'sd 8888) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_108;
assign conv_mac_108 = 
	( 14'sd 7311) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13800) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12813) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25446) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2915) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14997) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17181) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14107) * $signed(input_fmap_8[7:0]) +
	( 11'sd 1011) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15090) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16011) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14491) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6757) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27542) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2487) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1645) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28500) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21471) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27976) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15591) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1048) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7267) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28653) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1288) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13846) * $signed(input_fmap_27[7:0]) +
	( 11'sd 534) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9656) * $signed(input_fmap_29[7:0]) +
	( 14'sd 8122) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24694) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20841) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27599) * $signed(input_fmap_34[7:0]) +
	( 14'sd 8137) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1812) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17871) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24053) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3577) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15218) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1631) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3215) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3628) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31401) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9172) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13985) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18805) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11829) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28581) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18624) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16453) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23026) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11339) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29084) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24236) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27419) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14293) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31407) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4633) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18259) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20021) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12602) * $signed(input_fmap_63[7:0]) +
	( 9'sd 250) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12551) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12916) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18291) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17686) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29102) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6734) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23575) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4356) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6381) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10628) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4350) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22626) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18309) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31583) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19316) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13661) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27723) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22879) * $signed(input_fmap_83[7:0]) +
	( 14'sd 7154) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27032) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15653) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8821) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24703) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9111) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15640) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29104) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18013) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11589) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3254) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31605) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20477) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2170) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31741) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17980) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13978) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25402) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24145) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8364) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30728) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4960) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24202) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8366) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2523) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6795) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2928) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19280) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32442) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23040) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27475) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16474) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29150) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28796) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9485) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8870) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29512) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13209) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12447) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3982) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24632) * $signed(input_fmap_127[7:0]) +
	( 11'sd 529) * $signed(input_fmap_128[7:0]) +
	( 16'sd 30470) * $signed(input_fmap_129[7:0]) +
	( 11'sd 682) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13904) * $signed(input_fmap_131[7:0]) +
	( 15'sd 12464) * $signed(input_fmap_132[7:0]) +
	( 16'sd 25074) * $signed(input_fmap_133[7:0]) +
	( 10'sd 476) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23656) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25168) * $signed(input_fmap_136[7:0]) +
	( 11'sd 599) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32190) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11270) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_140[7:0]) +
	( 15'sd 16342) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27030) * $signed(input_fmap_142[7:0]) +
	( 16'sd 30320) * $signed(input_fmap_143[7:0]) +
	( 16'sd 17786) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27484) * $signed(input_fmap_145[7:0]) +
	( 16'sd 20064) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27638) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22739) * $signed(input_fmap_148[7:0]) +
	( 15'sd 9541) * $signed(input_fmap_149[7:0]) +
	( 14'sd 6142) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12610) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6040) * $signed(input_fmap_152[7:0]) +
	( 14'sd 7733) * $signed(input_fmap_153[7:0]) +
	( 15'sd 14821) * $signed(input_fmap_154[7:0]) +
	( 15'sd 9860) * $signed(input_fmap_155[7:0]) +
	( 16'sd 19976) * $signed(input_fmap_156[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4139) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2355) * $signed(input_fmap_159[7:0]) +
	( 16'sd 32708) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20107) * $signed(input_fmap_161[7:0]) +
	( 16'sd 19242) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10068) * $signed(input_fmap_164[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13033) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30504) * $signed(input_fmap_167[7:0]) +
	( 16'sd 18058) * $signed(input_fmap_168[7:0]) +
	( 13'sd 2620) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9619) * $signed(input_fmap_170[7:0]) +
	( 15'sd 8963) * $signed(input_fmap_171[7:0]) +
	( 16'sd 21187) * $signed(input_fmap_172[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_173[7:0]) +
	( 16'sd 31737) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28429) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10627) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24994) * $signed(input_fmap_177[7:0]) +
	( 14'sd 8173) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_179[7:0]) +
	( 16'sd 16713) * $signed(input_fmap_180[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_181[7:0]) +
	( 15'sd 13958) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30382) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14861) * $signed(input_fmap_184[7:0]) +
	( 16'sd 23635) * $signed(input_fmap_185[7:0]) +
	( 12'sd 1862) * $signed(input_fmap_186[7:0]) +
	( 16'sd 19858) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32361) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7538) * $signed(input_fmap_189[7:0]) +
	( 15'sd 8893) * $signed(input_fmap_190[7:0]) +
	( 15'sd 10104) * $signed(input_fmap_191[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9224) * $signed(input_fmap_193[7:0]) +
	( 12'sd 1404) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17391) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7769) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32485) * $signed(input_fmap_197[7:0]) +
	( 16'sd 16831) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6534) * $signed(input_fmap_199[7:0]) +
	( 16'sd 32333) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3461) * $signed(input_fmap_201[7:0]) +
	( 16'sd 30889) * $signed(input_fmap_202[7:0]) +
	( 16'sd 22252) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11777) * $signed(input_fmap_204[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12981) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28913) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28542) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20477) * $signed(input_fmap_209[7:0]) +
	( 16'sd 28411) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6726) * $signed(input_fmap_211[7:0]) +
	( 16'sd 25513) * $signed(input_fmap_212[7:0]) +
	( 16'sd 21218) * $signed(input_fmap_213[7:0]) +
	( 10'sd 486) * $signed(input_fmap_214[7:0]) +
	( 15'sd 13440) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23268) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17073) * $signed(input_fmap_217[7:0]) +
	( 15'sd 9485) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14137) * $signed(input_fmap_219[7:0]) +
	( 16'sd 20661) * $signed(input_fmap_220[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3675) * $signed(input_fmap_222[7:0]) +
	( 14'sd 5393) * $signed(input_fmap_223[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_224[7:0]) +
	( 16'sd 32406) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13513) * $signed(input_fmap_227[7:0]) +
	( 15'sd 13332) * $signed(input_fmap_228[7:0]) +
	( 15'sd 13156) * $signed(input_fmap_229[7:0]) +
	( 14'sd 4996) * $signed(input_fmap_230[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_231[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_232[7:0]) +
	( 16'sd 29848) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18087) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12322) * $signed(input_fmap_235[7:0]) +
	( 16'sd 17661) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20513) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_239[7:0]) +
	( 15'sd 12771) * $signed(input_fmap_240[7:0]) +
	( 15'sd 14111) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17259) * $signed(input_fmap_242[7:0]) +
	( 16'sd 24915) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1380) * $signed(input_fmap_244[7:0]) +
	( 15'sd 8702) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9116) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30464) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17977) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32445) * $signed(input_fmap_250[7:0]) +
	( 15'sd 10344) * $signed(input_fmap_251[7:0]) +
	( 16'sd 21671) * $signed(input_fmap_252[7:0]) +
	( 15'sd 9551) * $signed(input_fmap_253[7:0]) +
	( 11'sd 1005) * $signed(input_fmap_254[7:0]) +
	( 15'sd 16337) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_109;
assign conv_mac_109 = 
	( 16'sd 17698) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28506) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3425) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12021) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6301) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17131) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24135) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21213) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24055) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7772) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11955) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10384) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22222) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29406) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32741) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16462) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17662) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2651) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9255) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29372) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1706) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5369) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31059) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28069) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29900) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22349) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30828) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7625) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7782) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16473) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12821) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4288) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5279) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19444) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17617) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2378) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28927) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25732) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3046) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27441) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9501) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20526) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18995) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19037) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3039) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14795) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29533) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4922) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29564) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21552) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10822) * $signed(input_fmap_55[7:0]) +
	( 16'sd 24975) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4724) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5662) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18735) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3898) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11634) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27237) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15399) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14961) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6541) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4268) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32652) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21392) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30277) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16047) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30439) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25802) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11423) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31848) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26965) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23668) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26633) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4448) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22479) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24215) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17131) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19372) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21987) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30464) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3743) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25763) * $signed(input_fmap_89[7:0]) +
	( 14'sd 8054) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25646) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24447) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32249) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24608) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13562) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27239) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9125) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25266) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13806) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20480) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28216) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27587) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11309) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14415) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12647) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28719) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25644) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14600) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24598) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5759) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29422) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25464) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27781) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15967) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23771) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22714) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9036) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24050) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20395) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22633) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4548) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18900) * $signed(input_fmap_127[7:0]) +
	( 16'sd 20283) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27560) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22271) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19250) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5866) * $signed(input_fmap_132[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25470) * $signed(input_fmap_134[7:0]) +
	( 16'sd 29531) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8282) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13432) * $signed(input_fmap_137[7:0]) +
	( 15'sd 14754) * $signed(input_fmap_138[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_139[7:0]) +
	( 15'sd 11763) * $signed(input_fmap_140[7:0]) +
	( 14'sd 6680) * $signed(input_fmap_141[7:0]) +
	( 16'sd 29552) * $signed(input_fmap_142[7:0]) +
	( 16'sd 29385) * $signed(input_fmap_143[7:0]) +
	( 16'sd 23932) * $signed(input_fmap_144[7:0]) +
	( 14'sd 5899) * $signed(input_fmap_145[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30105) * $signed(input_fmap_147[7:0]) +
	( 15'sd 12230) * $signed(input_fmap_148[7:0]) +
	( 16'sd 16901) * $signed(input_fmap_149[7:0]) +
	( 16'sd 30192) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17709) * $signed(input_fmap_151[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11342) * $signed(input_fmap_153[7:0]) +
	( 16'sd 32714) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_155[7:0]) +
	( 15'sd 12202) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24080) * $signed(input_fmap_157[7:0]) +
	( 16'sd 21331) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6814) * $signed(input_fmap_159[7:0]) +
	( 14'sd 8144) * $signed(input_fmap_160[7:0]) +
	( 13'sd 3094) * $signed(input_fmap_161[7:0]) +
	( 16'sd 22063) * $signed(input_fmap_162[7:0]) +
	( 15'sd 11604) * $signed(input_fmap_163[7:0]) +
	( 14'sd 5496) * $signed(input_fmap_164[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_165[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_167[7:0]) +
	( 10'sd 351) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12016) * $signed(input_fmap_169[7:0]) +
	( 14'sd 6477) * $signed(input_fmap_170[7:0]) +
	( 16'sd 17359) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6654) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18386) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10726) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3418) * $signed(input_fmap_175[7:0]) +
	( 16'sd 17749) * $signed(input_fmap_176[7:0]) +
	( 15'sd 12130) * $signed(input_fmap_177[7:0]) +
	( 11'sd 1002) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18396) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_180[7:0]) +
	( 14'sd 5163) * $signed(input_fmap_181[7:0]) +
	( 12'sd 1121) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29359) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9901) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1685) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17793) * $signed(input_fmap_186[7:0]) +
	( 16'sd 29351) * $signed(input_fmap_187[7:0]) +
	( 16'sd 24314) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26021) * $signed(input_fmap_189[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24317) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15013) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26481) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18281) * $signed(input_fmap_194[7:0]) +
	( 14'sd 8089) * $signed(input_fmap_195[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_197[7:0]) +
	( 13'sd 3253) * $signed(input_fmap_198[7:0]) +
	( 16'sd 26442) * $signed(input_fmap_199[7:0]) +
	( 16'sd 28806) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6829) * $signed(input_fmap_201[7:0]) +
	( 15'sd 13431) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25294) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17825) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29739) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27606) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30481) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22961) * $signed(input_fmap_208[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1846) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30166) * $signed(input_fmap_211[7:0]) +
	( 15'sd 13727) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2436) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30013) * $signed(input_fmap_214[7:0]) +
	( 16'sd 19906) * $signed(input_fmap_215[7:0]) +
	( 16'sd 22618) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32238) * $signed(input_fmap_217[7:0]) +
	( 16'sd 25095) * $signed(input_fmap_218[7:0]) +
	( 13'sd 2830) * $signed(input_fmap_219[7:0]) +
	( 13'sd 2163) * $signed(input_fmap_220[7:0]) +
	( 16'sd 29117) * $signed(input_fmap_221[7:0]) +
	( 15'sd 9293) * $signed(input_fmap_222[7:0]) +
	( 16'sd 29103) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7224) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13543) * $signed(input_fmap_225[7:0]) +
	( 10'sd 292) * $signed(input_fmap_226[7:0]) +
	( 15'sd 16155) * $signed(input_fmap_227[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_228[7:0]) +
	( 13'sd 2774) * $signed(input_fmap_229[7:0]) +
	( 13'sd 2176) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18122) * $signed(input_fmap_231[7:0]) +
	( 12'sd 2027) * $signed(input_fmap_232[7:0]) +
	( 16'sd 26113) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23578) * $signed(input_fmap_234[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_235[7:0]) +
	( 16'sd 29265) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6871) * $signed(input_fmap_237[7:0]) +
	( 15'sd 10457) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31181) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29692) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27342) * $signed(input_fmap_242[7:0]) +
	( 16'sd 30676) * $signed(input_fmap_243[7:0]) +
	( 16'sd 31882) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3687) * $signed(input_fmap_245[7:0]) +
	( 14'sd 4765) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21056) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4475) * $signed(input_fmap_248[7:0]) +
	( 15'sd 13074) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30654) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14113) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20896) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_253[7:0]) +
	( 15'sd 12644) * $signed(input_fmap_254[7:0]) +
	( 15'sd 13180) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_110;
assign conv_mac_110 = 
	( 16'sd 17486) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2987) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21690) * $signed(input_fmap_2[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28532) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12033) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29033) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1203) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23509) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14112) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18600) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5230) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27875) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19479) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20845) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28502) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21563) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6745) * $signed(input_fmap_19[7:0]) +
	( 11'sd 849) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21023) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16249) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4358) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25712) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18206) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6754) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32473) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25693) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5482) * $signed(input_fmap_29[7:0]) +
	( 16'sd 28634) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18588) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25750) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6473) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8911) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5125) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24692) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25308) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10179) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5817) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20697) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17367) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6185) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19289) * $signed(input_fmap_44[7:0]) +
	( 10'sd 387) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12829) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26828) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7122) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2683) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23713) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13271) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18822) * $signed(input_fmap_52[7:0]) +
	( 11'sd 962) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15724) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27037) * $signed(input_fmap_55[7:0]) +
	( 16'sd 25831) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9664) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16200) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32311) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3169) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9902) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19712) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8936) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29439) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22136) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10445) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8511) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15913) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17106) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24146) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8590) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25072) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19114) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17877) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_78[7:0]) +
	( 9'sd 186) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30226) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8310) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5276) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13670) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31802) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23537) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21998) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25135) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7739) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10926) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27819) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29275) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9715) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25790) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27423) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7973) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8268) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29996) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19942) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5403) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9766) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27595) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25005) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17958) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17455) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31876) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27443) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14861) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27189) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25236) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30295) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18070) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5358) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32678) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20907) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19190) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8846) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17171) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13389) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1826) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25176) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19803) * $signed(input_fmap_126[7:0]) +
	( 10'sd 353) * $signed(input_fmap_127[7:0]) +
	( 14'sd 5927) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31188) * $signed(input_fmap_129[7:0]) +
	( 15'sd 15036) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_131[7:0]) +
	( 16'sd 26304) * $signed(input_fmap_132[7:0]) +
	( 16'sd 26520) * $signed(input_fmap_133[7:0]) +
	( 16'sd 26437) * $signed(input_fmap_134[7:0]) +
	( 16'sd 16981) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17437) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6608) * $signed(input_fmap_137[7:0]) +
	( 14'sd 5615) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21025) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9023) * $signed(input_fmap_140[7:0]) +
	( 12'sd 1031) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14636) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17997) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11883) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2302) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27632) * $signed(input_fmap_146[7:0]) +
	( 13'sd 2103) * $signed(input_fmap_147[7:0]) +
	( 14'sd 5485) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23433) * $signed(input_fmap_149[7:0]) +
	( 15'sd 13704) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4963) * $signed(input_fmap_151[7:0]) +
	( 14'sd 5797) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25296) * $signed(input_fmap_153[7:0]) +
	( 16'sd 26384) * $signed(input_fmap_154[7:0]) +
	( 16'sd 29367) * $signed(input_fmap_155[7:0]) +
	( 16'sd 31664) * $signed(input_fmap_156[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_157[7:0]) +
	( 14'sd 7801) * $signed(input_fmap_158[7:0]) +
	( 16'sd 29083) * $signed(input_fmap_159[7:0]) +
	( 13'sd 2955) * $signed(input_fmap_160[7:0]) +
	( 14'sd 6794) * $signed(input_fmap_161[7:0]) +
	( 16'sd 22657) * $signed(input_fmap_162[7:0]) +
	( 15'sd 14876) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11917) * $signed(input_fmap_164[7:0]) +
	( 16'sd 27621) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3351) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17792) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26564) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18453) * $signed(input_fmap_169[7:0]) +
	( 14'sd 6656) * $signed(input_fmap_170[7:0]) +
	( 16'sd 17515) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6991) * $signed(input_fmap_172[7:0]) +
	( 15'sd 16094) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10545) * $signed(input_fmap_174[7:0]) +
	( 15'sd 16244) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13945) * $signed(input_fmap_176[7:0]) +
	( 16'sd 17280) * $signed(input_fmap_177[7:0]) +
	( 14'sd 8025) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20923) * $signed(input_fmap_179[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_180[7:0]) +
	( 16'sd 24899) * $signed(input_fmap_181[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_182[7:0]) +
	( 15'sd 10632) * $signed(input_fmap_183[7:0]) +
	( 9'sd 254) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1873) * $signed(input_fmap_185[7:0]) +
	( 15'sd 10570) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1296) * $signed(input_fmap_187[7:0]) +
	( 16'sd 16748) * $signed(input_fmap_188[7:0]) +
	( 12'sd 1751) * $signed(input_fmap_189[7:0]) +
	( 16'sd 26627) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3263) * $signed(input_fmap_191[7:0]) +
	( 15'sd 16157) * $signed(input_fmap_192[7:0]) +
	( 16'sd 32432) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26636) * $signed(input_fmap_194[7:0]) +
	( 13'sd 2713) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20551) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24388) * $signed(input_fmap_197[7:0]) +
	( 16'sd 25594) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14456) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5505) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13050) * $signed(input_fmap_201[7:0]) +
	( 15'sd 10035) * $signed(input_fmap_202[7:0]) +
	( 11'sd 675) * $signed(input_fmap_203[7:0]) +
	( 14'sd 8081) * $signed(input_fmap_204[7:0]) +
	( 16'sd 17878) * $signed(input_fmap_205[7:0]) +
	( 15'sd 13982) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7066) * $signed(input_fmap_207[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26875) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5636) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23767) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29061) * $signed(input_fmap_212[7:0]) +
	( 16'sd 26531) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31225) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17293) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23968) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24596) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21540) * $signed(input_fmap_218[7:0]) +
	( 14'sd 7741) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22400) * $signed(input_fmap_220[7:0]) +
	( 14'sd 8164) * $signed(input_fmap_221[7:0]) +
	( 16'sd 30418) * $signed(input_fmap_222[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13264) * $signed(input_fmap_224[7:0]) +
	( 15'sd 10321) * $signed(input_fmap_225[7:0]) +
	( 16'sd 21224) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_228[7:0]) +
	( 15'sd 12119) * $signed(input_fmap_229[7:0]) +
	( 16'sd 20290) * $signed(input_fmap_230[7:0]) +
	( 16'sd 29949) * $signed(input_fmap_231[7:0]) +
	( 11'sd 771) * $signed(input_fmap_232[7:0]) +
	( 15'sd 9849) * $signed(input_fmap_233[7:0]) +
	( 16'sd 21582) * $signed(input_fmap_234[7:0]) +
	( 12'sd 1691) * $signed(input_fmap_235[7:0]) +
	( 16'sd 17743) * $signed(input_fmap_236[7:0]) +
	( 15'sd 16088) * $signed(input_fmap_237[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12637) * $signed(input_fmap_239[7:0]) +
	( 15'sd 15775) * $signed(input_fmap_240[7:0]) +
	( 16'sd 19437) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23359) * $signed(input_fmap_242[7:0]) +
	( 15'sd 14807) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_244[7:0]) +
	( 16'sd 20188) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22934) * $signed(input_fmap_246[7:0]) +
	( 14'sd 7224) * $signed(input_fmap_247[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_248[7:0]) +
	( 16'sd 27905) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26928) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_251[7:0]) +
	( 15'sd 14415) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17461) * $signed(input_fmap_253[7:0]) +
	( 16'sd 24650) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20273) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_111;
assign conv_mac_111 = 
	( 15'sd 12074) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17427) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25605) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21221) * $signed(input_fmap_5[7:0]) +
	( 10'sd 358) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2348) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30658) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23808) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15774) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29346) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14852) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14591) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18447) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31718) * $signed(input_fmap_16[7:0]) +
	( 11'sd 766) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13017) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25528) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5307) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16077) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22339) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11321) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17542) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13095) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17117) * $signed(input_fmap_26[7:0]) +
	( 11'sd 759) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21889) * $signed(input_fmap_28[7:0]) +
	( 11'sd 1023) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9303) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5702) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27146) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29724) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4858) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8794) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20345) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5490) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3925) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2311) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8412) * $signed(input_fmap_41[7:0]) +
	( 11'sd 798) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32443) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14677) * $signed(input_fmap_44[7:0]) +
	( 12'sd 2012) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22813) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16958) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15052) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13259) * $signed(input_fmap_50[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30708) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26432) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21591) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21602) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22860) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22964) * $signed(input_fmap_59[7:0]) +
	( 16'sd 21260) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29763) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14876) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11986) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30355) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11820) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7418) * $signed(input_fmap_66[7:0]) +
	( 12'sd 1283) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19609) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29844) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25835) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27159) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24862) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15634) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3531) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1792) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14303) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26380) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19543) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30061) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26965) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8418) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28929) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14859) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10700) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9373) * $signed(input_fmap_87[7:0]) +
	( 14'sd 4284) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29249) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7980) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14381) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25894) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17987) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5409) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3624) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30847) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13655) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9673) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31862) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27192) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22213) * $signed(input_fmap_105[7:0]) +
	( 5'sd 10) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15295) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8785) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23961) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3596) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6569) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25264) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2945) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6586) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30854) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_116[7:0]) +
	( 15'sd 16078) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19286) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13402) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6576) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31217) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21608) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21305) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_126[7:0]) +
	( 11'sd 793) * $signed(input_fmap_127[7:0]) +
	( 16'sd 25351) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27884) * $signed(input_fmap_129[7:0]) +
	( 15'sd 9008) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_131[7:0]) +
	( 16'sd 20885) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21791) * $signed(input_fmap_133[7:0]) +
	( 15'sd 13318) * $signed(input_fmap_134[7:0]) +
	( 13'sd 2050) * $signed(input_fmap_135[7:0]) +
	( 15'sd 10759) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27878) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7261) * $signed(input_fmap_138[7:0]) +
	( 16'sd 29682) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30960) * $signed(input_fmap_140[7:0]) +
	( 15'sd 8967) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31090) * $signed(input_fmap_142[7:0]) +
	( 15'sd 11460) * $signed(input_fmap_143[7:0]) +
	( 16'sd 21540) * $signed(input_fmap_144[7:0]) +
	( 15'sd 13250) * $signed(input_fmap_145[7:0]) +
	( 16'sd 26890) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18914) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11937) * $signed(input_fmap_148[7:0]) +
	( 16'sd 31917) * $signed(input_fmap_149[7:0]) +
	( 16'sd 19753) * $signed(input_fmap_150[7:0]) +
	( 13'sd 2628) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16832) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31459) * $signed(input_fmap_153[7:0]) +
	( 15'sd 15272) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17696) * $signed(input_fmap_156[7:0]) +
	( 10'sd 465) * $signed(input_fmap_157[7:0]) +
	( 16'sd 29652) * $signed(input_fmap_158[7:0]) +
	( 16'sd 25237) * $signed(input_fmap_159[7:0]) +
	( 15'sd 10569) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31952) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10669) * $signed(input_fmap_162[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_163[7:0]) +
	( 16'sd 21763) * $signed(input_fmap_164[7:0]) +
	( 16'sd 24455) * $signed(input_fmap_165[7:0]) +
	( 15'sd 11480) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17521) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12053) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_170[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_171[7:0]) +
	( 16'sd 28237) * $signed(input_fmap_172[7:0]) +
	( 9'sd 143) * $signed(input_fmap_173[7:0]) +
	( 13'sd 2654) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7743) * $signed(input_fmap_175[7:0]) +
	( 15'sd 14592) * $signed(input_fmap_176[7:0]) +
	( 10'sd 282) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9460) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18806) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26317) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30789) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2918) * $signed(input_fmap_183[7:0]) +
	( 14'sd 5321) * $signed(input_fmap_184[7:0]) +
	( 15'sd 9884) * $signed(input_fmap_185[7:0]) +
	( 16'sd 28026) * $signed(input_fmap_186[7:0]) +
	( 16'sd 26217) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21804) * $signed(input_fmap_188[7:0]) +
	( 16'sd 27813) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30318) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23516) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12031) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_193[7:0]) +
	( 15'sd 13396) * $signed(input_fmap_194[7:0]) +
	( 16'sd 20957) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25071) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10642) * $signed(input_fmap_197[7:0]) +
	( 16'sd 31411) * $signed(input_fmap_198[7:0]) +
	( 16'sd 31367) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3278) * $signed(input_fmap_200[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21135) * $signed(input_fmap_202[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14559) * $signed(input_fmap_204[7:0]) +
	( 15'sd 13637) * $signed(input_fmap_205[7:0]) +
	( 11'sd 867) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18510) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22302) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26084) * $signed(input_fmap_209[7:0]) +
	( 16'sd 26213) * $signed(input_fmap_210[7:0]) +
	( 16'sd 19047) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1766) * $signed(input_fmap_212[7:0]) +
	( 15'sd 14056) * $signed(input_fmap_213[7:0]) +
	( 9'sd 237) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1289) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23266) * $signed(input_fmap_216[7:0]) +
	( 14'sd 6882) * $signed(input_fmap_217[7:0]) +
	( 16'sd 24660) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21308) * $signed(input_fmap_219[7:0]) +
	( 16'sd 18874) * $signed(input_fmap_220[7:0]) +
	( 15'sd 9142) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12147) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2399) * $signed(input_fmap_223[7:0]) +
	( 16'sd 31657) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5379) * $signed(input_fmap_225[7:0]) +
	( 15'sd 9129) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20647) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31965) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6297) * $signed(input_fmap_229[7:0]) +
	( 15'sd 10642) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14710) * $signed(input_fmap_231[7:0]) +
	( 16'sd 24180) * $signed(input_fmap_232[7:0]) +
	( 16'sd 31310) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5814) * $signed(input_fmap_234[7:0]) +
	( 14'sd 6556) * $signed(input_fmap_235[7:0]) +
	( 14'sd 7274) * $signed(input_fmap_236[7:0]) +
	( 14'sd 4303) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22735) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12264) * $signed(input_fmap_239[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7150) * $signed(input_fmap_241[7:0]) +
	( 16'sd 32304) * $signed(input_fmap_242[7:0]) +
	( 16'sd 19030) * $signed(input_fmap_243[7:0]) +
	( 14'sd 8032) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10377) * $signed(input_fmap_245[7:0]) +
	( 14'sd 8133) * $signed(input_fmap_246[7:0]) +
	( 14'sd 5780) * $signed(input_fmap_247[7:0]) +
	( 16'sd 20700) * $signed(input_fmap_248[7:0]) +
	( 16'sd 16757) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30722) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13667) * $signed(input_fmap_251[7:0]) +
	( 16'sd 32213) * $signed(input_fmap_252[7:0]) +
	( 15'sd 16095) * $signed(input_fmap_253[7:0]) +
	( 16'sd 16984) * $signed(input_fmap_254[7:0]) +
	( 14'sd 4374) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_112;
assign conv_mac_112 = 
	( 16'sd 16450) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7544) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6417) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30908) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21172) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22056) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15194) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20811) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30521) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12411) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5132) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1958) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13863) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5919) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4813) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3967) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19161) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6309) * $signed(input_fmap_18[7:0]) +
	( 11'sd 834) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22107) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22503) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13399) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18962) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20716) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16617) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16679) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19009) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_30[7:0]) +
	( 9'sd 138) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10904) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16221) * $signed(input_fmap_33[7:0]) +
	( 10'sd 469) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23364) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32010) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3859) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19318) * $signed(input_fmap_38[7:0]) +
	( 8'sd 108) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7582) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4364) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30980) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10492) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20423) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3922) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3890) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5763) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15444) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16610) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3027) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22356) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7631) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14453) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21457) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17719) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18649) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29092) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12491) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29834) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11810) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15326) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7298) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24342) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1964) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31529) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21741) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25239) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20042) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4972) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12086) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23671) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30329) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8255) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27807) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30685) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25649) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14740) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_79[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22408) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11669) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6759) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24409) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24105) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17323) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9837) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28852) * $signed(input_fmap_90[7:0]) +
	( 14'sd 8026) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15498) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32506) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15209) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24991) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14428) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2173) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30524) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23852) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12584) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27211) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30073) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9628) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1699) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26753) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29562) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23879) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16064) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3862) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14403) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26671) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12579) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17650) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4989) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5413) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10098) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10435) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28493) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24328) * $signed(input_fmap_122[7:0]) +
	( 11'sd 609) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6939) * $signed(input_fmap_124[7:0]) +
	( 15'sd 8915) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23127) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19375) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8856) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1305) * $signed(input_fmap_129[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13389) * $signed(input_fmap_131[7:0]) +
	( 14'sd 4178) * $signed(input_fmap_132[7:0]) +
	( 14'sd 5904) * $signed(input_fmap_133[7:0]) +
	( 15'sd 10988) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19574) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23836) * $signed(input_fmap_136[7:0]) +
	( 12'sd 1136) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28580) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18600) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11339) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7192) * $signed(input_fmap_143[7:0]) +
	( 16'sd 32186) * $signed(input_fmap_144[7:0]) +
	( 15'sd 12344) * $signed(input_fmap_145[7:0]) +
	( 15'sd 11247) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19519) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3792) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4750) * $signed(input_fmap_149[7:0]) +
	( 16'sd 19126) * $signed(input_fmap_150[7:0]) +
	( 15'sd 9031) * $signed(input_fmap_151[7:0]) +
	( 15'sd 13763) * $signed(input_fmap_152[7:0]) +
	( 16'sd 26641) * $signed(input_fmap_153[7:0]) +
	( 16'sd 26245) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13101) * $signed(input_fmap_155[7:0]) +
	( 11'sd 856) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27396) * $signed(input_fmap_157[7:0]) +
	( 14'sd 6446) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5651) * $signed(input_fmap_159[7:0]) +
	( 16'sd 30751) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23974) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30190) * $signed(input_fmap_162[7:0]) +
	( 16'sd 29763) * $signed(input_fmap_163[7:0]) +
	( 15'sd 16272) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14077) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3498) * $signed(input_fmap_166[7:0]) +
	( 15'sd 15254) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6567) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17976) * $signed(input_fmap_170[7:0]) +
	( 15'sd 14824) * $signed(input_fmap_171[7:0]) +
	( 15'sd 10211) * $signed(input_fmap_172[7:0]) +
	( 15'sd 10536) * $signed(input_fmap_173[7:0]) +
	( 6'sd 19) * $signed(input_fmap_174[7:0]) +
	( 14'sd 6623) * $signed(input_fmap_175[7:0]) +
	( 15'sd 9094) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6929) * $signed(input_fmap_177[7:0]) +
	( 16'sd 19731) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_179[7:0]) +
	( 13'sd 2763) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15131) * $signed(input_fmap_181[7:0]) +
	( 16'sd 25593) * $signed(input_fmap_182[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22493) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27622) * $signed(input_fmap_185[7:0]) +
	( 16'sd 30828) * $signed(input_fmap_186[7:0]) +
	( 16'sd 20020) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21673) * $signed(input_fmap_188[7:0]) +
	( 15'sd 12269) * $signed(input_fmap_189[7:0]) +
	( 15'sd 16273) * $signed(input_fmap_190[7:0]) +
	( 15'sd 10034) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12360) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27075) * $signed(input_fmap_193[7:0]) +
	( 6'sd 21) * $signed(input_fmap_194[7:0]) +
	( 14'sd 4424) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12316) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14913) * $signed(input_fmap_197[7:0]) +
	( 15'sd 14866) * $signed(input_fmap_198[7:0]) +
	( 16'sd 16752) * $signed(input_fmap_199[7:0]) +
	( 16'sd 30646) * $signed(input_fmap_200[7:0]) +
	( 15'sd 16184) * $signed(input_fmap_201[7:0]) +
	( 16'sd 27793) * $signed(input_fmap_202[7:0]) +
	( 11'sd 620) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11148) * $signed(input_fmap_204[7:0]) +
	( 16'sd 23864) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12694) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3889) * $signed(input_fmap_207[7:0]) +
	( 15'sd 10306) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23383) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9310) * $signed(input_fmap_210[7:0]) +
	( 16'sd 24693) * $signed(input_fmap_211[7:0]) +
	( 13'sd 2690) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24067) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1616) * $signed(input_fmap_214[7:0]) +
	( 16'sd 31424) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20480) * $signed(input_fmap_216[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31552) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14723) * $signed(input_fmap_219[7:0]) +
	( 16'sd 32620) * $signed(input_fmap_220[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_221[7:0]) +
	( 15'sd 11442) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22434) * $signed(input_fmap_223[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_224[7:0]) +
	( 11'sd 689) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30142) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24439) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8640) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17824) * $signed(input_fmap_229[7:0]) +
	( 15'sd 12036) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13047) * $signed(input_fmap_231[7:0]) +
	( 15'sd 10671) * $signed(input_fmap_232[7:0]) +
	( 16'sd 19135) * $signed(input_fmap_233[7:0]) +
	( 16'sd 27986) * $signed(input_fmap_234[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12896) * $signed(input_fmap_236[7:0]) +
	( 16'sd 31281) * $signed(input_fmap_237[7:0]) +
	( 15'sd 15560) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9768) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19154) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3146) * $signed(input_fmap_241[7:0]) +
	( 15'sd 12077) * $signed(input_fmap_242[7:0]) +
	( 16'sd 21882) * $signed(input_fmap_243[7:0]) +
	( 16'sd 26668) * $signed(input_fmap_244[7:0]) +
	( 15'sd 15251) * $signed(input_fmap_245[7:0]) +
	( 14'sd 6704) * $signed(input_fmap_246[7:0]) +
	( 16'sd 23255) * $signed(input_fmap_247[7:0]) +
	( 16'sd 20842) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3443) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6656) * $signed(input_fmap_251[7:0]) +
	( 16'sd 25967) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13169) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26460) * $signed(input_fmap_254[7:0]) +
	( 16'sd 30281) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_113;
assign conv_mac_113 = 
	( 16'sd 31485) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26314) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31212) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5293) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17413) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12495) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20595) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15194) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12770) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21898) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5173) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31759) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24813) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19346) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14536) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30875) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27522) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22069) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3632) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18107) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15625) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2281) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21136) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26201) * $signed(input_fmap_25[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18346) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27661) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26679) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20704) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26590) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23667) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18338) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18866) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3326) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26007) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5093) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21269) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8476) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7755) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11704) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12398) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2095) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16667) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1627) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4643) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17254) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21482) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2246) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7966) * $signed(input_fmap_52[7:0]) +
	( 11'sd 778) * $signed(input_fmap_53[7:0]) +
	( 13'sd 4029) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25520) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2410) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31859) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4104) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12799) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19769) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11113) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7834) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29095) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24090) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2455) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29152) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15038) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27895) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21503) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19545) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20166) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31612) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31837) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30461) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15332) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19196) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12108) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11786) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16864) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29762) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32076) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18408) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27619) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19420) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31664) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6354) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7670) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23186) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32125) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23373) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24121) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17633) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21429) * $signed(input_fmap_97[7:0]) +
	( 16'sd 16705) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16302) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10984) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8853) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16467) * $signed(input_fmap_102[7:0]) +
	( 11'sd 764) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7485) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27413) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9594) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11063) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25571) * $signed(input_fmap_109[7:0]) +
	( 11'sd 579) * $signed(input_fmap_110[7:0]) +
	( 14'sd 8047) * $signed(input_fmap_111[7:0]) +
	( 10'sd 307) * $signed(input_fmap_112[7:0]) +
	( 11'sd 906) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3018) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15383) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14406) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26783) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3398) * $signed(input_fmap_118[7:0]) +
	( 10'sd 439) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26255) * $signed(input_fmap_120[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13695) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19037) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29624) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9699) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26284) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4826) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5479) * $signed(input_fmap_129[7:0]) +
	( 15'sd 11774) * $signed(input_fmap_130[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_131[7:0]) +
	( 15'sd 9704) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29776) * $signed(input_fmap_133[7:0]) +
	( 15'sd 12198) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32303) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15273) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24186) * $signed(input_fmap_137[7:0]) +
	( 16'sd 18411) * $signed(input_fmap_138[7:0]) +
	( 12'sd 1279) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15317) * $signed(input_fmap_140[7:0]) +
	( 16'sd 23276) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8727) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7019) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_144[7:0]) +
	( 16'sd 16402) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18459) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11516) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_148[7:0]) +
	( 16'sd 30231) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31261) * $signed(input_fmap_150[7:0]) +
	( 15'sd 8949) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22491) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24488) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24280) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13143) * $signed(input_fmap_155[7:0]) +
	( 14'sd 4737) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20134) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20446) * $signed(input_fmap_158[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5954) * $signed(input_fmap_160[7:0]) +
	( 16'sd 26992) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_163[7:0]) +
	( 16'sd 29117) * $signed(input_fmap_164[7:0]) +
	( 14'sd 8176) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3529) * $signed(input_fmap_166[7:0]) +
	( 16'sd 27972) * $signed(input_fmap_167[7:0]) +
	( 16'sd 28190) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7901) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12918) * $signed(input_fmap_171[7:0]) +
	( 16'sd 17782) * $signed(input_fmap_172[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19770) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1422) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13579) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1509) * $signed(input_fmap_177[7:0]) +
	( 16'sd 25403) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2904) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24001) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23350) * $signed(input_fmap_181[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25605) * $signed(input_fmap_183[7:0]) +
	( 16'sd 29312) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24414) * $signed(input_fmap_185[7:0]) +
	( 16'sd 24574) * $signed(input_fmap_186[7:0]) +
	( 16'sd 21449) * $signed(input_fmap_187[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30745) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28495) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32037) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28357) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28533) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9768) * $signed(input_fmap_194[7:0]) +
	( 14'sd 6574) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15034) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5366) * $signed(input_fmap_198[7:0]) +
	( 16'sd 18967) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13775) * $signed(input_fmap_200[7:0]) +
	( 12'sd 2020) * $signed(input_fmap_201[7:0]) +
	( 15'sd 9154) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5911) * $signed(input_fmap_203[7:0]) +
	( 11'sd 981) * $signed(input_fmap_204[7:0]) +
	( 16'sd 27949) * $signed(input_fmap_205[7:0]) +
	( 12'sd 2047) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17127) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8600) * $signed(input_fmap_208[7:0]) +
	( 16'sd 21081) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9164) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3731) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1727) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9919) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31076) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6813) * $signed(input_fmap_215[7:0]) +
	( 16'sd 27496) * $signed(input_fmap_216[7:0]) +
	( 15'sd 12824) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5313) * $signed(input_fmap_218[7:0]) +
	( 16'sd 22066) * $signed(input_fmap_219[7:0]) +
	( 16'sd 32032) * $signed(input_fmap_220[7:0]) +
	( 15'sd 11539) * $signed(input_fmap_221[7:0]) +
	( 12'sd 1197) * $signed(input_fmap_222[7:0]) +
	( 15'sd 13125) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14589) * $signed(input_fmap_224[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_225[7:0]) +
	( 11'sd 691) * $signed(input_fmap_226[7:0]) +
	( 11'sd 571) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25411) * $signed(input_fmap_228[7:0]) +
	( 15'sd 15577) * $signed(input_fmap_229[7:0]) +
	( 16'sd 19936) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24657) * $signed(input_fmap_231[7:0]) +
	( 16'sd 19014) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5476) * $signed(input_fmap_233[7:0]) +
	( 16'sd 22348) * $signed(input_fmap_234[7:0]) +
	( 13'sd 4041) * $signed(input_fmap_235[7:0]) +
	( 16'sd 29593) * $signed(input_fmap_236[7:0]) +
	( 16'sd 21409) * $signed(input_fmap_237[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21487) * $signed(input_fmap_239[7:0]) +
	( 16'sd 27118) * $signed(input_fmap_240[7:0]) +
	( 16'sd 22946) * $signed(input_fmap_241[7:0]) +
	( 15'sd 8267) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25776) * $signed(input_fmap_243[7:0]) +
	( 15'sd 11613) * $signed(input_fmap_244[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15503) * $signed(input_fmap_246[7:0]) +
	( 16'sd 28698) * $signed(input_fmap_247[7:0]) +
	( 15'sd 9593) * $signed(input_fmap_248[7:0]) +
	( 16'sd 23470) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7518) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6199) * $signed(input_fmap_251[7:0]) +
	( 16'sd 16385) * $signed(input_fmap_252[7:0]) +
	( 16'sd 21409) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1340) * $signed(input_fmap_254[7:0]) +
	( 16'sd 31703) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_114;
assign conv_mac_114 = 
	( 15'sd 15889) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32698) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27703) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20793) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22418) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20661) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16056) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4341) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21410) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21440) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22412) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9130) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4995) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3781) * $signed(input_fmap_13[7:0]) +
	( 10'sd 310) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23274) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4526) * $signed(input_fmap_18[7:0]) +
	( 14'sd 8022) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24974) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_22[7:0]) +
	( 14'sd 8008) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25325) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5039) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31430) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27193) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14165) * $signed(input_fmap_30[7:0]) +
	( 13'sd 4027) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12752) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26889) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23624) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2305) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1113) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13354) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21183) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26458) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3026) * $signed(input_fmap_42[7:0]) +
	( 14'sd 8153) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1040) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19750) * $signed(input_fmap_46[7:0]) +
	( 11'sd 900) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25571) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23053) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7872) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6966) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32507) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12590) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29442) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26647) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5290) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8167) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25521) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24005) * $signed(input_fmap_59[7:0]) +
	( 16'sd 16753) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8336) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21022) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7409) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14917) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25278) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21362) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32666) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11971) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3233) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7990) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28581) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4799) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19328) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7824) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22514) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12533) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24550) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28273) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8671) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7134) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3770) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11794) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25095) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13925) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10786) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30399) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8997) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3520) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16330) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14955) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2205) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23764) * $signed(input_fmap_96[7:0]) +
	( 10'sd 284) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3086) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5039) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2498) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6433) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18611) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19743) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31263) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1986) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30590) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11312) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11826) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6165) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17002) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13337) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18513) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27783) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1434) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21308) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31096) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14981) * $signed(input_fmap_118[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14275) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24798) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23261) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30999) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2256) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1917) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6636) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29695) * $signed(input_fmap_128[7:0]) +
	( 16'sd 16576) * $signed(input_fmap_129[7:0]) +
	( 13'sd 3586) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_131[7:0]) +
	( 11'sd 641) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31270) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_134[7:0]) +
	( 12'sd 1497) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25506) * $signed(input_fmap_136[7:0]) +
	( 14'sd 5611) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7311) * $signed(input_fmap_138[7:0]) +
	( 16'sd 26705) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17558) * $signed(input_fmap_140[7:0]) +
	( 15'sd 14353) * $signed(input_fmap_141[7:0]) +
	( 12'sd 1120) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4920) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6159) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26212) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21564) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9304) * $signed(input_fmap_147[7:0]) +
	( 15'sd 12099) * $signed(input_fmap_148[7:0]) +
	( 14'sd 5288) * $signed(input_fmap_149[7:0]) +
	( 13'sd 3007) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6389) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14328) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24818) * $signed(input_fmap_153[7:0]) +
	( 16'sd 28083) * $signed(input_fmap_154[7:0]) +
	( 11'sd 689) * $signed(input_fmap_155[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_156[7:0]) +
	( 16'sd 19754) * $signed(input_fmap_157[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14813) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_160[7:0]) +
	( 16'sd 18114) * $signed(input_fmap_161[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_162[7:0]) +
	( 16'sd 25586) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13602) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12323) * $signed(input_fmap_165[7:0]) +
	( 16'sd 23937) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7097) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20983) * $signed(input_fmap_168[7:0]) +
	( 15'sd 8507) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14137) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20420) * $signed(input_fmap_171[7:0]) +
	( 15'sd 16242) * $signed(input_fmap_172[7:0]) +
	( 13'sd 2198) * $signed(input_fmap_173[7:0]) +
	( 16'sd 18576) * $signed(input_fmap_174[7:0]) +
	( 16'sd 31070) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1765) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30519) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10726) * $signed(input_fmap_178[7:0]) +
	( 16'sd 17478) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21123) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18739) * $signed(input_fmap_181[7:0]) +
	( 16'sd 20387) * $signed(input_fmap_182[7:0]) +
	( 10'sd 493) * $signed(input_fmap_183[7:0]) +
	( 14'sd 5652) * $signed(input_fmap_184[7:0]) +
	( 15'sd 12706) * $signed(input_fmap_185[7:0]) +
	( 11'sd 576) * $signed(input_fmap_186[7:0]) +
	( 14'sd 6894) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17071) * $signed(input_fmap_188[7:0]) +
	( 16'sd 27416) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4887) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23634) * $signed(input_fmap_191[7:0]) +
	( 9'sd 135) * $signed(input_fmap_192[7:0]) +
	( 13'sd 2794) * $signed(input_fmap_193[7:0]) +
	( 16'sd 20214) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24392) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19267) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11032) * $signed(input_fmap_197[7:0]) +
	( 14'sd 7076) * $signed(input_fmap_198[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_199[7:0]) +
	( 15'sd 9965) * $signed(input_fmap_200[7:0]) +
	( 16'sd 23339) * $signed(input_fmap_201[7:0]) +
	( 15'sd 13324) * $signed(input_fmap_202[7:0]) +
	( 16'sd 22930) * $signed(input_fmap_203[7:0]) +
	( 16'sd 31369) * $signed(input_fmap_204[7:0]) +
	( 16'sd 20328) * $signed(input_fmap_205[7:0]) +
	( 11'sd 954) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12530) * $signed(input_fmap_207[7:0]) +
	( 16'sd 24720) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18616) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12820) * $signed(input_fmap_211[7:0]) +
	( 14'sd 4544) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24895) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20321) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2256) * $signed(input_fmap_215[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17993) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26921) * $signed(input_fmap_218[7:0]) +
	( 16'sd 16636) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19395) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23817) * $signed(input_fmap_221[7:0]) +
	( 16'sd 24671) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19864) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12137) * $signed(input_fmap_224[7:0]) +
	( 16'sd 29392) * $signed(input_fmap_225[7:0]) +
	( 15'sd 12735) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27758) * $signed(input_fmap_227[7:0]) +
	( 16'sd 23571) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3916) * $signed(input_fmap_229[7:0]) +
	( 16'sd 25381) * $signed(input_fmap_230[7:0]) +
	( 15'sd 12454) * $signed(input_fmap_231[7:0]) +
	( 16'sd 28557) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5642) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15439) * $signed(input_fmap_234[7:0]) +
	( 15'sd 13033) * $signed(input_fmap_235[7:0]) +
	( 12'sd 1088) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2956) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28513) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21277) * $signed(input_fmap_239[7:0]) +
	( 16'sd 32444) * $signed(input_fmap_240[7:0]) +
	( 16'sd 22907) * $signed(input_fmap_241[7:0]) +
	( 15'sd 10495) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23704) * $signed(input_fmap_243[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_244[7:0]) +
	( 16'sd 23709) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23496) * $signed(input_fmap_246[7:0]) +
	( 15'sd 10771) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4381) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30039) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24540) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21211) * $signed(input_fmap_251[7:0]) +
	( 15'sd 8838) * $signed(input_fmap_252[7:0]) +
	( 16'sd 19704) * $signed(input_fmap_253[7:0]) +
	( 16'sd 24172) * $signed(input_fmap_254[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_115;
assign conv_mac_115 = 
	( 5'sd 15) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24881) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18135) * $signed(input_fmap_2[7:0]) +
	( 8'sd 123) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7392) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25493) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23400) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9205) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21617) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31059) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28882) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11626) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20011) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9354) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25223) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31262) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1523) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3833) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18508) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12284) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16912) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31618) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25607) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15554) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19279) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25266) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13811) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26343) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24967) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3541) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26759) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17266) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13050) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18044) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8172) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24496) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30761) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1513) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5806) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29410) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27925) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28686) * $signed(input_fmap_53[7:0]) +
	( 10'sd 375) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9985) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2579) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31003) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16626) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2393) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13246) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28779) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31184) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6912) * $signed(input_fmap_65[7:0]) +
	( 10'sd 413) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3472) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29500) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10933) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2157) * $signed(input_fmap_70[7:0]) +
	( 11'sd 587) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29765) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11971) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15301) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17707) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11036) * $signed(input_fmap_76[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19996) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4647) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10004) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22825) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29342) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30560) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31681) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32737) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15923) * $signed(input_fmap_88[7:0]) +
	( 15'sd 11645) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15191) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30779) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17871) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31882) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25992) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27531) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8547) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15371) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30420) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22520) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19632) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31749) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4309) * $signed(input_fmap_102[7:0]) +
	( 10'sd 467) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16391) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9621) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21190) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15367) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15044) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8654) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21066) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14420) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29243) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29692) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2397) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9382) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16262) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30237) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30013) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5598) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6002) * $signed(input_fmap_120[7:0]) +
	( 16'sd 21667) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14738) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6376) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5232) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18350) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15563) * $signed(input_fmap_128[7:0]) +
	( 11'sd 1009) * $signed(input_fmap_129[7:0]) +
	( 14'sd 4138) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5238) * $signed(input_fmap_131[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_132[7:0]) +
	( 16'sd 32398) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24284) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_135[7:0]) +
	( 13'sd 4065) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24972) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19020) * $signed(input_fmap_138[7:0]) +
	( 14'sd 8005) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3188) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24227) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25557) * $signed(input_fmap_142[7:0]) +
	( 16'sd 21020) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8944) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14150) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24051) * $signed(input_fmap_147[7:0]) +
	( 14'sd 8157) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18004) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23163) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18812) * $signed(input_fmap_151[7:0]) +
	( 16'sd 26886) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22398) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27744) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28880) * $signed(input_fmap_156[7:0]) +
	( 15'sd 10385) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20407) * $signed(input_fmap_158[7:0]) +
	( 16'sd 29881) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24814) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4223) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24093) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26704) * $signed(input_fmap_163[7:0]) +
	( 16'sd 32436) * $signed(input_fmap_164[7:0]) +
	( 15'sd 16124) * $signed(input_fmap_165[7:0]) +
	( 11'sd 512) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31087) * $signed(input_fmap_167[7:0]) +
	( 16'sd 32540) * $signed(input_fmap_168[7:0]) +
	( 13'sd 2942) * $signed(input_fmap_169[7:0]) +
	( 14'sd 6475) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19177) * $signed(input_fmap_171[7:0]) +
	( 16'sd 32400) * $signed(input_fmap_172[7:0]) +
	( 16'sd 24814) * $signed(input_fmap_173[7:0]) +
	( 16'sd 31105) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25819) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27944) * $signed(input_fmap_176[7:0]) +
	( 16'sd 26019) * $signed(input_fmap_177[7:0]) +
	( 16'sd 24721) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2840) * $signed(input_fmap_179[7:0]) +
	( 15'sd 9299) * $signed(input_fmap_180[7:0]) +
	( 10'sd 426) * $signed(input_fmap_181[7:0]) +
	( 16'sd 18431) * $signed(input_fmap_182[7:0]) +
	( 15'sd 9066) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26696) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26380) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3022) * $signed(input_fmap_186[7:0]) +
	( 11'sd 572) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_188[7:0]) +
	( 16'sd 22553) * $signed(input_fmap_189[7:0]) +
	( 16'sd 32056) * $signed(input_fmap_190[7:0]) +
	( 14'sd 4807) * $signed(input_fmap_191[7:0]) +
	( 14'sd 4702) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27128) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14348) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29235) * $signed(input_fmap_195[7:0]) +
	( 16'sd 21510) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25674) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22557) * $signed(input_fmap_198[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_199[7:0]) +
	( 12'sd 1091) * $signed(input_fmap_200[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_201[7:0]) +
	( 16'sd 30357) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5414) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5744) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24142) * $signed(input_fmap_205[7:0]) +
	( 15'sd 14568) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1756) * $signed(input_fmap_207[7:0]) +
	( 9'sd 219) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24807) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9834) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17885) * $signed(input_fmap_211[7:0]) +
	( 15'sd 8467) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2862) * $signed(input_fmap_213[7:0]) +
	( 14'sd 6919) * $signed(input_fmap_214[7:0]) +
	( 9'sd 197) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11921) * $signed(input_fmap_216[7:0]) +
	( 15'sd 15381) * $signed(input_fmap_217[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12619) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26289) * $signed(input_fmap_220[7:0]) +
	( 15'sd 11752) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19564) * $signed(input_fmap_222[7:0]) +
	( 16'sd 23961) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19645) * $signed(input_fmap_224[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11005) * $signed(input_fmap_226[7:0]) +
	( 16'sd 18817) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22933) * $signed(input_fmap_228[7:0]) +
	( 16'sd 31265) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7075) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28015) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7038) * $signed(input_fmap_232[7:0]) +
	( 16'sd 29516) * $signed(input_fmap_233[7:0]) +
	( 15'sd 10330) * $signed(input_fmap_234[7:0]) +
	( 16'sd 17437) * $signed(input_fmap_235[7:0]) +
	( 16'sd 24138) * $signed(input_fmap_236[7:0]) +
	( 16'sd 21018) * $signed(input_fmap_237[7:0]) +
	( 16'sd 21005) * $signed(input_fmap_238[7:0]) +
	( 14'sd 4550) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23945) * $signed(input_fmap_241[7:0]) +
	( 15'sd 9197) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23515) * $signed(input_fmap_243[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_244[7:0]) +
	( 15'sd 15291) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17784) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17448) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3704) * $signed(input_fmap_248[7:0]) +
	( 12'sd 1767) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7871) * $signed(input_fmap_250[7:0]) +
	( 10'sd 379) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13792) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_253[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_254[7:0]) +
	( 16'sd 21470) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_116;
assign conv_mac_116 = 
	( 16'sd 21934) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5836) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12185) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25827) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11717) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_6[7:0]) +
	( 13'sd 2963) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15807) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11765) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10224) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13461) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23323) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4334) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3506) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5760) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2391) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20870) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10624) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31321) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32055) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15974) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24681) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4101) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11108) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1583) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17588) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12419) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26984) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3921) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14992) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24666) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15725) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10624) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15184) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31868) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13035) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25477) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3116) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2903) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17003) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32205) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13119) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22259) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28642) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19162) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31341) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16475) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14976) * $signed(input_fmap_56[7:0]) +
	( 7'sd 41) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19360) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7772) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6444) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25755) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14579) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17940) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31756) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25250) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18410) * $signed(input_fmap_66[7:0]) +
	( 16'sd 20515) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10083) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12021) * $signed(input_fmap_69[7:0]) +
	( 11'sd 822) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17577) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30565) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6006) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8906) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20299) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17821) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21301) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23737) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31583) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20890) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17667) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27707) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17283) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4464) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29350) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2853) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9024) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21317) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18174) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32583) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13062) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16159) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19163) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29050) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30424) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28462) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24036) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14784) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12295) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15955) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19652) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11989) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1423) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24480) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20061) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15880) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12400) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24049) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27197) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_118[7:0]) +
	( 10'sd 269) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17555) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20766) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6527) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31492) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29400) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26291) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21535) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27790) * $signed(input_fmap_127[7:0]) +
	( 14'sd 5219) * $signed(input_fmap_128[7:0]) +
	( 14'sd 4785) * $signed(input_fmap_129[7:0]) +
	( 15'sd 15565) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19494) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18764) * $signed(input_fmap_132[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24083) * $signed(input_fmap_134[7:0]) +
	( 16'sd 29845) * $signed(input_fmap_135[7:0]) +
	( 16'sd 29804) * $signed(input_fmap_136[7:0]) +
	( 16'sd 32569) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17469) * $signed(input_fmap_138[7:0]) +
	( 16'sd 19015) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26487) * $signed(input_fmap_140[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_141[7:0]) +
	( 15'sd 9597) * $signed(input_fmap_142[7:0]) +
	( 16'sd 18587) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9595) * $signed(input_fmap_144[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24400) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4624) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2049) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18055) * $signed(input_fmap_150[7:0]) +
	( 14'sd 7230) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20883) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10762) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6321) * $signed(input_fmap_154[7:0]) +
	( 14'sd 4732) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24445) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25544) * $signed(input_fmap_157[7:0]) +
	( 15'sd 10292) * $signed(input_fmap_158[7:0]) +
	( 15'sd 10653) * $signed(input_fmap_159[7:0]) +
	( 11'sd 588) * $signed(input_fmap_160[7:0]) +
	( 14'sd 5749) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14659) * $signed(input_fmap_162[7:0]) +
	( 10'sd 306) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8597) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12454) * $signed(input_fmap_165[7:0]) +
	( 15'sd 10154) * $signed(input_fmap_166[7:0]) +
	( 15'sd 12077) * $signed(input_fmap_167[7:0]) +
	( 16'sd 18958) * $signed(input_fmap_168[7:0]) +
	( 14'sd 5978) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24532) * $signed(input_fmap_171[7:0]) +
	( 14'sd 5798) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19470) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6734) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25089) * $signed(input_fmap_175[7:0]) +
	( 16'sd 28747) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31730) * $signed(input_fmap_177[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_178[7:0]) +
	( 15'sd 10013) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27846) * $signed(input_fmap_180[7:0]) +
	( 15'sd 9272) * $signed(input_fmap_181[7:0]) +
	( 15'sd 16134) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29788) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11613) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_185[7:0]) +
	( 16'sd 31425) * $signed(input_fmap_186[7:0]) +
	( 10'sd 438) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21251) * $signed(input_fmap_188[7:0]) +
	( 15'sd 14325) * $signed(input_fmap_189[7:0]) +
	( 16'sd 19067) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19150) * $signed(input_fmap_191[7:0]) +
	( 13'sd 3320) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12939) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3341) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29452) * $signed(input_fmap_195[7:0]) +
	( 15'sd 8637) * $signed(input_fmap_196[7:0]) +
	( 16'sd 29278) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10970) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24127) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6619) * $signed(input_fmap_200[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_201[7:0]) +
	( 16'sd 24145) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6239) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2193) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_205[7:0]) +
	( 14'sd 7365) * $signed(input_fmap_206[7:0]) +
	( 15'sd 16049) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17326) * $signed(input_fmap_208[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31566) * $signed(input_fmap_210[7:0]) +
	( 16'sd 27744) * $signed(input_fmap_211[7:0]) +
	( 15'sd 9910) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23137) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1433) * $signed(input_fmap_214[7:0]) +
	( 16'sd 24629) * $signed(input_fmap_215[7:0]) +
	( 16'sd 29164) * $signed(input_fmap_216[7:0]) +
	( 16'sd 23881) * $signed(input_fmap_217[7:0]) +
	( 14'sd 6591) * $signed(input_fmap_218[7:0]) +
	( 15'sd 11165) * $signed(input_fmap_219[7:0]) +
	( 15'sd 11048) * $signed(input_fmap_220[7:0]) +
	( 16'sd 18598) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15685) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2817) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12283) * $signed(input_fmap_224[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_225[7:0]) +
	( 15'sd 8921) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27838) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_229[7:0]) +
	( 16'sd 19156) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13417) * $signed(input_fmap_231[7:0]) +
	( 16'sd 26082) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23380) * $signed(input_fmap_233[7:0]) +
	( 16'sd 26216) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19946) * $signed(input_fmap_235[7:0]) +
	( 16'sd 18458) * $signed(input_fmap_236[7:0]) +
	( 15'sd 15412) * $signed(input_fmap_237[7:0]) +
	( 16'sd 32150) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5086) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26761) * $signed(input_fmap_240[7:0]) +
	( 15'sd 12188) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1067) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31295) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20100) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24114) * $signed(input_fmap_245[7:0]) +
	( 14'sd 6864) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_247[7:0]) +
	( 16'sd 23864) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21590) * $signed(input_fmap_249[7:0]) +
	( 15'sd 8855) * $signed(input_fmap_250[7:0]) +
	( 16'sd 29123) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6994) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25717) * $signed(input_fmap_253[7:0]) +
	( 15'sd 11869) * $signed(input_fmap_254[7:0]) +
	( 14'sd 6347) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_117;
assign conv_mac_117 = 
	( 16'sd 23042) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2917) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24833) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26390) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10115) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24769) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7093) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21624) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23320) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1839) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1980) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29497) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26758) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18882) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14488) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7119) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3202) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11091) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20209) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16030) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28447) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32133) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22957) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15954) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30733) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21414) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10991) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22533) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21695) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21622) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26126) * $signed(input_fmap_35[7:0]) +
	( 11'sd 662) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16824) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32478) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15910) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19118) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21900) * $signed(input_fmap_42[7:0]) +
	( 11'sd 691) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20711) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18719) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2748) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11892) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6668) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9876) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17767) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29368) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3184) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15581) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16184) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10271) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18834) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24078) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15589) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23538) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4307) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2921) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11626) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3586) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23034) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2281) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8867) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2429) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26459) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31484) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20251) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25462) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14139) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23286) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8957) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27746) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13535) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15026) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22721) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1207) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1029) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25685) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5985) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22980) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31793) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11370) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27884) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20496) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4277) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18746) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19042) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14116) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6611) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11904) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29079) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20412) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24148) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14241) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31643) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13645) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7940) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10283) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31816) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28845) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16512) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21598) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6541) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32397) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27827) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14210) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3151) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9397) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11847) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3257) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7803) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10460) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32027) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5543) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9674) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29664) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8500) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7950) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22510) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19593) * $signed(input_fmap_131[7:0]) +
	( 16'sd 24555) * $signed(input_fmap_132[7:0]) +
	( 14'sd 5914) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21171) * $signed(input_fmap_134[7:0]) +
	( 15'sd 9667) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12490) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4443) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17445) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20464) * $signed(input_fmap_139[7:0]) +
	( 16'sd 32397) * $signed(input_fmap_140[7:0]) +
	( 16'sd 32492) * $signed(input_fmap_141[7:0]) +
	( 15'sd 10012) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10274) * $signed(input_fmap_143[7:0]) +
	( 15'sd 10875) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7307) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3908) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14720) * $signed(input_fmap_147[7:0]) +
	( 15'sd 12382) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2193) * $signed(input_fmap_149[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23625) * $signed(input_fmap_151[7:0]) +
	( 14'sd 4564) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1331) * $signed(input_fmap_153[7:0]) +
	( 16'sd 20428) * $signed(input_fmap_154[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15780) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24611) * $signed(input_fmap_157[7:0]) +
	( 16'sd 22576) * $signed(input_fmap_158[7:0]) +
	( 16'sd 31337) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5708) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4483) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13040) * $signed(input_fmap_162[7:0]) +
	( 15'sd 13685) * $signed(input_fmap_163[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_164[7:0]) +
	( 16'sd 20664) * $signed(input_fmap_165[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_166[7:0]) +
	( 15'sd 16082) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29786) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6238) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2757) * $signed(input_fmap_170[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_171[7:0]) +
	( 16'sd 20192) * $signed(input_fmap_172[7:0]) +
	( 15'sd 11481) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10932) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21490) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7156) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5936) * $signed(input_fmap_177[7:0]) +
	( 16'sd 29024) * $signed(input_fmap_178[7:0]) +
	( 16'sd 27790) * $signed(input_fmap_179[7:0]) +
	( 13'sd 2150) * $signed(input_fmap_180[7:0]) +
	( 16'sd 22848) * $signed(input_fmap_181[7:0]) +
	( 16'sd 31256) * $signed(input_fmap_182[7:0]) +
	( 16'sd 28858) * $signed(input_fmap_183[7:0]) +
	( 14'sd 6769) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7629) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4910) * $signed(input_fmap_186[7:0]) +
	( 14'sd 6808) * $signed(input_fmap_187[7:0]) +
	( 14'sd 8030) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3716) * $signed(input_fmap_189[7:0]) +
	( 16'sd 18015) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32473) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14508) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30622) * $signed(input_fmap_193[7:0]) +
	( 15'sd 10661) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13092) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11683) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31298) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2315) * $signed(input_fmap_198[7:0]) +
	( 13'sd 3652) * $signed(input_fmap_199[7:0]) +
	( 14'sd 7311) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12358) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21332) * $signed(input_fmap_202[7:0]) +
	( 16'sd 23090) * $signed(input_fmap_203[7:0]) +
	( 16'sd 20428) * $signed(input_fmap_204[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_205[7:0]) +
	( 15'sd 10458) * $signed(input_fmap_206[7:0]) +
	( 11'sd 532) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28724) * $signed(input_fmap_208[7:0]) +
	( 16'sd 21167) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5618) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26990) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12501) * $signed(input_fmap_212[7:0]) +
	( 16'sd 22751) * $signed(input_fmap_213[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_214[7:0]) +
	( 16'sd 31034) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11521) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19551) * $signed(input_fmap_217[7:0]) +
	( 16'sd 17665) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31917) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23138) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2771) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2513) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27443) * $signed(input_fmap_224[7:0]) +
	( 15'sd 10584) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30446) * $signed(input_fmap_226[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_227[7:0]) +
	( 14'sd 7667) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10373) * $signed(input_fmap_229[7:0]) +
	( 16'sd 25847) * $signed(input_fmap_230[7:0]) +
	( 16'sd 16903) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7524) * $signed(input_fmap_232[7:0]) +
	( 16'sd 20091) * $signed(input_fmap_233[7:0]) +
	( 16'sd 30014) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21094) * $signed(input_fmap_235[7:0]) +
	( 15'sd 14006) * $signed(input_fmap_236[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16460) * $signed(input_fmap_238[7:0]) +
	( 14'sd 4170) * $signed(input_fmap_239[7:0]) +
	( 15'sd 14840) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7797) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15583) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6821) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13880) * $signed(input_fmap_244[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11955) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9816) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26167) * $signed(input_fmap_248[7:0]) +
	( 16'sd 20860) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24179) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2614) * $signed(input_fmap_251[7:0]) +
	( 11'sd 607) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31513) * $signed(input_fmap_254[7:0]) +
	( 15'sd 15083) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_118;
assign conv_mac_118 = 
	( 12'sd 1383) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10102) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22292) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13747) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27104) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5001) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8864) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13081) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14492) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18586) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6280) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1922) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29723) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3574) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7749) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15689) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31889) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27096) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20314) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22154) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23891) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5426) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16289) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20979) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18335) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26744) * $signed(input_fmap_27[7:0]) +
	( 14'sd 8022) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9242) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1535) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10957) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5279) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11150) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9009) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7852) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25216) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17678) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29419) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14153) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7556) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19352) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22601) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8769) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1223) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21782) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26089) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20508) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23705) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2274) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21270) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21415) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13526) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22698) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1834) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18054) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7436) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6654) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19025) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1298) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14832) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18212) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24587) * $signed(input_fmap_67[7:0]) +
	( 10'sd 333) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32446) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10671) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18921) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25102) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11476) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16713) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13075) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_76[7:0]) +
	( 11'sd 563) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20380) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29281) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20466) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20425) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31269) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4855) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7541) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4410) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20988) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28829) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13968) * $signed(input_fmap_90[7:0]) +
	( 11'sd 538) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19953) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11938) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_94[7:0]) +
	( 11'sd 761) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24111) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15166) * $signed(input_fmap_98[7:0]) +
	( 8'sd 115) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29401) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8567) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16251) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19840) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3927) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11864) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27227) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6519) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20901) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9807) * $signed(input_fmap_109[7:0]) +
	( 16'sd 16853) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27942) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13546) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28562) * $signed(input_fmap_113[7:0]) +
	( 13'sd 4082) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26981) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2472) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25291) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2076) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9483) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8039) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31057) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26807) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26747) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24891) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15110) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23682) * $signed(input_fmap_128[7:0]) +
	( 16'sd 32197) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18127) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20329) * $signed(input_fmap_131[7:0]) +
	( 16'sd 32341) * $signed(input_fmap_132[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31064) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31249) * $signed(input_fmap_135[7:0]) +
	( 16'sd 28828) * $signed(input_fmap_136[7:0]) +
	( 10'sd 433) * $signed(input_fmap_137[7:0]) +
	( 15'sd 12993) * $signed(input_fmap_138[7:0]) +
	( 16'sd 17422) * $signed(input_fmap_139[7:0]) +
	( 15'sd 13739) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12780) * $signed(input_fmap_141[7:0]) +
	( 16'sd 26239) * $signed(input_fmap_142[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31444) * $signed(input_fmap_144[7:0]) +
	( 16'sd 29705) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29876) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3187) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26324) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23879) * $signed(input_fmap_149[7:0]) +
	( 15'sd 8704) * $signed(input_fmap_150[7:0]) +
	( 16'sd 20394) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2863) * $signed(input_fmap_152[7:0]) +
	( 14'sd 6297) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30931) * $signed(input_fmap_154[7:0]) +
	( 16'sd 18236) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10022) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25741) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17112) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12806) * $signed(input_fmap_159[7:0]) +
	( 12'sd 1734) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1839) * $signed(input_fmap_161[7:0]) +
	( 15'sd 9159) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8830) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19586) * $signed(input_fmap_164[7:0]) +
	( 14'sd 8054) * $signed(input_fmap_165[7:0]) +
	( 15'sd 16155) * $signed(input_fmap_166[7:0]) +
	( 16'sd 32340) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20677) * $signed(input_fmap_168[7:0]) +
	( 16'sd 28211) * $signed(input_fmap_169[7:0]) +
	( 16'sd 26437) * $signed(input_fmap_170[7:0]) +
	( 16'sd 29767) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19999) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1591) * $signed(input_fmap_173[7:0]) +
	( 16'sd 22315) * $signed(input_fmap_174[7:0]) +
	( 15'sd 16293) * $signed(input_fmap_175[7:0]) +
	( 14'sd 4441) * $signed(input_fmap_176[7:0]) +
	( 13'sd 3162) * $signed(input_fmap_177[7:0]) +
	( 16'sd 25633) * $signed(input_fmap_178[7:0]) +
	( 14'sd 7079) * $signed(input_fmap_179[7:0]) +
	( 16'sd 19363) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30336) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29322) * $signed(input_fmap_182[7:0]) +
	( 15'sd 10875) * $signed(input_fmap_183[7:0]) +
	( 16'sd 27795) * $signed(input_fmap_184[7:0]) +
	( 16'sd 28286) * $signed(input_fmap_185[7:0]) +
	( 16'sd 20297) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27785) * $signed(input_fmap_187[7:0]) +
	( 15'sd 15207) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30069) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_190[7:0]) +
	( 15'sd 15400) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15552) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3363) * $signed(input_fmap_194[7:0]) +
	( 16'sd 23901) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25786) * $signed(input_fmap_196[7:0]) +
	( 16'sd 20573) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29533) * $signed(input_fmap_198[7:0]) +
	( 13'sd 4019) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25793) * $signed(input_fmap_200[7:0]) +
	( 16'sd 26046) * $signed(input_fmap_201[7:0]) +
	( 15'sd 13642) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25312) * $signed(input_fmap_203[7:0]) +
	( 16'sd 28232) * $signed(input_fmap_204[7:0]) +
	( 15'sd 14180) * $signed(input_fmap_205[7:0]) +
	( 16'sd 25830) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21410) * $signed(input_fmap_207[7:0]) +
	( 13'sd 3620) * $signed(input_fmap_208[7:0]) +
	( 10'sd 356) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15411) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26370) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_212[7:0]) +
	( 14'sd 4616) * $signed(input_fmap_213[7:0]) +
	( 15'sd 11690) * $signed(input_fmap_214[7:0]) +
	( 16'sd 24011) * $signed(input_fmap_215[7:0]) +
	( 14'sd 6165) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24765) * $signed(input_fmap_217[7:0]) +
	( 12'sd 1278) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19793) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15901) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10551) * $signed(input_fmap_222[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_223[7:0]) +
	( 13'sd 2392) * $signed(input_fmap_224[7:0]) +
	( 14'sd 4786) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27353) * $signed(input_fmap_226[7:0]) +
	( 16'sd 17367) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4879) * $signed(input_fmap_228[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28730) * $signed(input_fmap_230[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_231[7:0]) +
	( 16'sd 23355) * $signed(input_fmap_232[7:0]) +
	( 16'sd 30956) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13435) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5035) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2941) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_237[7:0]) +
	( 16'sd 20510) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20040) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10254) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29154) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13447) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13670) * $signed(input_fmap_244[7:0]) +
	( 16'sd 26015) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15042) * $signed(input_fmap_246[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13019) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14509) * $signed(input_fmap_249[7:0]) +
	( 12'sd 1447) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2761) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27527) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3896) * $signed(input_fmap_253[7:0]) +
	( 14'sd 6683) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11475) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_119;
assign conv_mac_119 = 
	( 14'sd 4375) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2133) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30218) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26719) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31951) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23264) * $signed(input_fmap_6[7:0]) +
	( 9'sd 198) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24196) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15817) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17191) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29721) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6893) * $signed(input_fmap_13[7:0]) +
	( 6'sd 27) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1371) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23189) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2769) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11751) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10180) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22133) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11912) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17487) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25834) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19514) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16895) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31142) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2056) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9979) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26639) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12841) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21587) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4527) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11360) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31832) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18273) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18081) * $signed(input_fmap_36[7:0]) +
	( 11'sd 624) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28926) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4228) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28704) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31199) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8440) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8310) * $signed(input_fmap_43[7:0]) +
	( 13'sd 4073) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19508) * $signed(input_fmap_47[7:0]) +
	( 6'sd 25) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24992) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6053) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18779) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17833) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30289) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19398) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20626) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26144) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16330) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16596) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16241) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32339) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8364) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7469) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28976) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29861) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26255) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25442) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7762) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15513) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21729) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25299) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17126) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29125) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4596) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25147) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16706) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27772) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2641) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7814) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27997) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20652) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2631) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18704) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15359) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9028) * $signed(input_fmap_85[7:0]) +
	( 13'sd 4011) * $signed(input_fmap_86[7:0]) +
	( 11'sd 1009) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20675) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5811) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17134) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15667) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18845) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7573) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25457) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10669) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31232) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14815) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22393) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29618) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5433) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7919) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12749) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28450) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1974) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5763) * $signed(input_fmap_110[7:0]) +
	( 11'sd 1008) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30628) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22762) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24364) * $signed(input_fmap_115[7:0]) +
	( 10'sd 298) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27145) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2689) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20822) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30413) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1626) * $signed(input_fmap_121[7:0]) +
	( 15'sd 11488) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25253) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21523) * $signed(input_fmap_124[7:0]) +
	( 14'sd 8004) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18367) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6687) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31302) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28816) * $signed(input_fmap_129[7:0]) +
	( 15'sd 16306) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10043) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32293) * $signed(input_fmap_134[7:0]) +
	( 15'sd 8615) * $signed(input_fmap_135[7:0]) +
	( 15'sd 11872) * $signed(input_fmap_136[7:0]) +
	( 16'sd 23796) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31211) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31966) * $signed(input_fmap_139[7:0]) +
	( 16'sd 21358) * $signed(input_fmap_140[7:0]) +
	( 16'sd 30417) * $signed(input_fmap_141[7:0]) +
	( 15'sd 16028) * $signed(input_fmap_142[7:0]) +
	( 15'sd 15198) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3867) * $signed(input_fmap_144[7:0]) +
	( 15'sd 11308) * $signed(input_fmap_145[7:0]) +
	( 15'sd 8259) * $signed(input_fmap_146[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22273) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17089) * $signed(input_fmap_149[7:0]) +
	( 16'sd 28691) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12471) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22778) * $signed(input_fmap_152[7:0]) +
	( 16'sd 20867) * $signed(input_fmap_153[7:0]) +
	( 15'sd 8484) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23155) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29281) * $signed(input_fmap_156[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17889) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21802) * $signed(input_fmap_159[7:0]) +
	( 16'sd 23486) * $signed(input_fmap_160[7:0]) +
	( 16'sd 29072) * $signed(input_fmap_161[7:0]) +
	( 16'sd 23407) * $signed(input_fmap_162[7:0]) +
	( 15'sd 13796) * $signed(input_fmap_163[7:0]) +
	( 16'sd 21691) * $signed(input_fmap_164[7:0]) +
	( 14'sd 5184) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9042) * $signed(input_fmap_166[7:0]) +
	( 13'sd 3046) * $signed(input_fmap_167[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26127) * $signed(input_fmap_169[7:0]) +
	( 16'sd 26553) * $signed(input_fmap_170[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12761) * $signed(input_fmap_172[7:0]) +
	( 16'sd 22708) * $signed(input_fmap_173[7:0]) +
	( 13'sd 2947) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15125) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10132) * $signed(input_fmap_176[7:0]) +
	( 13'sd 3929) * $signed(input_fmap_177[7:0]) +
	( 16'sd 20981) * $signed(input_fmap_178[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_179[7:0]) +
	( 16'sd 30219) * $signed(input_fmap_180[7:0]) +
	( 16'sd 22318) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5056) * $signed(input_fmap_182[7:0]) +
	( 16'sd 20873) * $signed(input_fmap_183[7:0]) +
	( 16'sd 21812) * $signed(input_fmap_184[7:0]) +
	( 15'sd 10868) * $signed(input_fmap_185[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_186[7:0]) +
	( 16'sd 16730) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13890) * $signed(input_fmap_188[7:0]) +
	( 16'sd 27881) * $signed(input_fmap_189[7:0]) +
	( 16'sd 25496) * $signed(input_fmap_190[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_191[7:0]) +
	( 16'sd 21880) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22525) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18653) * $signed(input_fmap_194[7:0]) +
	( 13'sd 4050) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6128) * $signed(input_fmap_196[7:0]) +
	( 16'sd 23267) * $signed(input_fmap_197[7:0]) +
	( 11'sd 836) * $signed(input_fmap_198[7:0]) +
	( 15'sd 9826) * $signed(input_fmap_199[7:0]) +
	( 12'sd 1040) * $signed(input_fmap_200[7:0]) +
	( 15'sd 14060) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17128) * $signed(input_fmap_202[7:0]) +
	( 15'sd 11845) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6375) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30354) * $signed(input_fmap_205[7:0]) +
	( 16'sd 23968) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12522) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4892) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22528) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4984) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14054) * $signed(input_fmap_212[7:0]) +
	( 16'sd 32708) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17978) * $signed(input_fmap_214[7:0]) +
	( 15'sd 15387) * $signed(input_fmap_215[7:0]) +
	( 15'sd 9824) * $signed(input_fmap_216[7:0]) +
	( 16'sd 20488) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21569) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21646) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26568) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27832) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12662) * $signed(input_fmap_222[7:0]) +
	( 16'sd 27392) * $signed(input_fmap_223[7:0]) +
	( 16'sd 23936) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27651) * $signed(input_fmap_225[7:0]) +
	( 14'sd 4241) * $signed(input_fmap_226[7:0]) +
	( 16'sd 18448) * $signed(input_fmap_227[7:0]) +
	( 15'sd 14627) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3152) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27923) * $signed(input_fmap_230[7:0]) +
	( 16'sd 21605) * $signed(input_fmap_231[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_232[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5371) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5865) * $signed(input_fmap_235[7:0]) +
	( 16'sd 32615) * $signed(input_fmap_236[7:0]) +
	( 14'sd 5212) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17075) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13112) * $signed(input_fmap_239[7:0]) +
	( 15'sd 15514) * $signed(input_fmap_240[7:0]) +
	( 15'sd 10687) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17649) * $signed(input_fmap_242[7:0]) +
	( 16'sd 16567) * $signed(input_fmap_243[7:0]) +
	( 14'sd 4881) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24057) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20012) * $signed(input_fmap_246[7:0]) +
	( 14'sd 7442) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32310) * $signed(input_fmap_248[7:0]) +
	( 16'sd 18003) * $signed(input_fmap_249[7:0]) +
	( 16'sd 31842) * $signed(input_fmap_250[7:0]) +
	( 15'sd 16242) * $signed(input_fmap_251[7:0]) +
	( 15'sd 11656) * $signed(input_fmap_252[7:0]) +
	( 16'sd 20099) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5036) * $signed(input_fmap_254[7:0]) +
	( 15'sd 13501) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_120;
assign conv_mac_120 = 
	( 15'sd 10077) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1444) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1575) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28568) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11638) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12523) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24760) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10290) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27074) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16771) * $signed(input_fmap_10[7:0]) +
	( 13'sd 3482) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29584) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25773) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17038) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5428) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14306) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22911) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10764) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13042) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32309) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23866) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4367) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28152) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24107) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1905) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30913) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31310) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23223) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32585) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11073) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30095) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22655) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11149) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21493) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9557) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30158) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28410) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24006) * $signed(input_fmap_41[7:0]) +
	( 9'sd 246) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26766) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2648) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16094) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6997) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27202) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29068) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6731) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22354) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8296) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11809) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15227) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3165) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3771) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7895) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12923) * $signed(input_fmap_58[7:0]) +
	( 11'sd 739) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10906) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14986) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22110) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23810) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7508) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21973) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12793) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15352) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7137) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28537) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5090) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2288) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26466) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21633) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11807) * $signed(input_fmap_79[7:0]) +
	( 10'sd 463) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27864) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16941) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12823) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28106) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16970) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15431) * $signed(input_fmap_87[7:0]) +
	( 12'sd 2022) * $signed(input_fmap_88[7:0]) +
	( 9'sd 194) * $signed(input_fmap_89[7:0]) +
	( 14'sd 8096) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20557) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14987) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29380) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21752) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16155) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7108) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16984) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21061) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11671) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3891) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22616) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25806) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21321) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18011) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24627) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12941) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29669) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10353) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18389) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24309) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8878) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21624) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17708) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11129) * $signed(input_fmap_118[7:0]) +
	( 14'sd 8190) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31558) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1849) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19296) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29918) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21739) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29265) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24576) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17592) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29551) * $signed(input_fmap_128[7:0]) +
	( 14'sd 4679) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6059) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_131[7:0]) +
	( 16'sd 19767) * $signed(input_fmap_132[7:0]) +
	( 14'sd 6040) * $signed(input_fmap_133[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_134[7:0]) +
	( 16'sd 17564) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_136[7:0]) +
	( 15'sd 10049) * $signed(input_fmap_137[7:0]) +
	( 13'sd 2631) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_139[7:0]) +
	( 15'sd 14625) * $signed(input_fmap_140[7:0]) +
	( 16'sd 30179) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8929) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20743) * $signed(input_fmap_143[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_144[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21388) * $signed(input_fmap_147[7:0]) +
	( 16'sd 18518) * $signed(input_fmap_148[7:0]) +
	( 16'sd 31846) * $signed(input_fmap_149[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17248) * $signed(input_fmap_151[7:0]) +
	( 15'sd 11427) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_153[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_154[7:0]) +
	( 15'sd 14396) * $signed(input_fmap_155[7:0]) +
	( 16'sd 16866) * $signed(input_fmap_156[7:0]) +
	( 13'sd 3779) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18313) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2687) * $signed(input_fmap_159[7:0]) +
	( 16'sd 20684) * $signed(input_fmap_160[7:0]) +
	( 15'sd 13391) * $signed(input_fmap_161[7:0]) +
	( 14'sd 8025) * $signed(input_fmap_162[7:0]) +
	( 14'sd 7204) * $signed(input_fmap_163[7:0]) +
	( 14'sd 5991) * $signed(input_fmap_164[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_165[7:0]) +
	( 15'sd 12452) * $signed(input_fmap_166[7:0]) +
	( 15'sd 15577) * $signed(input_fmap_167[7:0]) +
	( 16'sd 31747) * $signed(input_fmap_168[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17246) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31896) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22205) * $signed(input_fmap_172[7:0]) +
	( 15'sd 15887) * $signed(input_fmap_173[7:0]) +
	( 10'sd 381) * $signed(input_fmap_174[7:0]) +
	( 16'sd 18059) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1879) * $signed(input_fmap_177[7:0]) +
	( 13'sd 3892) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22507) * $signed(input_fmap_179[7:0]) +
	( 16'sd 22665) * $signed(input_fmap_180[7:0]) +
	( 16'sd 29695) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4708) * $signed(input_fmap_182[7:0]) +
	( 14'sd 7697) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30710) * $signed(input_fmap_184[7:0]) +
	( 16'sd 31875) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26590) * $signed(input_fmap_186[7:0]) +
	( 16'sd 24042) * $signed(input_fmap_187[7:0]) +
	( 15'sd 8885) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30133) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30319) * $signed(input_fmap_190[7:0]) +
	( 15'sd 12048) * $signed(input_fmap_191[7:0]) +
	( 10'sd 370) * $signed(input_fmap_192[7:0]) +
	( 12'sd 1065) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26230) * $signed(input_fmap_194[7:0]) +
	( 15'sd 10416) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6925) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_197[7:0]) +
	( 16'sd 25139) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6500) * $signed(input_fmap_199[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13623) * $signed(input_fmap_201[7:0]) +
	( 15'sd 16219) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30609) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11963) * $signed(input_fmap_204[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27107) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7705) * $signed(input_fmap_207[7:0]) +
	( 14'sd 7363) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24112) * $signed(input_fmap_209[7:0]) +
	( 16'sd 32117) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5866) * $signed(input_fmap_211[7:0]) +
	( 16'sd 30993) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9759) * $signed(input_fmap_213[7:0]) +
	( 16'sd 21535) * $signed(input_fmap_214[7:0]) +
	( 15'sd 8420) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24006) * $signed(input_fmap_216[7:0]) +
	( 11'sd 788) * $signed(input_fmap_217[7:0]) +
	( 14'sd 6593) * $signed(input_fmap_218[7:0]) +
	( 14'sd 4836) * $signed(input_fmap_219[7:0]) +
	( 15'sd 15018) * $signed(input_fmap_220[7:0]) +
	( 16'sd 32514) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_222[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_223[7:0]) +
	( 16'sd 28119) * $signed(input_fmap_224[7:0]) +
	( 15'sd 10160) * $signed(input_fmap_225[7:0]) +
	( 14'sd 5821) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26422) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23395) * $signed(input_fmap_229[7:0]) +
	( 16'sd 17475) * $signed(input_fmap_230[7:0]) +
	( 15'sd 9776) * $signed(input_fmap_231[7:0]) +
	( 16'sd 32571) * $signed(input_fmap_232[7:0]) +
	( 10'sd 380) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4414) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19697) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11135) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6646) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14097) * $signed(input_fmap_238[7:0]) +
	( 15'sd 8500) * $signed(input_fmap_239[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_240[7:0]) +
	( 15'sd 13656) * $signed(input_fmap_241[7:0]) +
	( 16'sd 31858) * $signed(input_fmap_242[7:0]) +
	( 12'sd 1055) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13543) * $signed(input_fmap_244[7:0]) +
	( 15'sd 13130) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28426) * $signed(input_fmap_246[7:0]) +
	( 16'sd 26337) * $signed(input_fmap_247[7:0]) +
	( 15'sd 15650) * $signed(input_fmap_248[7:0]) +
	( 15'sd 10545) * $signed(input_fmap_249[7:0]) +
	( 15'sd 11553) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21559) * $signed(input_fmap_251[7:0]) +
	( 16'sd 29199) * $signed(input_fmap_252[7:0]) +
	( 16'sd 19409) * $signed(input_fmap_253[7:0]) +
	( 14'sd 8147) * $signed(input_fmap_254[7:0]) +
	( 16'sd 17001) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_121;
assign conv_mac_121 = 
	( 13'sd 2826) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21974) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23059) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16068) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23146) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30943) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1650) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10065) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11446) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21332) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10820) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29069) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28587) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1812) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31310) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4617) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32013) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25399) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21463) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2824) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14936) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32736) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27489) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14546) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8945) * $signed(input_fmap_27[7:0]) +
	( 16'sd 29928) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9245) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21913) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19134) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29840) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14304) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5395) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1672) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31762) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23309) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28711) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2325) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18164) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24353) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_44[7:0]) +
	( 15'sd 8349) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12771) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24086) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31563) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9170) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16139) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25592) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15079) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7268) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24580) * $signed(input_fmap_54[7:0]) +
	( 13'sd 2664) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10807) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2790) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6121) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8226) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1819) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28637) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16331) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4909) * $signed(input_fmap_64[7:0]) +
	( 15'sd 14833) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18631) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27456) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31873) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6951) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9516) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15707) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7023) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26719) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22030) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8922) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32586) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28362) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10853) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29505) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24210) * $signed(input_fmap_81[7:0]) +
	( 16'sd 17081) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31835) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21534) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6510) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1780) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23357) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9851) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14458) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2576) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31343) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5872) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16277) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16677) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22446) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29990) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29726) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12164) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22454) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10640) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21513) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1670) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32451) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3673) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14967) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12219) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23472) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24039) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22267) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4214) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16021) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10019) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30855) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14760) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25669) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14727) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11598) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5728) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23822) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4170) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24738) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28268) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15032) * $signed(input_fmap_127[7:0]) +
	( 12'sd 1769) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14415) * $signed(input_fmap_129[7:0]) +
	( 15'sd 13889) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5903) * $signed(input_fmap_132[7:0]) +
	( 14'sd 7142) * $signed(input_fmap_133[7:0]) +
	( 15'sd 14284) * $signed(input_fmap_134[7:0]) +
	( 13'sd 2268) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23452) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9840) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11067) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9224) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3343) * $signed(input_fmap_141[7:0]) +
	( 11'sd 872) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12371) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31044) * $signed(input_fmap_144[7:0]) +
	( 13'sd 3526) * $signed(input_fmap_145[7:0]) +
	( 15'sd 11484) * $signed(input_fmap_146[7:0]) +
	( 15'sd 10407) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11415) * $signed(input_fmap_148[7:0]) +
	( 16'sd 32618) * $signed(input_fmap_149[7:0]) +
	( 15'sd 16337) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12786) * $signed(input_fmap_151[7:0]) +
	( 15'sd 12937) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27394) * $signed(input_fmap_153[7:0]) +
	( 15'sd 12035) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28790) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10112) * $signed(input_fmap_156[7:0]) +
	( 15'sd 12579) * $signed(input_fmap_157[7:0]) +
	( 16'sd 27030) * $signed(input_fmap_158[7:0]) +
	( 16'sd 28566) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26448) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2376) * $signed(input_fmap_162[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19951) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23394) * $signed(input_fmap_165[7:0]) +
	( 15'sd 11847) * $signed(input_fmap_166[7:0]) +
	( 15'sd 11024) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17482) * $signed(input_fmap_168[7:0]) +
	( 15'sd 8944) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14697) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12030) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31346) * $signed(input_fmap_172[7:0]) +
	( 14'sd 7589) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14220) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17615) * $signed(input_fmap_175[7:0]) +
	( 16'sd 24899) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6412) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1575) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25620) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24779) * $signed(input_fmap_180[7:0]) +
	( 15'sd 8391) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10842) * $signed(input_fmap_182[7:0]) +
	( 15'sd 15369) * $signed(input_fmap_183[7:0]) +
	( 16'sd 21885) * $signed(input_fmap_184[7:0]) +
	( 15'sd 12161) * $signed(input_fmap_185[7:0]) +
	( 16'sd 22651) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4898) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32046) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19234) * $signed(input_fmap_189[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_190[7:0]) +
	( 15'sd 10575) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31376) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20704) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30826) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_195[7:0]) +
	( 16'sd 30117) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21673) * $signed(input_fmap_197[7:0]) +
	( 15'sd 8711) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10363) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13466) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18229) * $signed(input_fmap_201[7:0]) +
	( 16'sd 26803) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25718) * $signed(input_fmap_203[7:0]) +
	( 16'sd 22206) * $signed(input_fmap_204[7:0]) +
	( 15'sd 14475) * $signed(input_fmap_205[7:0]) +
	( 16'sd 26074) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7830) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18937) * $signed(input_fmap_208[7:0]) +
	( 11'sd 561) * $signed(input_fmap_209[7:0]) +
	( 14'sd 6832) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23609) * $signed(input_fmap_211[7:0]) +
	( 16'sd 21913) * $signed(input_fmap_212[7:0]) +
	( 8'sd 100) * $signed(input_fmap_213[7:0]) +
	( 14'sd 6211) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29152) * $signed(input_fmap_215[7:0]) +
	( 16'sd 27803) * $signed(input_fmap_216[7:0]) +
	( 14'sd 7733) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7081) * $signed(input_fmap_218[7:0]) +
	( 15'sd 16106) * $signed(input_fmap_219[7:0]) +
	( 14'sd 5100) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5377) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28649) * $signed(input_fmap_222[7:0]) +
	( 16'sd 27243) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30228) * $signed(input_fmap_224[7:0]) +
	( 16'sd 25047) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14205) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5753) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4593) * $signed(input_fmap_228[7:0]) +
	( 14'sd 7763) * $signed(input_fmap_229[7:0]) +
	( 15'sd 11769) * $signed(input_fmap_230[7:0]) +
	( 16'sd 27976) * $signed(input_fmap_231[7:0]) +
	( 14'sd 4127) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1318) * $signed(input_fmap_233[7:0]) +
	( 16'sd 29356) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19023) * $signed(input_fmap_235[7:0]) +
	( 16'sd 29950) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6988) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_238[7:0]) +
	( 15'sd 11763) * $signed(input_fmap_239[7:0]) +
	( 16'sd 27303) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23511) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28892) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13512) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10703) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22666) * $signed(input_fmap_246[7:0]) +
	( 16'sd 25344) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4247) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14087) * $signed(input_fmap_249[7:0]) +
	( 13'sd 4011) * $signed(input_fmap_250[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_251[7:0]) +
	( 16'sd 22143) * $signed(input_fmap_252[7:0]) +
	( 14'sd 7605) * $signed(input_fmap_253[7:0]) +
	( 15'sd 15042) * $signed(input_fmap_254[7:0]) +
	( 16'sd 29386) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_122;
assign conv_mac_122 = 
	( 9'sd 182) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24698) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29626) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11332) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6731) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21519) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19128) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19676) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2846) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22176) * $signed(input_fmap_11[7:0]) +
	( 11'sd 645) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10155) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14940) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14537) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29793) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3853) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3199) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9859) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5738) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24426) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6229) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22742) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26513) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10261) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10975) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14616) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19628) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17313) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27478) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20258) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6786) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20766) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20396) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31743) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10049) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29532) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9413) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28169) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18596) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3066) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30252) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10653) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22754) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26371) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29699) * $signed(input_fmap_49[7:0]) +
	( 8'sd 68) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3872) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3366) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8219) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4440) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20169) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21670) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21981) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26551) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5018) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16458) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24620) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9055) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17736) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8757) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16939) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14163) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8620) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17593) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11450) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13523) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7803) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18974) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8621) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12301) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18293) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4905) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5230) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27889) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11432) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6374) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10812) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24281) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3893) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9909) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2062) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16570) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30060) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14042) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3787) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19525) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26295) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32725) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7724) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21390) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25179) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32541) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28246) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5828) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2222) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4235) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25034) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25005) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13338) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29266) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28797) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32647) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24235) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31241) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28309) * $signed(input_fmap_116[7:0]) +
	( 10'sd 443) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15144) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26580) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29547) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14966) * $signed(input_fmap_121[7:0]) +
	( 8'sd 82) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11200) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9076) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27781) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23211) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25075) * $signed(input_fmap_127[7:0]) +
	( 14'sd 7327) * $signed(input_fmap_128[7:0]) +
	( 16'sd 30460) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12337) * $signed(input_fmap_130[7:0]) +
	( 15'sd 12567) * $signed(input_fmap_131[7:0]) +
	( 16'sd 22212) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11344) * $signed(input_fmap_133[7:0]) +
	( 16'sd 23589) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19979) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31045) * $signed(input_fmap_136[7:0]) +
	( 9'sd 169) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22385) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20317) * $signed(input_fmap_139[7:0]) +
	( 16'sd 27357) * $signed(input_fmap_140[7:0]) +
	( 12'sd 1079) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19776) * $signed(input_fmap_142[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22965) * $signed(input_fmap_144[7:0]) +
	( 10'sd 479) * $signed(input_fmap_145[7:0]) +
	( 14'sd 5189) * $signed(input_fmap_146[7:0]) +
	( 15'sd 10162) * $signed(input_fmap_147[7:0]) +
	( 16'sd 24086) * $signed(input_fmap_148[7:0]) +
	( 16'sd 32038) * $signed(input_fmap_149[7:0]) +
	( 14'sd 4908) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19876) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14805) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24196) * $signed(input_fmap_153[7:0]) +
	( 13'sd 2253) * $signed(input_fmap_154[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17834) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24873) * $signed(input_fmap_157[7:0]) +
	( 15'sd 14423) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14767) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_160[7:0]) +
	( 15'sd 8525) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10330) * $signed(input_fmap_162[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13145) * $signed(input_fmap_164[7:0]) +
	( 16'sd 29361) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13914) * $signed(input_fmap_166[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29094) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21779) * $signed(input_fmap_169[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_170[7:0]) +
	( 15'sd 14682) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3161) * $signed(input_fmap_172[7:0]) +
	( 16'sd 16590) * $signed(input_fmap_173[7:0]) +
	( 15'sd 9527) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4104) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3315) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15081) * $signed(input_fmap_177[7:0]) +
	( 16'sd 23779) * $signed(input_fmap_178[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24874) * $signed(input_fmap_180[7:0]) +
	( 14'sd 7426) * $signed(input_fmap_181[7:0]) +
	( 16'sd 22432) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29491) * $signed(input_fmap_183[7:0]) +
	( 14'sd 7483) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_186[7:0]) +
	( 12'sd 2014) * $signed(input_fmap_187[7:0]) +
	( 16'sd 19871) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2964) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13901) * $signed(input_fmap_190[7:0]) +
	( 16'sd 30220) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26272) * $signed(input_fmap_193[7:0]) +
	( 15'sd 16350) * $signed(input_fmap_194[7:0]) +
	( 16'sd 20574) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6436) * $signed(input_fmap_196[7:0]) +
	( 16'sd 30845) * $signed(input_fmap_197[7:0]) +
	( 13'sd 3164) * $signed(input_fmap_198[7:0]) +
	( 14'sd 7359) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29245) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11266) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8656) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19069) * $signed(input_fmap_203[7:0]) +
	( 13'sd 3735) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29884) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21958) * $signed(input_fmap_206[7:0]) +
	( 16'sd 24652) * $signed(input_fmap_207[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19959) * $signed(input_fmap_209[7:0]) +
	( 16'sd 29140) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12767) * $signed(input_fmap_211[7:0]) +
	( 15'sd 8530) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2934) * $signed(input_fmap_213[7:0]) +
	( 16'sd 22556) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22238) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19885) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10108) * $signed(input_fmap_217[7:0]) +
	( 13'sd 3388) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12637) * $signed(input_fmap_219[7:0]) +
	( 16'sd 32581) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_221[7:0]) +
	( 12'sd 1116) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22996) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25962) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5553) * $signed(input_fmap_225[7:0]) +
	( 15'sd 16245) * $signed(input_fmap_226[7:0]) +
	( 15'sd 10037) * $signed(input_fmap_227[7:0]) +
	( 15'sd 16003) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29481) * $signed(input_fmap_229[7:0]) +
	( 16'sd 31549) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25178) * $signed(input_fmap_231[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18949) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_234[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2350) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28514) * $signed(input_fmap_238[7:0]) +
	( 16'sd 24698) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9059) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23396) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17888) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7484) * $signed(input_fmap_243[7:0]) +
	( 15'sd 10519) * $signed(input_fmap_244[7:0]) +
	( 15'sd 16094) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28604) * $signed(input_fmap_246[7:0]) +
	( 16'sd 25017) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13999) * $signed(input_fmap_248[7:0]) +
	( 16'sd 29775) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12607) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27486) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28696) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2816) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1277) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20840) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_123;
assign conv_mac_123 = 
	( 15'sd 13337) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28597) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6288) * $signed(input_fmap_2[7:0]) +
	( 14'sd 8149) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24448) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6309) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22953) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29418) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17512) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29149) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32512) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9101) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26050) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30966) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21097) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27041) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28802) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14666) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31238) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2821) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20596) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32160) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27172) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19592) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10432) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31735) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8281) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16432) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6683) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19593) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6632) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18477) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16190) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23850) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3715) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13726) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17935) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27824) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12837) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17191) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21820) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10571) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22590) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19038) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10950) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4447) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19413) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10369) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11599) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3353) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11788) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6535) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8300) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13347) * $signed(input_fmap_55[7:0]) +
	( 11'sd 921) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15156) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22515) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19889) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29333) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30906) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15253) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5614) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16416) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19124) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7144) * $signed(input_fmap_67[7:0]) +
	( 10'sd 292) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11290) * $signed(input_fmap_69[7:0]) +
	( 16'sd 31512) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20395) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29152) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21099) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19149) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6271) * $signed(input_fmap_76[7:0]) +
	( 13'sd 4022) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23496) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12877) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30563) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32219) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21135) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5540) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18328) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30796) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31603) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32496) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8788) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29569) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5916) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31958) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1691) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15492) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21072) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13810) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11598) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9758) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10413) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15951) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30469) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24797) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29700) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28410) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14958) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18835) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2592) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25775) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6678) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22969) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9812) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10174) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13738) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18211) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29357) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12784) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_123[7:0]) +
	( 10'sd 316) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22557) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_126[7:0]) +
	( 11'sd 817) * $signed(input_fmap_127[7:0]) +
	( 14'sd 5524) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27939) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_130[7:0]) +
	( 14'sd 7149) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14435) * $signed(input_fmap_132[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21341) * $signed(input_fmap_134[7:0]) +
	( 14'sd 6839) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13687) * $signed(input_fmap_136[7:0]) +
	( 10'sd 447) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22078) * $signed(input_fmap_138[7:0]) +
	( 12'sd 1856) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24035) * $signed(input_fmap_140[7:0]) +
	( 16'sd 32305) * $signed(input_fmap_141[7:0]) +
	( 14'sd 7940) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31104) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_144[7:0]) +
	( 15'sd 11311) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_146[7:0]) +
	( 10'sd 487) * $signed(input_fmap_147[7:0]) +
	( 15'sd 12757) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18192) * $signed(input_fmap_151[7:0]) +
	( 16'sd 17133) * $signed(input_fmap_152[7:0]) +
	( 16'sd 22079) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25279) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27884) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20220) * $signed(input_fmap_156[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_157[7:0]) +
	( 16'sd 21016) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14057) * $signed(input_fmap_159[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_160[7:0]) +
	( 16'sd 27176) * $signed(input_fmap_161[7:0]) +
	( 13'sd 3289) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22125) * $signed(input_fmap_163[7:0]) +
	( 16'sd 18402) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28444) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3488) * $signed(input_fmap_166[7:0]) +
	( 15'sd 11800) * $signed(input_fmap_167[7:0]) +
	( 16'sd 16842) * $signed(input_fmap_168[7:0]) +
	( 16'sd 19483) * $signed(input_fmap_169[7:0]) +
	( 13'sd 3903) * $signed(input_fmap_170[7:0]) +
	( 16'sd 21309) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15149) * $signed(input_fmap_172[7:0]) +
	( 16'sd 28115) * $signed(input_fmap_173[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1214) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22914) * $signed(input_fmap_177[7:0]) +
	( 16'sd 25553) * $signed(input_fmap_178[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6949) * $signed(input_fmap_180[7:0]) +
	( 16'sd 27665) * $signed(input_fmap_181[7:0]) +
	( 16'sd 22011) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2530) * $signed(input_fmap_183[7:0]) +
	( 12'sd 1763) * $signed(input_fmap_184[7:0]) +
	( 15'sd 14435) * $signed(input_fmap_185[7:0]) +
	( 15'sd 14669) * $signed(input_fmap_186[7:0]) +
	( 16'sd 16645) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31556) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3173) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28639) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3782) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24574) * $signed(input_fmap_192[7:0]) +
	( 15'sd 13484) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27928) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14377) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12368) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19238) * $signed(input_fmap_197[7:0]) +
	( 16'sd 28600) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14079) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31599) * $signed(input_fmap_200[7:0]) +
	( 16'sd 32457) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31077) * $signed(input_fmap_202[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_203[7:0]) +
	( 13'sd 3395) * $signed(input_fmap_204[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6637) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3841) * $signed(input_fmap_207[7:0]) +
	( 16'sd 20397) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14285) * $signed(input_fmap_209[7:0]) +
	( 15'sd 16056) * $signed(input_fmap_210[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1573) * $signed(input_fmap_212[7:0]) +
	( 16'sd 26196) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14349) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23022) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20654) * $signed(input_fmap_216[7:0]) +
	( 16'sd 29842) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10219) * $signed(input_fmap_218[7:0]) +
	( 11'sd 788) * $signed(input_fmap_219[7:0]) +
	( 15'sd 9264) * $signed(input_fmap_220[7:0]) +
	( 15'sd 14732) * $signed(input_fmap_221[7:0]) +
	( 16'sd 24109) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9981) * $signed(input_fmap_223[7:0]) +
	( 16'sd 27234) * $signed(input_fmap_224[7:0]) +
	( 16'sd 28303) * $signed(input_fmap_225[7:0]) +
	( 13'sd 2080) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27545) * $signed(input_fmap_227[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20378) * $signed(input_fmap_229[7:0]) +
	( 16'sd 25753) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10417) * $signed(input_fmap_231[7:0]) +
	( 16'sd 17152) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5511) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3782) * $signed(input_fmap_234[7:0]) +
	( 12'sd 1563) * $signed(input_fmap_235[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_236[7:0]) +
	( 14'sd 7935) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27375) * $signed(input_fmap_238[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31657) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7024) * $signed(input_fmap_241[7:0]) +
	( 15'sd 10601) * $signed(input_fmap_242[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28664) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22527) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10994) * $signed(input_fmap_246[7:0]) +
	( 16'sd 16391) * $signed(input_fmap_247[7:0]) +
	( 16'sd 19481) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21774) * $signed(input_fmap_249[7:0]) +
	( 15'sd 13136) * $signed(input_fmap_250[7:0]) +
	( 16'sd 31980) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6029) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2979) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20579) * $signed(input_fmap_254[7:0]) +
	( 14'sd 7024) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_124;
assign conv_mac_124 = 
	( 16'sd 18031) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9160) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1614) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7820) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12742) * $signed(input_fmap_4[7:0]) +
	( 10'sd 334) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22790) * $signed(input_fmap_6[7:0]) +
	( 8'sd 127) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27642) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29902) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1412) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11936) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16328) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11044) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11235) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7489) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28418) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5745) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18450) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30333) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1968) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17205) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1750) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12407) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2081) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15651) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27270) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12775) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17810) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28498) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9715) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28301) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9685) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26934) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29429) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28882) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29157) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9110) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18264) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30771) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24178) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31141) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2339) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17848) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31290) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31058) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15097) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19172) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4688) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4895) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16139) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10379) * $signed(input_fmap_58[7:0]) +
	( 14'sd 5286) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31577) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28498) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20710) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12096) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24465) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25282) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24064) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31272) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31723) * $signed(input_fmap_68[7:0]) +
	( 8'sd 77) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1556) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11428) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32107) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21417) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7508) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14249) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29209) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10895) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3037) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7144) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8304) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8438) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3147) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21044) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32094) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5095) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25340) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6516) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29470) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10284) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15269) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3972) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30186) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5777) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23186) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25561) * $signed(input_fmap_95[7:0]) +
	( 11'sd 569) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17062) * $signed(input_fmap_97[7:0]) +
	( 11'sd 533) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32330) * $signed(input_fmap_99[7:0]) +
	( 14'sd 8080) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18528) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23477) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31863) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16425) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12589) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7573) * $signed(input_fmap_107[7:0]) +
	( 9'sd 178) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15453) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21163) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2166) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8865) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10663) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11437) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17721) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25925) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4838) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22303) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11576) * $signed(input_fmap_119[7:0]) +
	( 16'sd 31680) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13287) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27202) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2494) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11490) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31492) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24425) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17909) * $signed(input_fmap_127[7:0]) +
	( 16'sd 27011) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18629) * $signed(input_fmap_130[7:0]) +
	( 15'sd 9056) * $signed(input_fmap_131[7:0]) +
	( 16'sd 30343) * $signed(input_fmap_132[7:0]) +
	( 16'sd 20046) * $signed(input_fmap_133[7:0]) +
	( 16'sd 22120) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28544) * $signed(input_fmap_135[7:0]) +
	( 16'sd 27808) * $signed(input_fmap_136[7:0]) +
	( 13'sd 2520) * $signed(input_fmap_137[7:0]) +
	( 13'sd 3384) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14845) * $signed(input_fmap_139[7:0]) +
	( 16'sd 21430) * $signed(input_fmap_140[7:0]) +
	( 15'sd 9205) * $signed(input_fmap_141[7:0]) +
	( 15'sd 10920) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2110) * $signed(input_fmap_144[7:0]) +
	( 16'sd 30950) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19591) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19084) * $signed(input_fmap_147[7:0]) +
	( 14'sd 5486) * $signed(input_fmap_148[7:0]) +
	( 15'sd 13495) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23744) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28640) * $signed(input_fmap_151[7:0]) +
	( 16'sd 29022) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10579) * $signed(input_fmap_153[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_154[7:0]) +
	( 15'sd 8574) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14447) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13807) * $signed(input_fmap_157[7:0]) +
	( 15'sd 10018) * $signed(input_fmap_158[7:0]) +
	( 12'sd 1779) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11080) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28546) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27965) * $signed(input_fmap_162[7:0]) +
	( 16'sd 19553) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8750) * $signed(input_fmap_164[7:0]) +
	( 15'sd 13296) * $signed(input_fmap_165[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_167[7:0]) +
	( 16'sd 22399) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30459) * $signed(input_fmap_169[7:0]) +
	( 15'sd 13749) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31186) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4980) * $signed(input_fmap_172[7:0]) +
	( 16'sd 16571) * $signed(input_fmap_173[7:0]) +
	( 16'sd 22805) * $signed(input_fmap_174[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_175[7:0]) +
	( 11'sd 853) * $signed(input_fmap_176[7:0]) +
	( 16'sd 20358) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6944) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29481) * $signed(input_fmap_180[7:0]) +
	( 16'sd 24138) * $signed(input_fmap_181[7:0]) +
	( 16'sd 17768) * $signed(input_fmap_182[7:0]) +
	( 9'sd 178) * $signed(input_fmap_183[7:0]) +
	( 11'sd 549) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5747) * $signed(input_fmap_185[7:0]) +
	( 16'sd 31759) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28987) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12149) * $signed(input_fmap_188[7:0]) +
	( 16'sd 16852) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27666) * $signed(input_fmap_190[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_191[7:0]) +
	( 15'sd 8392) * $signed(input_fmap_192[7:0]) +
	( 12'sd 1919) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29381) * $signed(input_fmap_194[7:0]) +
	( 16'sd 16475) * $signed(input_fmap_195[7:0]) +
	( 15'sd 10299) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25327) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18791) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13742) * $signed(input_fmap_200[7:0]) +
	( 16'sd 24809) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17704) * $signed(input_fmap_202[7:0]) +
	( 15'sd 15755) * $signed(input_fmap_203[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29589) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7620) * $signed(input_fmap_207[7:0]) +
	( 14'sd 5617) * $signed(input_fmap_208[7:0]) +
	( 14'sd 4705) * $signed(input_fmap_209[7:0]) +
	( 16'sd 21739) * $signed(input_fmap_210[7:0]) +
	( 16'sd 27900) * $signed(input_fmap_211[7:0]) +
	( 16'sd 20054) * $signed(input_fmap_212[7:0]) +
	( 15'sd 14543) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20188) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7831) * $signed(input_fmap_215[7:0]) +
	( 16'sd 21639) * $signed(input_fmap_216[7:0]) +
	( 14'sd 4939) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_218[7:0]) +
	( 16'sd 27009) * $signed(input_fmap_219[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12187) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5840) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_223[7:0]) +
	( 14'sd 5001) * $signed(input_fmap_224[7:0]) +
	( 16'sd 21012) * $signed(input_fmap_225[7:0]) +
	( 15'sd 13566) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18381) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17480) * $signed(input_fmap_229[7:0]) +
	( 15'sd 12657) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18083) * $signed(input_fmap_232[7:0]) +
	( 14'sd 4387) * $signed(input_fmap_233[7:0]) +
	( 15'sd 8769) * $signed(input_fmap_234[7:0]) +
	( 15'sd 15582) * $signed(input_fmap_235[7:0]) +
	( 16'sd 21541) * $signed(input_fmap_236[7:0]) +
	( 16'sd 30027) * $signed(input_fmap_237[7:0]) +
	( 15'sd 9084) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20623) * $signed(input_fmap_239[7:0]) +
	( 16'sd 21271) * $signed(input_fmap_240[7:0]) +
	( 15'sd 11629) * $signed(input_fmap_241[7:0]) +
	( 14'sd 6539) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25025) * $signed(input_fmap_243[7:0]) +
	( 16'sd 26893) * $signed(input_fmap_244[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_245[7:0]) +
	( 16'sd 27323) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18779) * $signed(input_fmap_247[7:0]) +
	( 16'sd 17022) * $signed(input_fmap_248[7:0]) +
	( 11'sd 520) * $signed(input_fmap_249[7:0]) +
	( 16'sd 21259) * $signed(input_fmap_250[7:0]) +
	( 16'sd 24836) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13487) * $signed(input_fmap_252[7:0]) +
	( 16'sd 26270) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_254[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_125;
assign conv_mac_125 = 
	( 15'sd 13732) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5925) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30406) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24250) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12165) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10326) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14971) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26959) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29156) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30786) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1905) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23528) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21387) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21076) * $signed(input_fmap_14[7:0]) +
	( 11'sd 569) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26122) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9308) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16984) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5158) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13955) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27342) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31406) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9687) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29104) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12824) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32089) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26442) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25747) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3012) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26423) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24285) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7936) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30712) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28343) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25168) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27310) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30591) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24466) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21425) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23644) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23364) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21019) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6350) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10551) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12710) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6744) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29877) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1950) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17877) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29643) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27323) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31272) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6854) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13069) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23754) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19693) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25973) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27955) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32500) * $signed(input_fmap_63[7:0]) +
	( 10'sd 459) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28759) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25331) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23757) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21931) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27519) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4706) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13990) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2481) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15660) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30715) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16239) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21423) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4501) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4357) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15634) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13219) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4354) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16493) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9663) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26094) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9585) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7761) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7749) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2230) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20959) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1452) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3859) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17430) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6205) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8750) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6037) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12252) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17395) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10777) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26060) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8701) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13703) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23937) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29870) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1816) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3630) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24441) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25725) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27370) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31601) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27515) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19887) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15151) * $signed(input_fmap_116[7:0]) +
	( 11'sd 776) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10234) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31875) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24444) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28484) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21429) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4182) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9903) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19042) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17568) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23085) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24481) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1930) * $signed(input_fmap_130[7:0]) +
	( 16'sd 32007) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14601) * $signed(input_fmap_132[7:0]) +
	( 12'sd 1882) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10175) * $signed(input_fmap_135[7:0]) +
	( 15'sd 14282) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13790) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17929) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8499) * $signed(input_fmap_139[7:0]) +
	( 13'sd 2926) * $signed(input_fmap_140[7:0]) +
	( 16'sd 23261) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11570) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4481) * $signed(input_fmap_143[7:0]) +
	( 16'sd 23738) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27829) * $signed(input_fmap_145[7:0]) +
	( 14'sd 5424) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14944) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20602) * $signed(input_fmap_148[7:0]) +
	( 13'sd 3623) * $signed(input_fmap_149[7:0]) +
	( 16'sd 17793) * $signed(input_fmap_150[7:0]) +
	( 15'sd 13434) * $signed(input_fmap_151[7:0]) +
	( 15'sd 12263) * $signed(input_fmap_152[7:0]) +
	( 16'sd 20173) * $signed(input_fmap_153[7:0]) +
	( 16'sd 32717) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5169) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28343) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30842) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28518) * $signed(input_fmap_158[7:0]) +
	( 15'sd 15994) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24710) * $signed(input_fmap_160[7:0]) +
	( 15'sd 15367) * $signed(input_fmap_161[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20258) * $signed(input_fmap_163[7:0]) +
	( 16'sd 21472) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4569) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2083) * $signed(input_fmap_166[7:0]) +
	( 14'sd 6802) * $signed(input_fmap_167[7:0]) +
	( 16'sd 24350) * $signed(input_fmap_168[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23031) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30368) * $signed(input_fmap_171[7:0]) +
	( 16'sd 26915) * $signed(input_fmap_172[7:0]) +
	( 16'sd 28325) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27096) * $signed(input_fmap_174[7:0]) +
	( 16'sd 19411) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15258) * $signed(input_fmap_177[7:0]) +
	( 15'sd 8241) * $signed(input_fmap_178[7:0]) +
	( 15'sd 9372) * $signed(input_fmap_179[7:0]) +
	( 14'sd 5180) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16736) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_183[7:0]) +
	( 13'sd 3388) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18833) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25172) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29268) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25998) * $signed(input_fmap_189[7:0]) +
	( 16'sd 32004) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26612) * $signed(input_fmap_191[7:0]) +
	( 14'sd 6904) * $signed(input_fmap_192[7:0]) +
	( 16'sd 21536) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13188) * $signed(input_fmap_195[7:0]) +
	( 16'sd 31952) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19848) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12385) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15832) * $signed(input_fmap_200[7:0]) +
	( 16'sd 17292) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2417) * $signed(input_fmap_202[7:0]) +
	( 16'sd 17919) * $signed(input_fmap_203[7:0]) +
	( 16'sd 22187) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_205[7:0]) +
	( 16'sd 26665) * $signed(input_fmap_206[7:0]) +
	( 14'sd 4822) * $signed(input_fmap_207[7:0]) +
	( 16'sd 27558) * $signed(input_fmap_208[7:0]) +
	( 16'sd 27320) * $signed(input_fmap_209[7:0]) +
	( 16'sd 22801) * $signed(input_fmap_210[7:0]) +
	( 16'sd 22633) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17700) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1695) * $signed(input_fmap_213[7:0]) +
	( 15'sd 13548) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22689) * $signed(input_fmap_215[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_216[7:0]) +
	( 14'sd 6047) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26754) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10959) * $signed(input_fmap_219[7:0]) +
	( 14'sd 7829) * $signed(input_fmap_220[7:0]) +
	( 16'sd 26603) * $signed(input_fmap_221[7:0]) +
	( 16'sd 24140) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25411) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12689) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14511) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10698) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2058) * $signed(input_fmap_227[7:0]) +
	( 15'sd 15795) * $signed(input_fmap_228[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_229[7:0]) +
	( 16'sd 25187) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18538) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29563) * $signed(input_fmap_232[7:0]) +
	( 15'sd 9011) * $signed(input_fmap_233[7:0]) +
	( 16'sd 25957) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22763) * $signed(input_fmap_235[7:0]) +
	( 16'sd 21023) * $signed(input_fmap_236[7:0]) +
	( 10'sd 321) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5185) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22659) * $signed(input_fmap_239[7:0]) +
	( 14'sd 7782) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15833) * $signed(input_fmap_241[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_242[7:0]) +
	( 14'sd 4842) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28759) * $signed(input_fmap_244[7:0]) +
	( 16'sd 20618) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11004) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20129) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18114) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30332) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25648) * $signed(input_fmap_250[7:0]) +
	( 16'sd 17414) * $signed(input_fmap_251[7:0]) +
	( 16'sd 21767) * $signed(input_fmap_252[7:0]) +
	( 15'sd 12604) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20239) * $signed(input_fmap_254[7:0]) +
	( 16'sd 21569) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_126;
assign conv_mac_126 = 
	( 15'sd 16355) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28860) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8779) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2647) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21649) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13143) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26068) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11546) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13838) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29811) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25971) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19901) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21316) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28226) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30086) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24011) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27137) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18993) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18538) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18681) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12668) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32453) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15084) * $signed(input_fmap_27[7:0]) +
	( 16'sd 21716) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13766) * $signed(input_fmap_29[7:0]) +
	( 7'sd 52) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30649) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26947) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1700) * $signed(input_fmap_33[7:0]) +
	( 12'sd 2044) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18491) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5753) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16554) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21360) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7218) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10342) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22624) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24274) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22259) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9855) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22366) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20213) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30020) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14033) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15847) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9924) * $signed(input_fmap_52[7:0]) +
	( 14'sd 8073) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3503) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24588) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20903) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16295) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22080) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24128) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21043) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24268) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17673) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31384) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11742) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21672) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6917) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29881) * $signed(input_fmap_71[7:0]) +
	( 15'sd 8448) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19130) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20653) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14277) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16404) * $signed(input_fmap_77[7:0]) +
	( 16'sd 16837) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18061) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10257) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11561) * $signed(input_fmap_81[7:0]) +
	( 11'sd 950) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1911) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19964) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27575) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24451) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16709) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30694) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30067) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10286) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25422) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9309) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28585) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14652) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24880) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15025) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29674) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30013) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26669) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23293) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19062) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3575) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30714) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19439) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9993) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15703) * $signed(input_fmap_109[7:0]) +
	( 16'sd 26889) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6134) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9600) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7217) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15703) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24844) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29249) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9147) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11763) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20134) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26593) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26185) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16920) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_123[7:0]) +
	( 11'sd 1005) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29832) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_127[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_128[7:0]) +
	( 14'sd 6967) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14898) * $signed(input_fmap_130[7:0]) +
	( 16'sd 29870) * $signed(input_fmap_131[7:0]) +
	( 16'sd 16952) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16676) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2906) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20661) * $signed(input_fmap_135[7:0]) +
	( 16'sd 24771) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26522) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11688) * $signed(input_fmap_138[7:0]) +
	( 14'sd 7552) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3313) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31054) * $signed(input_fmap_141[7:0]) +
	( 16'sd 26608) * $signed(input_fmap_142[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6872) * $signed(input_fmap_144[7:0]) +
	( 15'sd 13377) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15669) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24902) * $signed(input_fmap_147[7:0]) +
	( 12'sd 1585) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27009) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18670) * $signed(input_fmap_150[7:0]) +
	( 16'sd 29707) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23474) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17190) * $signed(input_fmap_153[7:0]) +
	( 16'sd 18232) * $signed(input_fmap_154[7:0]) +
	( 16'sd 18073) * $signed(input_fmap_155[7:0]) +
	( 12'sd 1834) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13474) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25395) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14408) * $signed(input_fmap_159[7:0]) +
	( 16'sd 25803) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_162[7:0]) +
	( 12'sd 1724) * $signed(input_fmap_163[7:0]) +
	( 16'sd 18150) * $signed(input_fmap_164[7:0]) +
	( 14'sd 6333) * $signed(input_fmap_165[7:0]) +
	( 14'sd 5739) * $signed(input_fmap_166[7:0]) +
	( 14'sd 6559) * $signed(input_fmap_167[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20265) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11217) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12279) * $signed(input_fmap_171[7:0]) +
	( 16'sd 17419) * $signed(input_fmap_172[7:0]) +
	( 16'sd 28523) * $signed(input_fmap_173[7:0]) +
	( 16'sd 30213) * $signed(input_fmap_174[7:0]) +
	( 16'sd 16828) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20927) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_177[7:0]) +
	( 16'sd 29965) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6008) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24838) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18606) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10220) * $signed(input_fmap_182[7:0]) +
	( 16'sd 32100) * $signed(input_fmap_183[7:0]) +
	( 15'sd 12382) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22711) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17736) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25246) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2176) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_189[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14276) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14248) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19772) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21970) * $signed(input_fmap_194[7:0]) +
	( 15'sd 15629) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12225) * $signed(input_fmap_196[7:0]) +
	( 14'sd 6239) * $signed(input_fmap_197[7:0]) +
	( 15'sd 15626) * $signed(input_fmap_198[7:0]) +
	( 13'sd 3264) * $signed(input_fmap_199[7:0]) +
	( 15'sd 14544) * $signed(input_fmap_200[7:0]) +
	( 16'sd 17613) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21826) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30456) * $signed(input_fmap_203[7:0]) +
	( 16'sd 23289) * $signed(input_fmap_204[7:0]) +
	( 15'sd 9913) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27438) * $signed(input_fmap_206[7:0]) +
	( 15'sd 8582) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17583) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24115) * $signed(input_fmap_209[7:0]) +
	( 16'sd 20535) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10428) * $signed(input_fmap_211[7:0]) +
	( 15'sd 10191) * $signed(input_fmap_212[7:0]) +
	( 16'sd 18799) * $signed(input_fmap_213[7:0]) +
	( 14'sd 4972) * $signed(input_fmap_214[7:0]) +
	( 13'sd 3297) * $signed(input_fmap_215[7:0]) +
	( 15'sd 12430) * $signed(input_fmap_216[7:0]) +
	( 13'sd 3630) * $signed(input_fmap_217[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20790) * $signed(input_fmap_219[7:0]) +
	( 16'sd 17000) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15644) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3106) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12747) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14496) * $signed(input_fmap_224[7:0]) +
	( 13'sd 4074) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22192) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9326) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22885) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6992) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18872) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3249) * $signed(input_fmap_231[7:0]) +
	( 16'sd 19964) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_233[7:0]) +
	( 16'sd 26283) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26055) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5473) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19528) * $signed(input_fmap_237[7:0]) +
	( 16'sd 20970) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23187) * $signed(input_fmap_239[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21808) * $signed(input_fmap_241[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_242[7:0]) +
	( 16'sd 29297) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18947) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30456) * $signed(input_fmap_245[7:0]) +
	( 16'sd 27854) * $signed(input_fmap_246[7:0]) +
	( 14'sd 5585) * $signed(input_fmap_247[7:0]) +
	( 13'sd 2715) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25715) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24997) * $signed(input_fmap_250[7:0]) +
	( 16'sd 31270) * $signed(input_fmap_251[7:0]) +
	( 11'sd 948) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2834) * $signed(input_fmap_253[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_254[7:0]) +
	( 15'sd 12077) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_127;
assign conv_mac_127 = 
	( 15'sd 10074) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16963) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12840) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5241) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24135) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14861) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32447) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9816) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20419) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28723) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9708) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31053) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32107) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13126) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23907) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31552) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25687) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26286) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21820) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4777) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23580) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24548) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32299) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27234) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7134) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_28[7:0]) +
	( 11'sd 830) * $signed(input_fmap_29[7:0]) +
	( 8'sd 66) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12888) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5607) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30760) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3741) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25464) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3344) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18144) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18688) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13150) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10754) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25945) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16214) * $signed(input_fmap_43[7:0]) +
	( 16'sd 31723) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24445) * $signed(input_fmap_45[7:0]) +
	( 7'sd 41) * $signed(input_fmap_46[7:0]) +
	( 15'sd 16129) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2782) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2563) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19348) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12840) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12546) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9816) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23512) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31752) * $signed(input_fmap_56[7:0]) +
	( 15'sd 16370) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17052) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12308) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17619) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2419) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4903) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27621) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12591) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14214) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11284) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20767) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28627) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13811) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12477) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13518) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18397) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13551) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26204) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15544) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14819) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29907) * $signed(input_fmap_83[7:0]) +
	( 10'sd 508) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27922) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23945) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31883) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13966) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9378) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23601) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14662) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5984) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9668) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11160) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16404) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24301) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_97[7:0]) +
	( 7'sd 36) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13103) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16961) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32002) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19099) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19717) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30914) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19004) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30983) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9557) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1445) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13010) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8716) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14884) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30583) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16666) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17137) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2505) * $signed(input_fmap_117[7:0]) +
	( 11'sd 566) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14588) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11898) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17163) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3224) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18168) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18664) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1553) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19989) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13165) * $signed(input_fmap_127[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_128[7:0]) +
	( 16'sd 23316) * $signed(input_fmap_129[7:0]) +
	( 13'sd 2615) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24225) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10203) * $signed(input_fmap_132[7:0]) +
	( 11'sd 901) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21105) * $signed(input_fmap_134[7:0]) +
	( 16'sd 29473) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21872) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25308) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29523) * $signed(input_fmap_138[7:0]) +
	( 15'sd 15073) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15072) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22350) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30762) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12813) * $signed(input_fmap_143[7:0]) +
	( 15'sd 14847) * $signed(input_fmap_144[7:0]) +
	( 16'sd 18639) * $signed(input_fmap_145[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18684) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11696) * $signed(input_fmap_148[7:0]) +
	( 15'sd 11346) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25479) * $signed(input_fmap_150[7:0]) +
	( 14'sd 7142) * $signed(input_fmap_151[7:0]) +
	( 16'sd 28226) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10243) * $signed(input_fmap_153[7:0]) +
	( 15'sd 9422) * $signed(input_fmap_154[7:0]) +
	( 10'sd 399) * $signed(input_fmap_155[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_156[7:0]) +
	( 16'sd 17881) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4667) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14855) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31757) * $signed(input_fmap_160[7:0]) +
	( 16'sd 27265) * $signed(input_fmap_161[7:0]) +
	( 16'sd 17375) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15090) * $signed(input_fmap_163[7:0]) +
	( 16'sd 16486) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30107) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2427) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13004) * $signed(input_fmap_167[7:0]) +
	( 16'sd 16421) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_169[7:0]) +
	( 15'sd 8525) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31166) * $signed(input_fmap_171[7:0]) +
	( 16'sd 24208) * $signed(input_fmap_172[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_173[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_174[7:0]) +
	( 16'sd 24436) * $signed(input_fmap_175[7:0]) +
	( 16'sd 31127) * $signed(input_fmap_176[7:0]) +
	( 15'sd 14802) * $signed(input_fmap_177[7:0]) +
	( 16'sd 26826) * $signed(input_fmap_178[7:0]) +
	( 16'sd 29446) * $signed(input_fmap_179[7:0]) +
	( 15'sd 13892) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15434) * $signed(input_fmap_181[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12091) * $signed(input_fmap_183[7:0]) +
	( 14'sd 4967) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17933) * $signed(input_fmap_185[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_186[7:0]) +
	( 15'sd 12175) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17607) * $signed(input_fmap_188[7:0]) +
	( 15'sd 15337) * $signed(input_fmap_189[7:0]) +
	( 16'sd 32618) * $signed(input_fmap_190[7:0]) +
	( 16'sd 21212) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20624) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_194[7:0]) +
	( 15'sd 12394) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20175) * $signed(input_fmap_196[7:0]) +
	( 14'sd 7715) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27051) * $signed(input_fmap_198[7:0]) +
	( 16'sd 26801) * $signed(input_fmap_199[7:0]) +
	( 16'sd 16766) * $signed(input_fmap_200[7:0]) +
	( 16'sd 25263) * $signed(input_fmap_201[7:0]) +
	( 12'sd 1949) * $signed(input_fmap_202[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15034) * $signed(input_fmap_204[7:0]) +
	( 16'sd 27584) * $signed(input_fmap_205[7:0]) +
	( 14'sd 7327) * $signed(input_fmap_206[7:0]) +
	( 16'sd 32270) * $signed(input_fmap_207[7:0]) +
	( 16'sd 32176) * $signed(input_fmap_208[7:0]) +
	( 16'sd 17998) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31787) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20418) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_212[7:0]) +
	( 15'sd 8346) * $signed(input_fmap_213[7:0]) +
	( 15'sd 8751) * $signed(input_fmap_214[7:0]) +
	( 16'sd 26321) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17848) * $signed(input_fmap_216[7:0]) +
	( 15'sd 11201) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8943) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19617) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1745) * $signed(input_fmap_220[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28276) * $signed(input_fmap_222[7:0]) +
	( 12'sd 2037) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17621) * $signed(input_fmap_224[7:0]) +
	( 16'sd 30294) * $signed(input_fmap_225[7:0]) +
	( 15'sd 15004) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_227[7:0]) +
	( 16'sd 20417) * $signed(input_fmap_228[7:0]) +
	( 16'sd 22662) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14747) * $signed(input_fmap_230[7:0]) +
	( 8'sd 102) * $signed(input_fmap_231[7:0]) +
	( 16'sd 21956) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27029) * $signed(input_fmap_233[7:0]) +
	( 16'sd 26566) * $signed(input_fmap_234[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_235[7:0]) +
	( 16'sd 16559) * $signed(input_fmap_236[7:0]) +
	( 16'sd 25826) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28379) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19650) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23174) * $signed(input_fmap_240[7:0]) +
	( 15'sd 10573) * $signed(input_fmap_241[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_242[7:0]) +
	( 16'sd 16477) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20335) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19412) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1810) * $signed(input_fmap_246[7:0]) +
	( 14'sd 4401) * $signed(input_fmap_247[7:0]) +
	( 15'sd 16097) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3959) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12778) * $signed(input_fmap_251[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24634) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23700) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_128;
assign conv_mac_128 = 
	( 16'sd 30887) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24974) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2286) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10487) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27145) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14428) * $signed(input_fmap_6[7:0]) +
	( 14'sd 8127) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9269) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31150) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6208) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5895) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7822) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5156) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7769) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15638) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8929) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4335) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26351) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31376) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22050) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12171) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18441) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31918) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27274) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23197) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27062) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7109) * $signed(input_fmap_29[7:0]) +
	( 14'sd 8017) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3794) * $signed(input_fmap_31[7:0]) +
	( 11'sd 721) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24218) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30498) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4553) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25373) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17739) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2506) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15691) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6812) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5285) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21842) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32302) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20162) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29859) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6615) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28383) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31047) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20825) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4630) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18892) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23133) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17874) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20078) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4111) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17136) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3183) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_61[7:0]) +
	( 10'sd 458) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8699) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30864) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4691) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15801) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26542) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6224) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10952) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5344) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12156) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3577) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6520) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20423) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14318) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18832) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19405) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18981) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5613) * $signed(input_fmap_80[7:0]) +
	( 10'sd 496) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12818) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20022) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5042) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14727) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10653) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16537) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15799) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24259) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15703) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5359) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27524) * $signed(input_fmap_92[7:0]) +
	( 16'sd 29700) * $signed(input_fmap_93[7:0]) +
	( 15'sd 8252) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9317) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5925) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11282) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6462) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12162) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31984) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8520) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22867) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28934) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17571) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8743) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16975) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4192) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1145) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9586) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10968) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21751) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26391) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31124) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1052) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11890) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30641) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31922) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22688) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12877) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31226) * $signed(input_fmap_121[7:0]) +
	( 16'sd 16956) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9698) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3163) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10990) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25663) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5952) * $signed(input_fmap_127[7:0]) +
	( 15'sd 10764) * $signed(input_fmap_128[7:0]) +
	( 9'sd 201) * $signed(input_fmap_129[7:0]) +
	( 16'sd 24965) * $signed(input_fmap_130[7:0]) +
	( 16'sd 30725) * $signed(input_fmap_131[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_132[7:0]) +
	( 14'sd 6400) * $signed(input_fmap_133[7:0]) +
	( 16'sd 22966) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20589) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25481) * $signed(input_fmap_136[7:0]) +
	( 15'sd 10065) * $signed(input_fmap_137[7:0]) +
	( 14'sd 4607) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24816) * $signed(input_fmap_139[7:0]) +
	( 15'sd 8677) * $signed(input_fmap_140[7:0]) +
	( 11'sd 546) * $signed(input_fmap_141[7:0]) +
	( 16'sd 17009) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31182) * $signed(input_fmap_143[7:0]) +
	( 16'sd 30655) * $signed(input_fmap_144[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_145[7:0]) +
	( 16'sd 20110) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26201) * $signed(input_fmap_148[7:0]) +
	( 12'sd 1834) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15330) * $signed(input_fmap_150[7:0]) +
	( 16'sd 32016) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24955) * $signed(input_fmap_152[7:0]) +
	( 15'sd 9754) * $signed(input_fmap_153[7:0]) +
	( 12'sd 1327) * $signed(input_fmap_154[7:0]) +
	( 15'sd 15483) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13114) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22849) * $signed(input_fmap_157[7:0]) +
	( 16'sd 30869) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20584) * $signed(input_fmap_159[7:0]) +
	( 16'sd 20484) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4577) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_162[7:0]) +
	( 14'sd 5331) * $signed(input_fmap_163[7:0]) +
	( 16'sd 22307) * $signed(input_fmap_164[7:0]) +
	( 16'sd 21332) * $signed(input_fmap_165[7:0]) +
	( 16'sd 16536) * $signed(input_fmap_166[7:0]) +
	( 13'sd 3289) * $signed(input_fmap_167[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17021) * $signed(input_fmap_169[7:0]) +
	( 15'sd 10168) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3922) * $signed(input_fmap_171[7:0]) +
	( 16'sd 17034) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29880) * $signed(input_fmap_173[7:0]) +
	( 15'sd 13642) * $signed(input_fmap_174[7:0]) +
	( 15'sd 8654) * $signed(input_fmap_175[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31720) * $signed(input_fmap_177[7:0]) +
	( 16'sd 21677) * $signed(input_fmap_178[7:0]) +
	( 15'sd 12628) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27127) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11009) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19169) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30899) * $signed(input_fmap_183[7:0]) +
	( 16'sd 27681) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25474) * $signed(input_fmap_185[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2527) * $signed(input_fmap_187[7:0]) +
	( 16'sd 16706) * $signed(input_fmap_188[7:0]) +
	( 16'sd 31120) * $signed(input_fmap_189[7:0]) +
	( 12'sd 1543) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_191[7:0]) +
	( 13'sd 2374) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26851) * $signed(input_fmap_193[7:0]) +
	( 12'sd 1816) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25843) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20309) * $signed(input_fmap_196[7:0]) +
	( 16'sd 16443) * $signed(input_fmap_197[7:0]) +
	( 12'sd 1061) * $signed(input_fmap_198[7:0]) +
	( 16'sd 22279) * $signed(input_fmap_199[7:0]) +
	( 16'sd 32282) * $signed(input_fmap_200[7:0]) +
	( 15'sd 10378) * $signed(input_fmap_201[7:0]) +
	( 16'sd 26326) * $signed(input_fmap_202[7:0]) +
	( 16'sd 22341) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32368) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27348) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13092) * $signed(input_fmap_207[7:0]) +
	( 13'sd 2742) * $signed(input_fmap_208[7:0]) +
	( 16'sd 21769) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30542) * $signed(input_fmap_210[7:0]) +
	( 16'sd 31619) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12805) * $signed(input_fmap_212[7:0]) +
	( 16'sd 22457) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23398) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10708) * $signed(input_fmap_215[7:0]) +
	( 14'sd 6139) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32527) * $signed(input_fmap_217[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_218[7:0]) +
	( 15'sd 8768) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25120) * $signed(input_fmap_220[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_221[7:0]) +
	( 16'sd 23176) * $signed(input_fmap_222[7:0]) +
	( 16'sd 18038) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12018) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5053) * $signed(input_fmap_225[7:0]) +
	( 14'sd 4352) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22939) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2332) * $signed(input_fmap_228[7:0]) +
	( 15'sd 16360) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_230[7:0]) +
	( 16'sd 32742) * $signed(input_fmap_231[7:0]) +
	( 14'sd 5840) * $signed(input_fmap_232[7:0]) +
	( 16'sd 25317) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19120) * $signed(input_fmap_234[7:0]) +
	( 15'sd 10608) * $signed(input_fmap_235[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_236[7:0]) +
	( 11'sd 554) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19895) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20885) * $signed(input_fmap_239[7:0]) +
	( 15'sd 14378) * $signed(input_fmap_240[7:0]) +
	( 16'sd 24592) * $signed(input_fmap_241[7:0]) +
	( 16'sd 24273) * $signed(input_fmap_242[7:0]) +
	( 16'sd 20929) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12038) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5747) * $signed(input_fmap_245[7:0]) +
	( 16'sd 16766) * $signed(input_fmap_246[7:0]) +
	( 14'sd 7366) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10276) * $signed(input_fmap_248[7:0]) +
	( 14'sd 5619) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9257) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2274) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2564) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24521) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2547) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14369) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_129;
assign conv_mac_129 = 
	( 16'sd 24221) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_1[7:0]) +
	( 10'sd 358) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10315) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19119) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9061) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21040) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15717) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5258) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3481) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2996) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18897) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1235) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20572) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26775) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11348) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2446) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32617) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5719) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7463) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17946) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26268) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17191) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27347) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17274) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24351) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24065) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32667) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27385) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18046) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25498) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8463) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30395) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17714) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2268) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31623) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7700) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9396) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8320) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21896) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12185) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30925) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13697) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10632) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20517) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19788) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32635) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3732) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15471) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30916) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32667) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22517) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13275) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27311) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13886) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2294) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30934) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8366) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30115) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25934) * $signed(input_fmap_62[7:0]) +
	( 15'sd 16362) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11204) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9948) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5596) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32130) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25530) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16954) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19556) * $signed(input_fmap_71[7:0]) +
	( 10'sd 325) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21863) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14227) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20889) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26907) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21594) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15110) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18586) * $signed(input_fmap_79[7:0]) +
	( 9'sd 196) * $signed(input_fmap_80[7:0]) +
	( 9'sd 231) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21683) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10102) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12144) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8825) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29171) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16828) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30534) * $signed(input_fmap_88[7:0]) +
	( 13'sd 4017) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29589) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28462) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27297) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31690) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7142) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19989) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1341) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31406) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23178) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4618) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24341) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31520) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24849) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18565) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31368) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19441) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3358) * $signed(input_fmap_106[7:0]) +
	( 11'sd 737) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25326) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30007) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1262) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20434) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8760) * $signed(input_fmap_112[7:0]) +
	( 10'sd 258) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8910) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11301) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16381) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8615) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14556) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9623) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27899) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3636) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16733) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29429) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23974) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30924) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18135) * $signed(input_fmap_128[7:0]) +
	( 16'sd 22547) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27379) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1523) * $signed(input_fmap_132[7:0]) +
	( 16'sd 23189) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4803) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21900) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15120) * $signed(input_fmap_136[7:0]) +
	( 15'sd 10214) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27148) * $signed(input_fmap_138[7:0]) +
	( 10'sd 361) * $signed(input_fmap_139[7:0]) +
	( 16'sd 22746) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24809) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12032) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18841) * $signed(input_fmap_144[7:0]) +
	( 16'sd 32377) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15316) * $signed(input_fmap_146[7:0]) +
	( 15'sd 12688) * $signed(input_fmap_147[7:0]) +
	( 16'sd 27550) * $signed(input_fmap_148[7:0]) +
	( 16'sd 24345) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5723) * $signed(input_fmap_150[7:0]) +
	( 16'sd 25448) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23012) * $signed(input_fmap_152[7:0]) +
	( 16'sd 32087) * $signed(input_fmap_153[7:0]) +
	( 13'sd 2157) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13602) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28221) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6304) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9552) * $signed(input_fmap_158[7:0]) +
	( 15'sd 9802) * $signed(input_fmap_159[7:0]) +
	( 16'sd 23378) * $signed(input_fmap_160[7:0]) +
	( 16'sd 30011) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4192) * $signed(input_fmap_162[7:0]) +
	( 11'sd 676) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10084) * $signed(input_fmap_164[7:0]) +
	( 16'sd 26007) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4609) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24531) * $signed(input_fmap_167[7:0]) +
	( 16'sd 24599) * $signed(input_fmap_168[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_169[7:0]) +
	( 16'sd 29257) * $signed(input_fmap_170[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_171[7:0]) +
	( 16'sd 25287) * $signed(input_fmap_172[7:0]) +
	( 16'sd 26819) * $signed(input_fmap_173[7:0]) +
	( 16'sd 31224) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28020) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3636) * $signed(input_fmap_176[7:0]) +
	( 15'sd 13353) * $signed(input_fmap_177[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_178[7:0]) +
	( 16'sd 23381) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28451) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6976) * $signed(input_fmap_181[7:0]) +
	( 16'sd 28526) * $signed(input_fmap_182[7:0]) +
	( 12'sd 1785) * $signed(input_fmap_183[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13983) * $signed(input_fmap_186[7:0]) +
	( 15'sd 14702) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1899) * $signed(input_fmap_188[7:0]) +
	( 16'sd 22136) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20755) * $signed(input_fmap_190[7:0]) +
	( 13'sd 2802) * $signed(input_fmap_191[7:0]) +
	( 16'sd 30451) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28078) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9080) * $signed(input_fmap_194[7:0]) +
	( 16'sd 32228) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25069) * $signed(input_fmap_197[7:0]) +
	( 16'sd 17996) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5619) * $signed(input_fmap_199[7:0]) +
	( 16'sd 21925) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18363) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_202[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_203[7:0]) +
	( 11'sd 841) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31996) * $signed(input_fmap_205[7:0]) +
	( 16'sd 18374) * $signed(input_fmap_206[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17478) * $signed(input_fmap_208[7:0]) +
	( 15'sd 15972) * $signed(input_fmap_209[7:0]) +
	( 14'sd 6466) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30947) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17973) * $signed(input_fmap_212[7:0]) +
	( 15'sd 15456) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20074) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23720) * $signed(input_fmap_215[7:0]) +
	( 16'sd 29157) * $signed(input_fmap_216[7:0]) +
	( 14'sd 4246) * $signed(input_fmap_217[7:0]) +
	( 11'sd 899) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14644) * $signed(input_fmap_219[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_220[7:0]) +
	( 15'sd 10519) * $signed(input_fmap_221[7:0]) +
	( 16'sd 26956) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15569) * $signed(input_fmap_223[7:0]) +
	( 13'sd 2448) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18795) * $signed(input_fmap_225[7:0]) +
	( 15'sd 12343) * $signed(input_fmap_226[7:0]) +
	( 16'sd 26479) * $signed(input_fmap_227[7:0]) +
	( 15'sd 13070) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6216) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28301) * $signed(input_fmap_230[7:0]) +
	( 16'sd 26789) * $signed(input_fmap_231[7:0]) +
	( 15'sd 13369) * $signed(input_fmap_232[7:0]) +
	( 13'sd 2753) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15952) * $signed(input_fmap_234[7:0]) +
	( 15'sd 10987) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25241) * $signed(input_fmap_236[7:0]) +
	( 16'sd 31731) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22354) * $signed(input_fmap_238[7:0]) +
	( 16'sd 32261) * $signed(input_fmap_239[7:0]) +
	( 16'sd 24190) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5776) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29621) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13328) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24220) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6282) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20140) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13522) * $signed(input_fmap_247[7:0]) +
	( 16'sd 19848) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3773) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7912) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18547) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27813) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29979) * $signed(input_fmap_253[7:0]) +
	( 15'sd 11580) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23245) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_130;
assign conv_mac_130 = 
	( 16'sd 18895) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14980) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4837) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6701) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8904) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10472) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3499) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13417) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30381) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21534) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1794) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29781) * $signed(input_fmap_16[7:0]) +
	( 9'sd 204) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13314) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10182) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24943) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28214) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4378) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7273) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1481) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29713) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24493) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22716) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20074) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15785) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25810) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14822) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1936) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21172) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21209) * $signed(input_fmap_36[7:0]) +
	( 11'sd 710) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10367) * $signed(input_fmap_38[7:0]) +
	( 16'sd 21876) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27481) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18806) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15154) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6893) * $signed(input_fmap_43[7:0]) +
	( 13'sd 4092) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26476) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3859) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5450) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5923) * $signed(input_fmap_48[7:0]) +
	( 13'sd 4043) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18134) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12733) * $signed(input_fmap_51[7:0]) +
	( 12'sd 2024) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12235) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7077) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30863) * $signed(input_fmap_55[7:0]) +
	( 10'sd 442) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32462) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12460) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15774) * $signed(input_fmap_59[7:0]) +
	( 11'sd 989) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23605) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10846) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12409) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21145) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18447) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30280) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17604) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23609) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32604) * $signed(input_fmap_69[7:0]) +
	( 15'sd 16359) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24331) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15442) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3763) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25972) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13052) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7673) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3599) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26298) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20820) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14438) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11130) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6008) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21247) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16791) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25855) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30851) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10638) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24396) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7088) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4096) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13571) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26005) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27745) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8417) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1256) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17171) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18868) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4662) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32577) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6459) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3705) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10872) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14213) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13599) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18328) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2886) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5691) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16134) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21453) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27660) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3039) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18226) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20885) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4424) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30628) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30911) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17403) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24480) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31906) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7625) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31345) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29806) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22218) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19383) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7823) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29920) * $signed(input_fmap_128[7:0]) +
	( 14'sd 6618) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22189) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31618) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5213) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10444) * $signed(input_fmap_133[7:0]) +
	( 14'sd 6096) * $signed(input_fmap_134[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17999) * $signed(input_fmap_136[7:0]) +
	( 16'sd 23718) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_138[7:0]) +
	( 15'sd 12648) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3028) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13594) * $signed(input_fmap_141[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5313) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19300) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25170) * $signed(input_fmap_145[7:0]) +
	( 16'sd 17668) * $signed(input_fmap_146[7:0]) +
	( 14'sd 5751) * $signed(input_fmap_147[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27829) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_150[7:0]) +
	( 16'sd 32276) * $signed(input_fmap_151[7:0]) +
	( 15'sd 8330) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10900) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20079) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14805) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5453) * $signed(input_fmap_157[7:0]) +
	( 16'sd 22073) * $signed(input_fmap_158[7:0]) +
	( 15'sd 13435) * $signed(input_fmap_159[7:0]) +
	( 15'sd 15621) * $signed(input_fmap_160[7:0]) +
	( 13'sd 3387) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2326) * $signed(input_fmap_162[7:0]) +
	( 14'sd 5270) * $signed(input_fmap_163[7:0]) +
	( 13'sd 2257) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22914) * $signed(input_fmap_165[7:0]) +
	( 9'sd 243) * $signed(input_fmap_166[7:0]) +
	( 12'sd 1072) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4507) * $signed(input_fmap_168[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_169[7:0]) +
	( 15'sd 8375) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14187) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19052) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26397) * $signed(input_fmap_174[7:0]) +
	( 16'sd 23632) * $signed(input_fmap_175[7:0]) +
	( 13'sd 2902) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15854) * $signed(input_fmap_177[7:0]) +
	( 16'sd 16557) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25471) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23243) * $signed(input_fmap_180[7:0]) +
	( 15'sd 16211) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19468) * $signed(input_fmap_182[7:0]) +
	( 16'sd 22241) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13896) * $signed(input_fmap_184[7:0]) +
	( 15'sd 10097) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26809) * $signed(input_fmap_186[7:0]) +
	( 16'sd 23446) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21426) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2309) * $signed(input_fmap_189[7:0]) +
	( 16'sd 18327) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24320) * $signed(input_fmap_191[7:0]) +
	( 9'sd 155) * $signed(input_fmap_192[7:0]) +
	( 16'sd 18494) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29597) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19453) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11337) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1437) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10377) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5797) * $signed(input_fmap_199[7:0]) +
	( 16'sd 28100) * $signed(input_fmap_200[7:0]) +
	( 16'sd 31507) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14888) * $signed(input_fmap_202[7:0]) +
	( 15'sd 15331) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4851) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28267) * $signed(input_fmap_205[7:0]) +
	( 15'sd 14668) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18192) * $signed(input_fmap_207[7:0]) +
	( 16'sd 19159) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3913) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31174) * $signed(input_fmap_210[7:0]) +
	( 16'sd 21170) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1855) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28212) * $signed(input_fmap_213[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_215[7:0]) +
	( 15'sd 15053) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10920) * $signed(input_fmap_217[7:0]) +
	( 12'sd 1547) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3857) * $signed(input_fmap_219[7:0]) +
	( 13'sd 3574) * $signed(input_fmap_220[7:0]) +
	( 14'sd 4904) * $signed(input_fmap_221[7:0]) +
	( 14'sd 7021) * $signed(input_fmap_222[7:0]) +
	( 16'sd 16452) * $signed(input_fmap_223[7:0]) +
	( 15'sd 15818) * $signed(input_fmap_224[7:0]) +
	( 16'sd 29453) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18490) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_227[7:0]) +
	( 15'sd 14442) * $signed(input_fmap_228[7:0]) +
	( 16'sd 32639) * $signed(input_fmap_229[7:0]) +
	( 16'sd 19195) * $signed(input_fmap_230[7:0]) +
	( 14'sd 6987) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20729) * $signed(input_fmap_232[7:0]) +
	( 16'sd 30160) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14452) * $signed(input_fmap_234[7:0]) +
	( 15'sd 10657) * $signed(input_fmap_235[7:0]) +
	( 15'sd 13554) * $signed(input_fmap_236[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27311) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9032) * $signed(input_fmap_239[7:0]) +
	( 16'sd 20313) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_242[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28907) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14172) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31838) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18192) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10033) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3190) * $signed(input_fmap_249[7:0]) +
	( 16'sd 29989) * $signed(input_fmap_250[7:0]) +
	( 16'sd 24325) * $signed(input_fmap_251[7:0]) +
	( 15'sd 11165) * $signed(input_fmap_252[7:0]) +
	( 14'sd 4971) * $signed(input_fmap_253[7:0]) +
	( 16'sd 30562) * $signed(input_fmap_254[7:0]) +
	( 14'sd 8147) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_131;
assign conv_mac_131 = 
	( 3'sd 2) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22087) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10250) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24322) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14475) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16770) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2694) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22239) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5060) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16246) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30322) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22049) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29804) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26575) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30174) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18730) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14140) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9194) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21228) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1513) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9900) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15620) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31969) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9635) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23298) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32551) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11564) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6570) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9130) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20178) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23223) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11123) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23274) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26503) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15370) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14953) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15044) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21469) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17120) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7413) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1297) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32025) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7586) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18185) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16866) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4917) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10824) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17807) * $signed(input_fmap_50[7:0]) +
	( 11'sd 585) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17375) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23128) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8571) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_55[7:0]) +
	( 10'sd 384) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17122) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15414) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9239) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3979) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10877) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9502) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29512) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31281) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2187) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31572) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22051) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20625) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2600) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5223) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30037) * $signed(input_fmap_74[7:0]) +
	( 16'sd 26657) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16035) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17884) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30087) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14593) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30909) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4451) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18679) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22013) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11122) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21685) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12506) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3494) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8202) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1170) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12461) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15504) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25022) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6970) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22187) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24671) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18585) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13148) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29202) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9903) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19823) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27570) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6720) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24351) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14116) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18754) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6870) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26621) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3864) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1379) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14661) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4860) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16983) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16923) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22308) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2194) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9800) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27165) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31234) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12212) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8871) * $signed(input_fmap_127[7:0]) +
	( 16'sd 26415) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17155) * $signed(input_fmap_129[7:0]) +
	( 13'sd 3043) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19414) * $signed(input_fmap_131[7:0]) +
	( 15'sd 9991) * $signed(input_fmap_132[7:0]) +
	( 15'sd 13443) * $signed(input_fmap_133[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21309) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_136[7:0]) +
	( 16'sd 23273) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29514) * $signed(input_fmap_138[7:0]) +
	( 4'sd 7) * $signed(input_fmap_139[7:0]) +
	( 14'sd 7657) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3268) * $signed(input_fmap_141[7:0]) +
	( 15'sd 12450) * $signed(input_fmap_142[7:0]) +
	( 16'sd 19906) * $signed(input_fmap_143[7:0]) +
	( 15'sd 14154) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26691) * $signed(input_fmap_145[7:0]) +
	( 14'sd 5466) * $signed(input_fmap_146[7:0]) +
	( 16'sd 20139) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22087) * $signed(input_fmap_148[7:0]) +
	( 16'sd 21733) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18772) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6989) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16606) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17276) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7719) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23479) * $signed(input_fmap_155[7:0]) +
	( 15'sd 12428) * $signed(input_fmap_156[7:0]) +
	( 10'sd 448) * $signed(input_fmap_157[7:0]) +
	( 13'sd 2396) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12169) * $signed(input_fmap_159[7:0]) +
	( 15'sd 9129) * $signed(input_fmap_160[7:0]) +
	( 14'sd 6988) * $signed(input_fmap_161[7:0]) +
	( 14'sd 7982) * $signed(input_fmap_162[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_163[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28824) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9763) * $signed(input_fmap_166[7:0]) +
	( 14'sd 5539) * $signed(input_fmap_167[7:0]) +
	( 16'sd 25514) * $signed(input_fmap_168[7:0]) +
	( 16'sd 29761) * $signed(input_fmap_169[7:0]) +
	( 16'sd 30208) * $signed(input_fmap_170[7:0]) +
	( 14'sd 5443) * $signed(input_fmap_171[7:0]) +
	( 16'sd 32394) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12808) * $signed(input_fmap_173[7:0]) +
	( 15'sd 13767) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1652) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15094) * $signed(input_fmap_176[7:0]) +
	( 16'sd 23095) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_178[7:0]) +
	( 15'sd 12408) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3373) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28777) * $signed(input_fmap_181[7:0]) +
	( 16'sd 23841) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25419) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_184[7:0]) +
	( 16'sd 16611) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23979) * $signed(input_fmap_186[7:0]) +
	( 14'sd 6559) * $signed(input_fmap_187[7:0]) +
	( 15'sd 14260) * $signed(input_fmap_188[7:0]) +
	( 14'sd 4418) * $signed(input_fmap_189[7:0]) +
	( 16'sd 21658) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31779) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12563) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5961) * $signed(input_fmap_193[7:0]) +
	( 16'sd 17073) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25095) * $signed(input_fmap_195[7:0]) +
	( 15'sd 10152) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19501) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29602) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23564) * $signed(input_fmap_199[7:0]) +
	( 16'sd 27796) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18032) * $signed(input_fmap_201[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24374) * $signed(input_fmap_203[7:0]) +
	( 16'sd 30531) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2558) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3610) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25853) * $signed(input_fmap_208[7:0]) +
	( 16'sd 21095) * $signed(input_fmap_209[7:0]) +
	( 15'sd 12589) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20795) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26426) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2552) * $signed(input_fmap_213[7:0]) +
	( 16'sd 25783) * $signed(input_fmap_214[7:0]) +
	( 16'sd 21307) * $signed(input_fmap_215[7:0]) +
	( 16'sd 25206) * $signed(input_fmap_216[7:0]) +
	( 16'sd 20935) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8705) * $signed(input_fmap_218[7:0]) +
	( 15'sd 8514) * $signed(input_fmap_219[7:0]) +
	( 16'sd 18386) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5333) * $signed(input_fmap_221[7:0]) +
	( 16'sd 17064) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15668) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12992) * $signed(input_fmap_224[7:0]) +
	( 11'sd 793) * $signed(input_fmap_225[7:0]) +
	( 16'sd 25072) * $signed(input_fmap_226[7:0]) +
	( 16'sd 31086) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10537) * $signed(input_fmap_228[7:0]) +
	( 13'sd 2745) * $signed(input_fmap_229[7:0]) +
	( 15'sd 10001) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25108) * $signed(input_fmap_231[7:0]) +
	( 16'sd 24584) * $signed(input_fmap_232[7:0]) +
	( 16'sd 19875) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4215) * $signed(input_fmap_234[7:0]) +
	( 16'sd 23017) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_236[7:0]) +
	( 16'sd 24654) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17582) * $signed(input_fmap_238[7:0]) +
	( 15'sd 16146) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19117) * $signed(input_fmap_240[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_241[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_242[7:0]) +
	( 16'sd 27128) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1946) * $signed(input_fmap_244[7:0]) +
	( 11'sd 538) * $signed(input_fmap_245[7:0]) +
	( 15'sd 13452) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_247[7:0]) +
	( 16'sd 28958) * $signed(input_fmap_248[7:0]) +
	( 16'sd 18181) * $signed(input_fmap_249[7:0]) +
	( 16'sd 18171) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13210) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12936) * $signed(input_fmap_252[7:0]) +
	( 16'sd 23781) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31243) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23688) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_132;
assign conv_mac_132 = 
	( 16'sd 17141) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25564) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18977) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18937) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19627) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17556) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31964) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18521) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1193) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25051) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31533) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3922) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13004) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30748) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28658) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8647) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28890) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19293) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15362) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29053) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2438) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11318) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5276) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30263) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20486) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30992) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4118) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_30[7:0]) +
	( 14'sd 8034) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19922) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2690) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9137) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17807) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32601) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20408) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13650) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26597) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11768) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17229) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21580) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31400) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30594) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9838) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5144) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25491) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10943) * $signed(input_fmap_53[7:0]) +
	( 11'sd 566) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_55[7:0]) +
	( 13'sd 4032) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32460) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25980) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13398) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20727) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13645) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27191) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26941) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24333) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20370) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14295) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27081) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2232) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6684) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1153) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32319) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24643) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28638) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18623) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28927) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2287) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1440) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1236) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31319) * $signed(input_fmap_81[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26058) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28379) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17935) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4745) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19975) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2352) * $signed(input_fmap_88[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6227) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28766) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24349) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24429) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25743) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8622) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9371) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13392) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15431) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14965) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22745) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5870) * $signed(input_fmap_103[7:0]) +
	( 11'sd 708) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29556) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21674) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1757) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7594) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31414) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32509) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31678) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25521) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6390) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23529) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8728) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17823) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27658) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10328) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24515) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20335) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31369) * $signed(input_fmap_123[7:0]) +
	( 2'sd 1) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23436) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19750) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19158) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2561) * $signed(input_fmap_128[7:0]) +
	( 13'sd 2277) * $signed(input_fmap_129[7:0]) +
	( 16'sd 28183) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24944) * $signed(input_fmap_131[7:0]) +
	( 11'sd 531) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28027) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24213) * $signed(input_fmap_134[7:0]) +
	( 16'sd 24836) * $signed(input_fmap_135[7:0]) +
	( 15'sd 14184) * $signed(input_fmap_136[7:0]) +
	( 16'sd 19889) * $signed(input_fmap_137[7:0]) +
	( 16'sd 20254) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3769) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30020) * $signed(input_fmap_140[7:0]) +
	( 16'sd 26537) * $signed(input_fmap_141[7:0]) +
	( 16'sd 18598) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10701) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28418) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25003) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1739) * $signed(input_fmap_146[7:0]) +
	( 12'sd 1481) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17402) * $signed(input_fmap_148[7:0]) +
	( 16'sd 21921) * $signed(input_fmap_149[7:0]) +
	( 16'sd 30997) * $signed(input_fmap_150[7:0]) +
	( 14'sd 5626) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24485) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14524) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4862) * $signed(input_fmap_154[7:0]) +
	( 15'sd 11328) * $signed(input_fmap_155[7:0]) +
	( 13'sd 3821) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23919) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25631) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27669) * $signed(input_fmap_159[7:0]) +
	( 15'sd 14585) * $signed(input_fmap_160[7:0]) +
	( 15'sd 13048) * $signed(input_fmap_161[7:0]) +
	( 14'sd 6496) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8923) * $signed(input_fmap_164[7:0]) +
	( 16'sd 16574) * $signed(input_fmap_165[7:0]) +
	( 16'sd 23044) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7178) * $signed(input_fmap_167[7:0]) +
	( 14'sd 7569) * $signed(input_fmap_168[7:0]) +
	( 14'sd 4496) * $signed(input_fmap_169[7:0]) +
	( 16'sd 19881) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12128) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15335) * $signed(input_fmap_172[7:0]) +
	( 15'sd 15728) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6094) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4222) * $signed(input_fmap_175[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1643) * $signed(input_fmap_177[7:0]) +
	( 16'sd 28236) * $signed(input_fmap_178[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_179[7:0]) +
	( 11'sd 600) * $signed(input_fmap_180[7:0]) +
	( 16'sd 19108) * $signed(input_fmap_181[7:0]) +
	( 6'sd 23) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17945) * $signed(input_fmap_183[7:0]) +
	( 16'sd 28754) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5167) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4910) * $signed(input_fmap_187[7:0]) +
	( 16'sd 19413) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17496) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_190[7:0]) +
	( 14'sd 7843) * $signed(input_fmap_191[7:0]) +
	( 15'sd 8666) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6877) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26900) * $signed(input_fmap_194[7:0]) +
	( 16'sd 21360) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6381) * $signed(input_fmap_196[7:0]) +
	( 13'sd 3341) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2978) * $signed(input_fmap_198[7:0]) +
	( 15'sd 11323) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18342) * $signed(input_fmap_200[7:0]) +
	( 16'sd 26377) * $signed(input_fmap_201[7:0]) +
	( 14'sd 4163) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25533) * $signed(input_fmap_203[7:0]) +
	( 16'sd 27623) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_205[7:0]) +
	( 16'sd 22597) * $signed(input_fmap_206[7:0]) +
	( 15'sd 15556) * $signed(input_fmap_207[7:0]) +
	( 13'sd 4018) * $signed(input_fmap_208[7:0]) +
	( 16'sd 25473) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4817) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15545) * $signed(input_fmap_211[7:0]) +
	( 15'sd 9431) * $signed(input_fmap_212[7:0]) +
	( 16'sd 31839) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30962) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7644) * $signed(input_fmap_215[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_216[7:0]) +
	( 15'sd 14034) * $signed(input_fmap_217[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20525) * $signed(input_fmap_219[7:0]) +
	( 15'sd 8940) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19384) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28051) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25353) * $signed(input_fmap_223[7:0]) +
	( 15'sd 11274) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1454) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6880) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9893) * $signed(input_fmap_227[7:0]) +
	( 16'sd 30336) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17483) * $signed(input_fmap_229[7:0]) +
	( 14'sd 5505) * $signed(input_fmap_230[7:0]) +
	( 15'sd 8563) * $signed(input_fmap_231[7:0]) +
	( 15'sd 10915) * $signed(input_fmap_232[7:0]) +
	( 13'sd 2937) * $signed(input_fmap_233[7:0]) +
	( 15'sd 12141) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21056) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10278) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10148) * $signed(input_fmap_237[7:0]) +
	( 14'sd 8108) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5491) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26877) * $signed(input_fmap_240[7:0]) +
	( 16'sd 24075) * $signed(input_fmap_241[7:0]) +
	( 16'sd 32759) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6388) * $signed(input_fmap_243[7:0]) +
	( 13'sd 3667) * $signed(input_fmap_244[7:0]) +
	( 12'sd 1873) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30605) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27846) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21619) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12447) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_250[7:0]) +
	( 16'sd 16520) * $signed(input_fmap_251[7:0]) +
	( 16'sd 18403) * $signed(input_fmap_252[7:0]) +
	( 16'sd 30491) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10239) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11785) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_133;
assign conv_mac_133 = 
	( 16'sd 16796) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10413) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28122) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2567) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31730) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3011) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1724) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28550) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24915) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28390) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26123) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22016) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19301) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2457) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7302) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31044) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28298) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19349) * $signed(input_fmap_19[7:0]) +
	( 10'sd 464) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9765) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21301) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13672) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5063) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32514) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28595) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11572) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25253) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21168) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25985) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28113) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17357) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6487) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15186) * $signed(input_fmap_37[7:0]) +
	( 10'sd 257) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28392) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13025) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32213) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19693) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29995) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19562) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26114) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3898) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6751) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22745) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16949) * $signed(input_fmap_50[7:0]) +
	( 11'sd 666) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23143) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5957) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22210) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15477) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19375) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1087) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9395) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19391) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27447) * $signed(input_fmap_64[7:0]) +
	( 14'sd 8097) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9060) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22404) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18170) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17444) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8222) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28387) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24600) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10866) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30767) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13547) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28024) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14576) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15943) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10304) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15038) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26759) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30784) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14491) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_87[7:0]) +
	( 14'sd 8044) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7847) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15949) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26246) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2928) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8195) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25222) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29292) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12376) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21880) * $signed(input_fmap_98[7:0]) +
	( 15'sd 14974) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32345) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4396) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19424) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28300) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18645) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1487) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8985) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16972) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27186) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9197) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13831) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20090) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2554) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24672) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5944) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30856) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15145) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31065) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5438) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32335) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12438) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10774) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3919) * $signed(input_fmap_126[7:0]) +
	( 11'sd 959) * $signed(input_fmap_127[7:0]) +
	( 14'sd 7005) * $signed(input_fmap_128[7:0]) +
	( 8'sd 118) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1825) * $signed(input_fmap_130[7:0]) +
	( 16'sd 27830) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5820) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31163) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31635) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32209) * $signed(input_fmap_135[7:0]) +
	( 16'sd 24373) * $signed(input_fmap_136[7:0]) +
	( 12'sd 1687) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11116) * $signed(input_fmap_138[7:0]) +
	( 16'sd 16512) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28085) * $signed(input_fmap_140[7:0]) +
	( 15'sd 15728) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30539) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12191) * $signed(input_fmap_143[7:0]) +
	( 16'sd 30297) * $signed(input_fmap_144[7:0]) +
	( 16'sd 20093) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7396) * $signed(input_fmap_146[7:0]) +
	( 16'sd 23175) * $signed(input_fmap_147[7:0]) +
	( 16'sd 18055) * $signed(input_fmap_148[7:0]) +
	( 15'sd 10687) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9848) * $signed(input_fmap_150[7:0]) +
	( 15'sd 9442) * $signed(input_fmap_151[7:0]) +
	( 15'sd 15607) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4963) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22370) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19919) * $signed(input_fmap_155[7:0]) +
	( 16'sd 16961) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30797) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11898) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3656) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18305) * $signed(input_fmap_160[7:0]) +
	( 14'sd 7441) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24427) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8316) * $signed(input_fmap_164[7:0]) +
	( 15'sd 8428) * $signed(input_fmap_165[7:0]) +
	( 15'sd 11506) * $signed(input_fmap_166[7:0]) +
	( 14'sd 4964) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14403) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10112) * $signed(input_fmap_169[7:0]) +
	( 14'sd 4275) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15785) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7579) * $signed(input_fmap_172[7:0]) +
	( 14'sd 8054) * $signed(input_fmap_173[7:0]) +
	( 14'sd 4228) * $signed(input_fmap_174[7:0]) +
	( 11'sd 555) * $signed(input_fmap_175[7:0]) +
	( 16'sd 19599) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24164) * $signed(input_fmap_177[7:0]) +
	( 16'sd 21024) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15806) * $signed(input_fmap_179[7:0]) +
	( 16'sd 18323) * $signed(input_fmap_180[7:0]) +
	( 16'sd 27563) * $signed(input_fmap_181[7:0]) +
	( 16'sd 32747) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12229) * $signed(input_fmap_183[7:0]) +
	( 13'sd 2624) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3097) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9248) * $signed(input_fmap_186[7:0]) +
	( 16'sd 20535) * $signed(input_fmap_187[7:0]) +
	( 6'sd 25) * $signed(input_fmap_188[7:0]) +
	( 13'sd 4048) * $signed(input_fmap_189[7:0]) +
	( 15'sd 14334) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31778) * $signed(input_fmap_191[7:0]) +
	( 16'sd 30953) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11316) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21394) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19105) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7937) * $signed(input_fmap_196[7:0]) +
	( 15'sd 13656) * $signed(input_fmap_197[7:0]) +
	( 15'sd 12949) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23732) * $signed(input_fmap_199[7:0]) +
	( 16'sd 16847) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6480) * $signed(input_fmap_201[7:0]) +
	( 16'sd 32370) * $signed(input_fmap_202[7:0]) +
	( 16'sd 31590) * $signed(input_fmap_203[7:0]) +
	( 16'sd 25834) * $signed(input_fmap_204[7:0]) +
	( 13'sd 4072) * $signed(input_fmap_205[7:0]) +
	( 15'sd 11793) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29222) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4576) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20150) * $signed(input_fmap_209[7:0]) +
	( 16'sd 32697) * $signed(input_fmap_210[7:0]) +
	( 16'sd 22269) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17929) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1147) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5116) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9599) * $signed(input_fmap_217[7:0]) +
	( 13'sd 2812) * $signed(input_fmap_218[7:0]) +
	( 14'sd 7316) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28147) * $signed(input_fmap_220[7:0]) +
	( 16'sd 30413) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3186) * $signed(input_fmap_222[7:0]) +
	( 16'sd 21336) * $signed(input_fmap_223[7:0]) +
	( 16'sd 26445) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2546) * $signed(input_fmap_225[7:0]) +
	( 16'sd 24718) * $signed(input_fmap_226[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31349) * $signed(input_fmap_228[7:0]) +
	( 14'sd 7518) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14822) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31633) * $signed(input_fmap_231[7:0]) +
	( 16'sd 30039) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18048) * $signed(input_fmap_233[7:0]) +
	( 16'sd 31775) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11467) * $signed(input_fmap_235[7:0]) +
	( 14'sd 4742) * $signed(input_fmap_236[7:0]) +
	( 15'sd 12167) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3866) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_239[7:0]) +
	( 16'sd 27097) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7825) * $signed(input_fmap_241[7:0]) +
	( 14'sd 4714) * $signed(input_fmap_242[7:0]) +
	( 11'sd 686) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12120) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12343) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14267) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8627) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4322) * $signed(input_fmap_248[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7115) * $signed(input_fmap_250[7:0]) +
	( 16'sd 29882) * $signed(input_fmap_251[7:0]) +
	( 13'sd 3653) * $signed(input_fmap_252[7:0]) +
	( 15'sd 14778) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13456) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11117) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_134;
assign conv_mac_134 = 
	( 16'sd 20746) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31301) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25181) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29185) * $signed(input_fmap_3[7:0]) +
	( 5'sd 12) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13616) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20585) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3396) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18078) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7314) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16584) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18315) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30375) * $signed(input_fmap_13[7:0]) +
	( 11'sd 1010) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21941) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14350) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27745) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26145) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17939) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8217) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9505) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17541) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17344) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12169) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20845) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13684) * $signed(input_fmap_26[7:0]) +
	( 13'sd 4015) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24298) * $signed(input_fmap_28[7:0]) +
	( 16'sd 29089) * $signed(input_fmap_29[7:0]) +
	( 14'sd 7558) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24708) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7059) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18887) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25568) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10521) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26698) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4580) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9638) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8932) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13156) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15802) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28280) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9906) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29653) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5433) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9356) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22156) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27257) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3637) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13878) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29579) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28806) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21613) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30469) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27903) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32334) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19207) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24917) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14353) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27559) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6915) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10789) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3106) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17941) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7125) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16699) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13340) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9107) * $signed(input_fmap_71[7:0]) +
	( 9'sd 225) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32118) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12538) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15906) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12496) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23255) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10803) * $signed(input_fmap_80[7:0]) +
	( 11'sd 633) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19765) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21782) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16654) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1576) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20734) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12574) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18669) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19291) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19748) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17257) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5269) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31931) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12909) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9303) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10312) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4566) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4741) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2835) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19049) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26532) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8793) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21615) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29676) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22314) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22825) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28371) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21653) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25483) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20542) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6236) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17950) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8193) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19441) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25517) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12873) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23825) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17634) * $signed(input_fmap_121[7:0]) +
	( 11'sd 695) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12258) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8816) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5016) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26763) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22494) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30637) * $signed(input_fmap_128[7:0]) +
	( 16'sd 30653) * $signed(input_fmap_129[7:0]) +
	( 15'sd 16297) * $signed(input_fmap_130[7:0]) +
	( 11'sd 781) * $signed(input_fmap_131[7:0]) +
	( 15'sd 15518) * $signed(input_fmap_132[7:0]) +
	( 13'sd 2693) * $signed(input_fmap_133[7:0]) +
	( 16'sd 30949) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20365) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7998) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9156) * $signed(input_fmap_137[7:0]) +
	( 16'sd 21441) * $signed(input_fmap_138[7:0]) +
	( 16'sd 29021) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24754) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13363) * $signed(input_fmap_141[7:0]) +
	( 12'sd 1126) * $signed(input_fmap_142[7:0]) +
	( 16'sd 19155) * $signed(input_fmap_143[7:0]) +
	( 15'sd 8335) * $signed(input_fmap_144[7:0]) +
	( 16'sd 19916) * $signed(input_fmap_145[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_146[7:0]) +
	( 16'sd 26424) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6320) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2163) * $signed(input_fmap_149[7:0]) +
	( 16'sd 28134) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3291) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6043) * $signed(input_fmap_152[7:0]) +
	( 14'sd 7433) * $signed(input_fmap_153[7:0]) +
	( 16'sd 21271) * $signed(input_fmap_154[7:0]) +
	( 15'sd 9917) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25358) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31657) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17240) * $signed(input_fmap_158[7:0]) +
	( 16'sd 29567) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26237) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20104) * $signed(input_fmap_161[7:0]) +
	( 16'sd 19144) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27005) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14009) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3463) * $signed(input_fmap_166[7:0]) +
	( 16'sd 19320) * $signed(input_fmap_167[7:0]) +
	( 16'sd 32158) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26359) * $signed(input_fmap_169[7:0]) +
	( 13'sd 3066) * $signed(input_fmap_170[7:0]) +
	( 15'sd 14543) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19546) * $signed(input_fmap_172[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_173[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_174[7:0]) +
	( 11'sd 987) * $signed(input_fmap_175[7:0]) +
	( 16'sd 32317) * $signed(input_fmap_176[7:0]) +
	( 15'sd 10665) * $signed(input_fmap_177[7:0]) +
	( 16'sd 19678) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20560) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15998) * $signed(input_fmap_180[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_181[7:0]) +
	( 11'sd 778) * $signed(input_fmap_182[7:0]) +
	( 14'sd 7073) * $signed(input_fmap_183[7:0]) +
	( 13'sd 3677) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7270) * $signed(input_fmap_185[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_186[7:0]) +
	( 15'sd 10289) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1582) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30812) * $signed(input_fmap_189[7:0]) +
	( 16'sd 26399) * $signed(input_fmap_190[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27091) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19384) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12430) * $signed(input_fmap_194[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_195[7:0]) +
	( 13'sd 2796) * $signed(input_fmap_196[7:0]) +
	( 15'sd 8434) * $signed(input_fmap_197[7:0]) +
	( 15'sd 12764) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28463) * $signed(input_fmap_199[7:0]) +
	( 14'sd 4927) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1604) * $signed(input_fmap_201[7:0]) +
	( 16'sd 29027) * $signed(input_fmap_202[7:0]) +
	( 16'sd 31173) * $signed(input_fmap_203[7:0]) +
	( 14'sd 7486) * $signed(input_fmap_204[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27649) * $signed(input_fmap_206[7:0]) +
	( 16'sd 27373) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25103) * $signed(input_fmap_208[7:0]) +
	( 16'sd 30201) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18840) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26759) * $signed(input_fmap_211[7:0]) +
	( 14'sd 6065) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1288) * $signed(input_fmap_213[7:0]) +
	( 16'sd 24840) * $signed(input_fmap_214[7:0]) +
	( 13'sd 3867) * $signed(input_fmap_215[7:0]) +
	( 13'sd 3549) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_217[7:0]) +
	( 16'sd 18649) * $signed(input_fmap_218[7:0]) +
	( 16'sd 27806) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4958) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15734) * $signed(input_fmap_221[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_222[7:0]) +
	( 15'sd 11034) * $signed(input_fmap_223[7:0]) +
	( 16'sd 23422) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1662) * $signed(input_fmap_225[7:0]) +
	( 15'sd 12892) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22785) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19798) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23777) * $signed(input_fmap_229[7:0]) +
	( 16'sd 26434) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24264) * $signed(input_fmap_231[7:0]) +
	( 16'sd 21985) * $signed(input_fmap_232[7:0]) +
	( 16'sd 31420) * $signed(input_fmap_233[7:0]) +
	( 15'sd 10755) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11140) * $signed(input_fmap_235[7:0]) +
	( 16'sd 32076) * $signed(input_fmap_236[7:0]) +
	( 14'sd 8064) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_238[7:0]) +
	( 10'sd 408) * $signed(input_fmap_239[7:0]) +
	( 15'sd 14755) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32641) * $signed(input_fmap_241[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_242[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_243[7:0]) +
	( 14'sd 4917) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19924) * $signed(input_fmap_245[7:0]) +
	( 13'sd 2260) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11571) * $signed(input_fmap_247[7:0]) +
	( 16'sd 28633) * $signed(input_fmap_248[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_249[7:0]) +
	( 16'sd 28894) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28940) * $signed(input_fmap_252[7:0]) +
	( 15'sd 16292) * $signed(input_fmap_253[7:0]) +
	( 16'sd 22425) * $signed(input_fmap_254[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_135;
assign conv_mac_135 = 
	( 13'sd 3419) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28081) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30242) * $signed(input_fmap_2[7:0]) +
	( 15'sd 11483) * $signed(input_fmap_3[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31216) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20874) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12609) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3350) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12568) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11631) * $signed(input_fmap_11[7:0]) +
	( 12'sd 2040) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12305) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32324) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10197) * $signed(input_fmap_15[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10869) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23130) * $signed(input_fmap_18[7:0]) +
	( 15'sd 16279) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5342) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19200) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15578) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14203) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26077) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1334) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26960) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5012) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3807) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13777) * $signed(input_fmap_31[7:0]) +
	( 10'sd 292) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21723) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19761) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32660) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7709) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17038) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27100) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6557) * $signed(input_fmap_40[7:0]) +
	( 16'sd 23417) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19810) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11640) * $signed(input_fmap_44[7:0]) +
	( 11'sd 648) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11521) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3463) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25414) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32066) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4578) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25750) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4112) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31267) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31603) * $signed(input_fmap_54[7:0]) +
	( 14'sd 8185) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2104) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32238) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25292) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18406) * $signed(input_fmap_59[7:0]) +
	( 11'sd 699) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13852) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24474) * $signed(input_fmap_62[7:0]) +
	( 11'sd 936) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11789) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25967) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17635) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11268) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10717) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1111) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17522) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20965) * $signed(input_fmap_71[7:0]) +
	( 11'sd 966) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21277) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17979) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30458) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16863) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21055) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8788) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9161) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23316) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2151) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25245) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25622) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7063) * $signed(input_fmap_85[7:0]) +
	( 14'sd 8171) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27219) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13050) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20872) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18719) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4540) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30454) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_93[7:0]) +
	( 12'sd 2045) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26853) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16323) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9290) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8969) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30482) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7201) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18174) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27517) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5278) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18906) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24647) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22524) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24488) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11887) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19715) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15915) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14590) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6276) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11365) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32030) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19357) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2599) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13577) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10758) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12519) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3835) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32594) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2695) * $signed(input_fmap_124[7:0]) +
	( 14'sd 8045) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18157) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28940) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30257) * $signed(input_fmap_128[7:0]) +
	( 16'sd 20414) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27569) * $signed(input_fmap_130[7:0]) +
	( 16'sd 21216) * $signed(input_fmap_131[7:0]) +
	( 16'sd 29038) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16487) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_134[7:0]) +
	( 14'sd 7900) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_136[7:0]) +
	( 16'sd 31761) * $signed(input_fmap_137[7:0]) +
	( 15'sd 13623) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3205) * $signed(input_fmap_139[7:0]) +
	( 16'sd 31543) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20090) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19652) * $signed(input_fmap_142[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6221) * $signed(input_fmap_144[7:0]) +
	( 11'sd 977) * $signed(input_fmap_145[7:0]) +
	( 14'sd 6373) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3215) * $signed(input_fmap_147[7:0]) +
	( 11'sd 582) * $signed(input_fmap_148[7:0]) +
	( 11'sd 713) * $signed(input_fmap_149[7:0]) +
	( 15'sd 11487) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14956) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14446) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14877) * $signed(input_fmap_153[7:0]) +
	( 16'sd 21847) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10003) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24588) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14016) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20212) * $signed(input_fmap_158[7:0]) +
	( 16'sd 30890) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17138) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20347) * $signed(input_fmap_161[7:0]) +
	( 15'sd 15338) * $signed(input_fmap_162[7:0]) +
	( 16'sd 17309) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3043) * $signed(input_fmap_164[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_165[7:0]) +
	( 10'sd 371) * $signed(input_fmap_166[7:0]) +
	( 16'sd 27997) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5045) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3384) * $signed(input_fmap_169[7:0]) +
	( 15'sd 15225) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3538) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3279) * $signed(input_fmap_172[7:0]) +
	( 16'sd 22047) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10623) * $signed(input_fmap_174[7:0]) +
	( 15'sd 14428) * $signed(input_fmap_175[7:0]) +
	( 11'sd 932) * $signed(input_fmap_176[7:0]) +
	( 15'sd 13748) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10463) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3183) * $signed(input_fmap_180[7:0]) +
	( 16'sd 32731) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5069) * $signed(input_fmap_182[7:0]) +
	( 15'sd 8677) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13356) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27382) * $signed(input_fmap_185[7:0]) +
	( 16'sd 29435) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25633) * $signed(input_fmap_187[7:0]) +
	( 16'sd 19981) * $signed(input_fmap_188[7:0]) +
	( 15'sd 13440) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27602) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31845) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27901) * $signed(input_fmap_192[7:0]) +
	( 12'sd 1870) * $signed(input_fmap_193[7:0]) +
	( 16'sd 22675) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19643) * $signed(input_fmap_195[7:0]) +
	( 16'sd 27180) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22958) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12588) * $signed(input_fmap_199[7:0]) +
	( 16'sd 23338) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15143) * $signed(input_fmap_201[7:0]) +
	( 13'sd 3398) * $signed(input_fmap_202[7:0]) +
	( 15'sd 11634) * $signed(input_fmap_203[7:0]) +
	( 16'sd 18433) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12454) * $signed(input_fmap_205[7:0]) +
	( 15'sd 14820) * $signed(input_fmap_206[7:0]) +
	( 11'sd 740) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18035) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23486) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10097) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3584) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11734) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30826) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1245) * $signed(input_fmap_215[7:0]) +
	( 16'sd 21866) * $signed(input_fmap_216[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_217[7:0]) +
	( 14'sd 8096) * $signed(input_fmap_218[7:0]) +
	( 16'sd 23459) * $signed(input_fmap_219[7:0]) +
	( 13'sd 3959) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23239) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2487) * $signed(input_fmap_222[7:0]) +
	( 11'sd 941) * $signed(input_fmap_223[7:0]) +
	( 16'sd 21276) * $signed(input_fmap_224[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_225[7:0]) +
	( 15'sd 12711) * $signed(input_fmap_226[7:0]) +
	( 15'sd 8996) * $signed(input_fmap_227[7:0]) +
	( 15'sd 15417) * $signed(input_fmap_228[7:0]) +
	( 16'sd 30365) * $signed(input_fmap_229[7:0]) +
	( 14'sd 5801) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_231[7:0]) +
	( 15'sd 10482) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1550) * $signed(input_fmap_233[7:0]) +
	( 16'sd 28585) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29254) * $signed(input_fmap_235[7:0]) +
	( 16'sd 17205) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6205) * $signed(input_fmap_237[7:0]) +
	( 16'sd 25332) * $signed(input_fmap_238[7:0]) +
	( 16'sd 24114) * $signed(input_fmap_239[7:0]) +
	( 16'sd 24320) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20066) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26722) * $signed(input_fmap_242[7:0]) +
	( 15'sd 16001) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7731) * $signed(input_fmap_245[7:0]) +
	( 16'sd 24475) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18808) * $signed(input_fmap_247[7:0]) +
	( 14'sd 8122) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14790) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32057) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27980) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10768) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24211) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9289) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24348) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_136;
assign conv_mac_136 = 
	( 13'sd 3383) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16694) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10847) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15976) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18842) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7370) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4587) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29029) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1168) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4596) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24541) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6148) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7100) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1307) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24837) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9343) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13476) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32360) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22314) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18711) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10791) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27406) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10449) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19608) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6205) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28459) * $signed(input_fmap_27[7:0]) +
	( 10'sd 483) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26995) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31365) * $signed(input_fmap_31[7:0]) +
	( 11'sd 819) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13233) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25791) * $signed(input_fmap_34[7:0]) +
	( 14'sd 4384) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18781) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29962) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7455) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30103) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29338) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7462) * $signed(input_fmap_41[7:0]) +
	( 14'sd 8099) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23351) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29535) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30641) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18334) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8968) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11386) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28850) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11402) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28576) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9768) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31459) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22561) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19362) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25957) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29472) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30778) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7258) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3002) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15641) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30086) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3952) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16501) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29268) * $signed(input_fmap_70[7:0]) +
	( 7'sd 46) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28574) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6565) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10625) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27156) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15782) * $signed(input_fmap_76[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_77[7:0]) +
	( 11'sd 996) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30996) * $signed(input_fmap_79[7:0]) +
	( 11'sd 737) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17538) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21201) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20924) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30956) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4735) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9743) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10004) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24680) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3557) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7996) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27575) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28612) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21476) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17021) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7081) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27924) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13867) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23211) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26002) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4493) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29301) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4862) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9811) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10663) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31812) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8895) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5331) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20696) * $signed(input_fmap_112[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11785) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15594) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32663) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10860) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1747) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27907) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4505) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17190) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2774) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12389) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23898) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23994) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31385) * $signed(input_fmap_128[7:0]) +
	( 14'sd 6723) * $signed(input_fmap_129[7:0]) +
	( 15'sd 9953) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15932) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11205) * $signed(input_fmap_132[7:0]) +
	( 16'sd 19668) * $signed(input_fmap_133[7:0]) +
	( 15'sd 13494) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21349) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_136[7:0]) +
	( 16'sd 30376) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19666) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24415) * $signed(input_fmap_139[7:0]) +
	( 16'sd 21609) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10121) * $signed(input_fmap_141[7:0]) +
	( 15'sd 13825) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12516) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_144[7:0]) +
	( 16'sd 29145) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18646) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29108) * $signed(input_fmap_147[7:0]) +
	( 15'sd 13997) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23920) * $signed(input_fmap_149[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12525) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22465) * $signed(input_fmap_152[7:0]) +
	( 16'sd 20923) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25046) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12800) * $signed(input_fmap_155[7:0]) +
	( 12'sd 1789) * $signed(input_fmap_156[7:0]) +
	( 14'sd 4519) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26275) * $signed(input_fmap_159[7:0]) +
	( 15'sd 13504) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1628) * $signed(input_fmap_161[7:0]) +
	( 15'sd 9238) * $signed(input_fmap_162[7:0]) +
	( 16'sd 21644) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24469) * $signed(input_fmap_164[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_165[7:0]) +
	( 16'sd 16871) * $signed(input_fmap_166[7:0]) +
	( 15'sd 15624) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5873) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30275) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18498) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11870) * $signed(input_fmap_171[7:0]) +
	( 16'sd 24797) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23688) * $signed(input_fmap_173[7:0]) +
	( 16'sd 21482) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5741) * $signed(input_fmap_175[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5651) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2739) * $signed(input_fmap_178[7:0]) +
	( 15'sd 9373) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26394) * $signed(input_fmap_180[7:0]) +
	( 14'sd 4581) * $signed(input_fmap_181[7:0]) +
	( 16'sd 28077) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29252) * $signed(input_fmap_183[7:0]) +
	( 11'sd 745) * $signed(input_fmap_184[7:0]) +
	( 16'sd 31940) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3534) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2215) * $signed(input_fmap_187[7:0]) +
	( 13'sd 3664) * $signed(input_fmap_188[7:0]) +
	( 15'sd 14904) * $signed(input_fmap_189[7:0]) +
	( 8'sd 107) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29664) * $signed(input_fmap_191[7:0]) +
	( 16'sd 17222) * $signed(input_fmap_192[7:0]) +
	( 15'sd 13704) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30255) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24176) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22292) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22643) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29123) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29224) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15734) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3842) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8808) * $signed(input_fmap_202[7:0]) +
	( 13'sd 3839) * $signed(input_fmap_203[7:0]) +
	( 11'sd 712) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18431) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6845) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_207[7:0]) +
	( 16'sd 27766) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1660) * $signed(input_fmap_210[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19833) * $signed(input_fmap_212[7:0]) +
	( 15'sd 8455) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15196) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5078) * $signed(input_fmap_215[7:0]) +
	( 16'sd 26703) * $signed(input_fmap_216[7:0]) +
	( 15'sd 15218) * $signed(input_fmap_217[7:0]) +
	( 15'sd 12907) * $signed(input_fmap_218[7:0]) +
	( 16'sd 27719) * $signed(input_fmap_219[7:0]) +
	( 14'sd 6570) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6752) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3626) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17688) * $signed(input_fmap_223[7:0]) +
	( 16'sd 32532) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32280) * $signed(input_fmap_226[7:0]) +
	( 16'sd 25126) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24766) * $signed(input_fmap_228[7:0]) +
	( 16'sd 28857) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24147) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12713) * $signed(input_fmap_232[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_233[7:0]) +
	( 15'sd 12579) * $signed(input_fmap_234[7:0]) +
	( 11'sd 748) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30792) * $signed(input_fmap_236[7:0]) +
	( 15'sd 15631) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5375) * $signed(input_fmap_238[7:0]) +
	( 16'sd 24393) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22199) * $signed(input_fmap_240[7:0]) +
	( 16'sd 28297) * $signed(input_fmap_241[7:0]) +
	( 14'sd 4875) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13961) * $signed(input_fmap_243[7:0]) +
	( 16'sd 16537) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5243) * $signed(input_fmap_245[7:0]) +
	( 16'sd 32305) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18245) * $signed(input_fmap_247[7:0]) +
	( 15'sd 9100) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_249[7:0]) +
	( 13'sd 2430) * $signed(input_fmap_250[7:0]) +
	( 16'sd 16454) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4819) * $signed(input_fmap_252[7:0]) +
	( 16'sd 21804) * $signed(input_fmap_253[7:0]) +
	( 16'sd 30252) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14794) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_137;
assign conv_mac_137 = 
	( 16'sd 18917) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9563) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11027) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26713) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12739) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21224) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6872) * $signed(input_fmap_6[7:0]) +
	( 10'sd 290) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6679) * $signed(input_fmap_8[7:0]) +
	( 16'sd 32362) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12889) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14431) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12509) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9722) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6359) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26931) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7581) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28854) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6774) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7612) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17026) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28967) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29008) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2212) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10909) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30915) * $signed(input_fmap_26[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1059) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21089) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9585) * $signed(input_fmap_30[7:0]) +
	( 15'sd 16002) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28251) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2334) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18661) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21418) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2550) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4766) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16890) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21101) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24138) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32411) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1646) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2961) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7872) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30785) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24614) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21776) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23497) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24604) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5898) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6221) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17549) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3038) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20759) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29362) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14817) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10531) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7381) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12682) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15517) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27549) * $signed(input_fmap_64[7:0]) +
	( 10'sd 332) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10887) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7564) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3558) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18494) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26705) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2138) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24428) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11507) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24362) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32703) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25299) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28416) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19735) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4887) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22688) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31251) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29899) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21403) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11146) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24741) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12010) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26432) * $signed(input_fmap_88[7:0]) +
	( 7'sd 48) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15758) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28739) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8562) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22756) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16260) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27161) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27391) * $signed(input_fmap_96[7:0]) +
	( 15'sd 16031) * $signed(input_fmap_97[7:0]) +
	( 11'sd 670) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15611) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15502) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1802) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17049) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7857) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31136) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29229) * $signed(input_fmap_105[7:0]) +
	( 11'sd 604) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7205) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32341) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3957) * $signed(input_fmap_109[7:0]) +
	( 10'sd 470) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31793) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21228) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29704) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26214) * $signed(input_fmap_114[7:0]) +
	( 16'sd 32680) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1401) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17506) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1203) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16396) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20300) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11095) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30477) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24097) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25773) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4228) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17685) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13941) * $signed(input_fmap_128[7:0]) +
	( 16'sd 23561) * $signed(input_fmap_129[7:0]) +
	( 10'sd 335) * $signed(input_fmap_130[7:0]) +
	( 15'sd 11590) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1109) * $signed(input_fmap_132[7:0]) +
	( 15'sd 8553) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25206) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21555) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_136[7:0]) +
	( 16'sd 32443) * $signed(input_fmap_137[7:0]) +
	( 16'sd 21069) * $signed(input_fmap_138[7:0]) +
	( 14'sd 7206) * $signed(input_fmap_139[7:0]) +
	( 16'sd 32763) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5559) * $signed(input_fmap_141[7:0]) +
	( 14'sd 4141) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26399) * $signed(input_fmap_143[7:0]) +
	( 14'sd 6559) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23339) * $signed(input_fmap_145[7:0]) +
	( 15'sd 11007) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30020) * $signed(input_fmap_147[7:0]) +
	( 15'sd 12169) * $signed(input_fmap_148[7:0]) +
	( 16'sd 22231) * $signed(input_fmap_149[7:0]) +
	( 16'sd 26920) * $signed(input_fmap_150[7:0]) +
	( 15'sd 13215) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23162) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25191) * $signed(input_fmap_153[7:0]) +
	( 16'sd 21699) * $signed(input_fmap_154[7:0]) +
	( 16'sd 29118) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18971) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13193) * $signed(input_fmap_157[7:0]) +
	( 16'sd 22586) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12079) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21907) * $signed(input_fmap_160[7:0]) +
	( 14'sd 7040) * $signed(input_fmap_161[7:0]) +
	( 14'sd 5450) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30054) * $signed(input_fmap_163[7:0]) +
	( 16'sd 30427) * $signed(input_fmap_164[7:0]) +
	( 15'sd 13325) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2528) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17718) * $signed(input_fmap_167[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_168[7:0]) +
	( 15'sd 15228) * $signed(input_fmap_169[7:0]) +
	( 16'sd 26051) * $signed(input_fmap_170[7:0]) +
	( 14'sd 4277) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_172[7:0]) +
	( 16'sd 26675) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19519) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25343) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3045) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19995) * $signed(input_fmap_177[7:0]) +
	( 16'sd 23671) * $signed(input_fmap_178[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6905) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3187) * $signed(input_fmap_181[7:0]) +
	( 16'sd 20141) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2348) * $signed(input_fmap_183[7:0]) +
	( 16'sd 25100) * $signed(input_fmap_184[7:0]) +
	( 16'sd 23454) * $signed(input_fmap_185[7:0]) +
	( 15'sd 11511) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22494) * $signed(input_fmap_187[7:0]) +
	( 14'sd 6720) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17597) * $signed(input_fmap_189[7:0]) +
	( 16'sd 16984) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19459) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14439) * $signed(input_fmap_192[7:0]) +
	( 14'sd 4585) * $signed(input_fmap_193[7:0]) +
	( 16'sd 25003) * $signed(input_fmap_194[7:0]) +
	( 16'sd 30870) * $signed(input_fmap_195[7:0]) +
	( 16'sd 18093) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5854) * $signed(input_fmap_197[7:0]) +
	( 16'sd 32278) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5826) * $signed(input_fmap_199[7:0]) +
	( 16'sd 30233) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18840) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8766) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30019) * $signed(input_fmap_203[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_204[7:0]) +
	( 16'sd 16635) * $signed(input_fmap_205[7:0]) +
	( 10'sd 508) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5736) * $signed(input_fmap_207[7:0]) +
	( 16'sd 27024) * $signed(input_fmap_208[7:0]) +
	( 15'sd 12806) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4649) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30593) * $signed(input_fmap_211[7:0]) +
	( 16'sd 32004) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_213[7:0]) +
	( 13'sd 3216) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29829) * $signed(input_fmap_215[7:0]) +
	( 10'sd 376) * $signed(input_fmap_216[7:0]) +
	( 12'sd 1615) * $signed(input_fmap_217[7:0]) +
	( 13'sd 2058) * $signed(input_fmap_218[7:0]) +
	( 12'sd 1631) * $signed(input_fmap_219[7:0]) +
	( 15'sd 16278) * $signed(input_fmap_220[7:0]) +
	( 13'sd 2191) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19092) * $signed(input_fmap_222[7:0]) +
	( 16'sd 18128) * $signed(input_fmap_223[7:0]) +
	( 15'sd 16019) * $signed(input_fmap_224[7:0]) +
	( 14'sd 8116) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18549) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5767) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_228[7:0]) +
	( 16'sd 31090) * $signed(input_fmap_229[7:0]) +
	( 16'sd 16738) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1413) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18331) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14764) * $signed(input_fmap_233[7:0]) +
	( 15'sd 11940) * $signed(input_fmap_234[7:0]) +
	( 15'sd 9182) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31656) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10127) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3260) * $signed(input_fmap_238[7:0]) +
	( 12'sd 1682) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23635) * $signed(input_fmap_240[7:0]) +
	( 15'sd 14415) * $signed(input_fmap_241[7:0]) +
	( 15'sd 9504) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10173) * $signed(input_fmap_243[7:0]) +
	( 15'sd 14849) * $signed(input_fmap_244[7:0]) +
	( 16'sd 16872) * $signed(input_fmap_245[7:0]) +
	( 16'sd 26923) * $signed(input_fmap_246[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_247[7:0]) +
	( 15'sd 12243) * $signed(input_fmap_248[7:0]) +
	( 11'sd 636) * $signed(input_fmap_249[7:0]) +
	( 12'sd 1482) * $signed(input_fmap_250[7:0]) +
	( 10'sd 352) * $signed(input_fmap_251[7:0]) +
	( 11'sd 620) * $signed(input_fmap_252[7:0]) +
	( 16'sd 18241) * $signed(input_fmap_253[7:0]) +
	( 16'sd 27176) * $signed(input_fmap_254[7:0]) +
	( 16'sd 16389) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_138;
assign conv_mac_138 = 
	( 15'sd 14769) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4567) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21093) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27614) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9071) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22155) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19195) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11591) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27311) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14380) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26741) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27800) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31831) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32081) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27843) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26606) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29176) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10485) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32000) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7179) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10974) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_24[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14365) * $signed(input_fmap_26[7:0]) +
	( 10'sd 352) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16670) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10368) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9629) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28324) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9405) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13276) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19845) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19434) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8442) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32342) * $signed(input_fmap_39[7:0]) +
	( 10'sd 312) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21981) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11124) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10095) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16905) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26295) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9471) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3888) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4983) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25240) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2980) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5956) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26985) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8892) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24982) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10916) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29236) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22966) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22905) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18302) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18837) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31782) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31801) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11730) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18402) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28631) * $signed(input_fmap_72[7:0]) +
	( 11'sd 1009) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15413) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5948) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13890) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12907) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13392) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29349) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10574) * $signed(input_fmap_81[7:0]) +
	( 15'sd 10004) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10154) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28587) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20550) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1252) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19458) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8308) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10689) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19018) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24227) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18812) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27611) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30896) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12099) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1027) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24665) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32043) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11370) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8267) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11268) * $signed(input_fmap_102[7:0]) +
	( 8'sd 70) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1541) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6322) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25956) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20843) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20967) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16254) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5954) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21171) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4438) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28116) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1505) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20762) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13374) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15999) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23548) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22498) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9616) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14244) * $signed(input_fmap_122[7:0]) +
	( 10'sd 500) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20280) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22414) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12577) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15503) * $signed(input_fmap_128[7:0]) +
	( 15'sd 12064) * $signed(input_fmap_129[7:0]) +
	( 15'sd 9645) * $signed(input_fmap_130[7:0]) +
	( 16'sd 26099) * $signed(input_fmap_131[7:0]) +
	( 16'sd 28554) * $signed(input_fmap_132[7:0]) +
	( 12'sd 1503) * $signed(input_fmap_133[7:0]) +
	( 16'sd 30431) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27368) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7407) * $signed(input_fmap_136[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_137[7:0]) +
	( 15'sd 12706) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8575) * $signed(input_fmap_139[7:0]) +
	( 14'sd 4400) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10305) * $signed(input_fmap_141[7:0]) +
	( 11'sd 779) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10900) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9881) * $signed(input_fmap_144[7:0]) +
	( 15'sd 12492) * $signed(input_fmap_145[7:0]) +
	( 16'sd 25648) * $signed(input_fmap_146[7:0]) +
	( 14'sd 7596) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23321) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12140) * $signed(input_fmap_149[7:0]) +
	( 16'sd 32738) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3784) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23993) * $signed(input_fmap_154[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_155[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23028) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9306) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12446) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27730) * $signed(input_fmap_160[7:0]) +
	( 16'sd 29481) * $signed(input_fmap_161[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8619) * $signed(input_fmap_163[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10703) * $signed(input_fmap_165[7:0]) +
	( 16'sd 32205) * $signed(input_fmap_166[7:0]) +
	( 10'sd 486) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17459) * $signed(input_fmap_168[7:0]) +
	( 14'sd 4614) * $signed(input_fmap_169[7:0]) +
	( 14'sd 6767) * $signed(input_fmap_170[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_171[7:0]) +
	( 16'sd 24915) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29130) * $signed(input_fmap_173[7:0]) +
	( 11'sd 961) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15577) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27331) * $signed(input_fmap_176[7:0]) +
	( 15'sd 10639) * $signed(input_fmap_177[7:0]) +
	( 16'sd 28190) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2707) * $signed(input_fmap_179[7:0]) +
	( 13'sd 2181) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11816) * $signed(input_fmap_181[7:0]) +
	( 15'sd 11223) * $signed(input_fmap_182[7:0]) +
	( 14'sd 7128) * $signed(input_fmap_183[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26724) * $signed(input_fmap_185[7:0]) +
	( 16'sd 29935) * $signed(input_fmap_186[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_187[7:0]) +
	( 15'sd 9313) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3116) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28902) * $signed(input_fmap_190[7:0]) +
	( 16'sd 25236) * $signed(input_fmap_191[7:0]) +
	( 12'sd 1916) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30084) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21162) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25779) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19471) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22304) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31903) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_201[7:0]) +
	( 13'sd 3961) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19996) * $signed(input_fmap_203[7:0]) +
	( 16'sd 29727) * $signed(input_fmap_204[7:0]) +
	( 16'sd 21582) * $signed(input_fmap_205[7:0]) +
	( 15'sd 10630) * $signed(input_fmap_206[7:0]) +
	( 14'sd 6352) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17655) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24056) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31134) * $signed(input_fmap_210[7:0]) +
	( 15'sd 13587) * $signed(input_fmap_211[7:0]) +
	( 15'sd 9344) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1803) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18167) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_216[7:0]) +
	( 15'sd 15307) * $signed(input_fmap_217[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_218[7:0]) +
	( 16'sd 27669) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26151) * $signed(input_fmap_220[7:0]) +
	( 16'sd 24489) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5874) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24631) * $signed(input_fmap_223[7:0]) +
	( 16'sd 18036) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3707) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11591) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24281) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19387) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24977) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18737) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3045) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9240) * $signed(input_fmap_232[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_233[7:0]) +
	( 13'sd 2300) * $signed(input_fmap_234[7:0]) +
	( 16'sd 18468) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10800) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17839) * $signed(input_fmap_238[7:0]) +
	( 16'sd 29131) * $signed(input_fmap_239[7:0]) +
	( 14'sd 7224) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21142) * $signed(input_fmap_241[7:0]) +
	( 16'sd 25385) * $signed(input_fmap_242[7:0]) +
	( 16'sd 21468) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1171) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20041) * $signed(input_fmap_246[7:0]) +
	( 12'sd 1754) * $signed(input_fmap_247[7:0]) +
	( 11'sd 880) * $signed(input_fmap_248[7:0]) +
	( 16'sd 16503) * $signed(input_fmap_249[7:0]) +
	( 14'sd 5197) * $signed(input_fmap_250[7:0]) +
	( 16'sd 30267) * $signed(input_fmap_251[7:0]) +
	( 16'sd 32362) * $signed(input_fmap_252[7:0]) +
	( 16'sd 21389) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5612) * $signed(input_fmap_254[7:0]) +
	( 14'sd 7192) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_139;
assign conv_mac_139 = 
	( 16'sd 30938) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25566) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2512) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9302) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30173) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3252) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14975) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27503) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17893) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23296) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27009) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4380) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3103) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12541) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10082) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31538) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29012) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7829) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30521) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30783) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22520) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31689) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15531) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17116) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19537) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6073) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24804) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25421) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5714) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6171) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9431) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5436) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21391) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12472) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22483) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7436) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28384) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24867) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31726) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8374) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6022) * $signed(input_fmap_45[7:0]) +
	( 16'sd 20685) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22118) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10608) * $signed(input_fmap_48[7:0]) +
	( 16'sd 25009) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9696) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24628) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23383) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1112) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19702) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18412) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14652) * $signed(input_fmap_56[7:0]) +
	( 16'sd 26372) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13688) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21386) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32239) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17772) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11347) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29692) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21844) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3741) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26390) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21649) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15143) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3160) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25698) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30993) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20164) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22272) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1302) * $signed(input_fmap_75[7:0]) +
	( 11'sd 703) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21989) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9893) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2293) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13743) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26452) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2303) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31367) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30191) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7367) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32079) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10796) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16227) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24052) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26612) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8547) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6788) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9084) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21196) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14828) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17894) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2551) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31412) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8393) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17150) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9331) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7536) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2183) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13125) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10328) * $signed(input_fmap_109[7:0]) +
	( 14'sd 8001) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30005) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16566) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24191) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31455) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10287) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20923) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26688) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6929) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20352) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32543) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9753) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8609) * $signed(input_fmap_123[7:0]) +
	( 11'sd 947) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21030) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2842) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5984) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4323) * $signed(input_fmap_128[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_129[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24808) * $signed(input_fmap_131[7:0]) +
	( 10'sd 497) * $signed(input_fmap_132[7:0]) +
	( 16'sd 30819) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24718) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21446) * $signed(input_fmap_135[7:0]) +
	( 16'sd 16818) * $signed(input_fmap_136[7:0]) +
	( 16'sd 31801) * $signed(input_fmap_137[7:0]) +
	( 16'sd 18786) * $signed(input_fmap_138[7:0]) +
	( 16'sd 29432) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10467) * $signed(input_fmap_141[7:0]) +
	( 16'sd 18018) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17914) * $signed(input_fmap_143[7:0]) +
	( 16'sd 16588) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27509) * $signed(input_fmap_145[7:0]) +
	( 13'sd 2687) * $signed(input_fmap_146[7:0]) +
	( 16'sd 28343) * $signed(input_fmap_147[7:0]) +
	( 16'sd 24142) * $signed(input_fmap_148[7:0]) +
	( 12'sd 1235) * $signed(input_fmap_149[7:0]) +
	( 12'sd 2020) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4543) * $signed(input_fmap_151[7:0]) +
	( 16'sd 25780) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3921) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11604) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12311) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7828) * $signed(input_fmap_156[7:0]) +
	( 13'sd 2984) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28216) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6020) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_160[7:0]) +
	( 16'sd 24520) * $signed(input_fmap_161[7:0]) +
	( 13'sd 3078) * $signed(input_fmap_162[7:0]) +
	( 14'sd 8029) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10643) * $signed(input_fmap_164[7:0]) +
	( 13'sd 3095) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9041) * $signed(input_fmap_166[7:0]) +
	( 16'sd 21330) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20828) * $signed(input_fmap_168[7:0]) +
	( 16'sd 31779) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5329) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19399) * $signed(input_fmap_171[7:0]) +
	( 16'sd 18222) * $signed(input_fmap_172[7:0]) +
	( 15'sd 9341) * $signed(input_fmap_173[7:0]) +
	( 16'sd 25606) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21893) * $signed(input_fmap_175[7:0]) +
	( 16'sd 24737) * $signed(input_fmap_176[7:0]) +
	( 16'sd 20990) * $signed(input_fmap_177[7:0]) +
	( 16'sd 28618) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25728) * $signed(input_fmap_179[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_180[7:0]) +
	( 15'sd 13073) * $signed(input_fmap_181[7:0]) +
	( 16'sd 31304) * $signed(input_fmap_182[7:0]) +
	( 16'sd 16837) * $signed(input_fmap_183[7:0]) +
	( 16'sd 18546) * $signed(input_fmap_184[7:0]) +
	( 15'sd 9650) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26081) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25128) * $signed(input_fmap_187[7:0]) +
	( 14'sd 7663) * $signed(input_fmap_188[7:0]) +
	( 16'sd 22513) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13459) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20240) * $signed(input_fmap_191[7:0]) +
	( 16'sd 18984) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11284) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27163) * $signed(input_fmap_194[7:0]) +
	( 16'sd 18257) * $signed(input_fmap_195[7:0]) +
	( 16'sd 18019) * $signed(input_fmap_196[7:0]) +
	( 16'sd 16882) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29954) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14663) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26527) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_201[7:0]) +
	( 11'sd 838) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13072) * $signed(input_fmap_203[7:0]) +
	( 16'sd 23092) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6618) * $signed(input_fmap_205[7:0]) +
	( 16'sd 22723) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1143) * $signed(input_fmap_207[7:0]) +
	( 8'sd 82) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26760) * $signed(input_fmap_209[7:0]) +
	( 16'sd 26217) * $signed(input_fmap_210[7:0]) +
	( 10'sd 342) * $signed(input_fmap_211[7:0]) +
	( 16'sd 20873) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5435) * $signed(input_fmap_213[7:0]) +
	( 16'sd 24874) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1114) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28936) * $signed(input_fmap_216[7:0]) +
	( 13'sd 3392) * $signed(input_fmap_217[7:0]) +
	( 15'sd 14062) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10222) * $signed(input_fmap_219[7:0]) +
	( 10'sd 412) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25346) * $signed(input_fmap_221[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12651) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7365) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5091) * $signed(input_fmap_225[7:0]) +
	( 14'sd 4207) * $signed(input_fmap_226[7:0]) +
	( 16'sd 23509) * $signed(input_fmap_227[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_228[7:0]) +
	( 12'sd 1102) * $signed(input_fmap_229[7:0]) +
	( 13'sd 2782) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24820) * $signed(input_fmap_231[7:0]) +
	( 16'sd 27643) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11124) * $signed(input_fmap_233[7:0]) +
	( 16'sd 16811) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5231) * $signed(input_fmap_235[7:0]) +
	( 16'sd 19255) * $signed(input_fmap_236[7:0]) +
	( 16'sd 18289) * $signed(input_fmap_237[7:0]) +
	( 14'sd 4977) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23206) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19594) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_241[7:0]) +
	( 16'sd 18095) * $signed(input_fmap_242[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_243[7:0]) +
	( 15'sd 9879) * $signed(input_fmap_244[7:0]) +
	( 9'sd 138) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11982) * $signed(input_fmap_246[7:0]) +
	( 13'sd 2982) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26652) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17305) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22436) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22121) * $signed(input_fmap_251[7:0]) +
	( 16'sd 19747) * $signed(input_fmap_252[7:0]) +
	( 14'sd 4166) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5568) * $signed(input_fmap_254[7:0]) +
	( 15'sd 13360) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_140;
assign conv_mac_140 = 
	( 15'sd 13079) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25804) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20806) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1032) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8660) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13607) * $signed(input_fmap_6[7:0]) +
	( 11'sd 979) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29742) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23403) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30173) * $signed(input_fmap_10[7:0]) +
	( 13'sd 4042) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29197) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8689) * $signed(input_fmap_13[7:0]) +
	( 11'sd 746) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1812) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12979) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6440) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23658) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10853) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_20[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27477) * $signed(input_fmap_22[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24991) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31118) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29177) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9498) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21540) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2244) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15482) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2287) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3227) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19904) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28097) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27183) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5402) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2756) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31715) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11666) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16440) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26696) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19634) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21554) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18658) * $signed(input_fmap_46[7:0]) +
	( 12'sd 1929) * $signed(input_fmap_47[7:0]) +
	( 16'sd 23512) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24673) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28072) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31041) * $signed(input_fmap_51[7:0]) +
	( 14'sd 8031) * $signed(input_fmap_52[7:0]) +
	( 11'sd 986) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5016) * $signed(input_fmap_54[7:0]) +
	( 12'sd 2008) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29389) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12597) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13338) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16739) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1739) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25471) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22648) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11711) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14672) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11963) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12014) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32355) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25430) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10847) * $signed(input_fmap_70[7:0]) +
	( 11'sd 631) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26857) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8910) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7270) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22272) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19377) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11841) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13141) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16217) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26475) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13681) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18213) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16768) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17892) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28014) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21343) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30343) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9492) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15180) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21065) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2317) * $signed(input_fmap_93[7:0]) +
	( 11'sd 872) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16084) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14812) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9348) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4253) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28310) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4889) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9072) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7311) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27583) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25926) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18986) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24595) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_108[7:0]) +
	( 10'sd 319) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18419) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1358) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28896) * $signed(input_fmap_113[7:0]) +
	( 15'sd 10939) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18027) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5700) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6675) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7514) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27032) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21033) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19673) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10144) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29765) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24017) * $signed(input_fmap_125[7:0]) +
	( 15'sd 16248) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27362) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8812) * $signed(input_fmap_128[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_129[7:0]) +
	( 14'sd 7372) * $signed(input_fmap_130[7:0]) +
	( 16'sd 17412) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18136) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10241) * $signed(input_fmap_133[7:0]) +
	( 16'sd 27812) * $signed(input_fmap_134[7:0]) +
	( 15'sd 12787) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23242) * $signed(input_fmap_136[7:0]) +
	( 16'sd 23588) * $signed(input_fmap_137[7:0]) +
	( 16'sd 23873) * $signed(input_fmap_138[7:0]) +
	( 16'sd 22961) * $signed(input_fmap_139[7:0]) +
	( 15'sd 8309) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22566) * $signed(input_fmap_141[7:0]) +
	( 14'sd 4297) * $signed(input_fmap_142[7:0]) +
	( 16'sd 16519) * $signed(input_fmap_143[7:0]) +
	( 16'sd 29807) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17079) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3537) * $signed(input_fmap_146[7:0]) +
	( 12'sd 1767) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6074) * $signed(input_fmap_148[7:0]) +
	( 12'sd 1792) * $signed(input_fmap_149[7:0]) +
	( 16'sd 32565) * $signed(input_fmap_150[7:0]) +
	( 12'sd 1275) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14532) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2769) * $signed(input_fmap_153[7:0]) +
	( 13'sd 3044) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13014) * $signed(input_fmap_155[7:0]) +
	( 11'sd 593) * $signed(input_fmap_156[7:0]) +
	( 16'sd 17329) * $signed(input_fmap_157[7:0]) +
	( 15'sd 15579) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12477) * $signed(input_fmap_159[7:0]) +
	( 13'sd 3503) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1483) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10407) * $signed(input_fmap_162[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_165[7:0]) +
	( 16'sd 17361) * $signed(input_fmap_166[7:0]) +
	( 15'sd 10999) * $signed(input_fmap_167[7:0]) +
	( 16'sd 19464) * $signed(input_fmap_168[7:0]) +
	( 16'sd 16634) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9750) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19687) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14529) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1258) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10649) * $signed(input_fmap_174[7:0]) +
	( 11'sd 1014) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1358) * $signed(input_fmap_176[7:0]) +
	( 15'sd 10349) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27251) * $signed(input_fmap_178[7:0]) +
	( 15'sd 13825) * $signed(input_fmap_179[7:0]) +
	( 15'sd 14971) * $signed(input_fmap_180[7:0]) +
	( 14'sd 4802) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30184) * $signed(input_fmap_182[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31430) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5696) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25425) * $signed(input_fmap_187[7:0]) +
	( 16'sd 18119) * $signed(input_fmap_188[7:0]) +
	( 16'sd 21170) * $signed(input_fmap_189[7:0]) +
	( 15'sd 14799) * $signed(input_fmap_190[7:0]) +
	( 14'sd 4540) * $signed(input_fmap_191[7:0]) +
	( 16'sd 25906) * $signed(input_fmap_192[7:0]) +
	( 15'sd 8214) * $signed(input_fmap_193[7:0]) +
	( 14'sd 5433) * $signed(input_fmap_194[7:0]) +
	( 16'sd 26482) * $signed(input_fmap_195[7:0]) +
	( 15'sd 8644) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26513) * $signed(input_fmap_197[7:0]) +
	( 16'sd 16987) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10806) * $signed(input_fmap_199[7:0]) +
	( 16'sd 17194) * $signed(input_fmap_200[7:0]) +
	( 16'sd 32568) * $signed(input_fmap_201[7:0]) +
	( 15'sd 12532) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25319) * $signed(input_fmap_203[7:0]) +
	( 16'sd 24542) * $signed(input_fmap_204[7:0]) +
	( 16'sd 16775) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6181) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3368) * $signed(input_fmap_207[7:0]) +
	( 16'sd 26407) * $signed(input_fmap_208[7:0]) +
	( 12'sd 1709) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19292) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_211[7:0]) +
	( 15'sd 15615) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_213[7:0]) +
	( 16'sd 19232) * $signed(input_fmap_214[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23589) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17598) * $signed(input_fmap_217[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17556) * $signed(input_fmap_219[7:0]) +
	( 16'sd 27776) * $signed(input_fmap_220[7:0]) +
	( 15'sd 14579) * $signed(input_fmap_221[7:0]) +
	( 15'sd 13853) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14562) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19872) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14322) * $signed(input_fmap_225[7:0]) +
	( 16'sd 26405) * $signed(input_fmap_226[7:0]) +
	( 15'sd 10159) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26378) * $signed(input_fmap_228[7:0]) +
	( 14'sd 4719) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6779) * $signed(input_fmap_230[7:0]) +
	( 15'sd 9088) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7301) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27504) * $signed(input_fmap_233[7:0]) +
	( 16'sd 20990) * $signed(input_fmap_234[7:0]) +
	( 16'sd 30132) * $signed(input_fmap_235[7:0]) +
	( 14'sd 7890) * $signed(input_fmap_236[7:0]) +
	( 15'sd 15290) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16968) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21705) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23392) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5156) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_242[7:0]) +
	( 13'sd 3994) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28553) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19606) * $signed(input_fmap_245[7:0]) +
	( 16'sd 26727) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21824) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26574) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15938) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30558) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18968) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4459) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6361) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13329) * $signed(input_fmap_254[7:0]) +
	( 13'sd 3427) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_141;
assign conv_mac_141 = 
	( 13'sd 3880) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27950) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1663) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26267) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18728) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15528) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13124) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20475) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31154) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15653) * $signed(input_fmap_9[7:0]) +
	( 9'sd 134) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9414) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20426) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3552) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16464) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11137) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17472) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13159) * $signed(input_fmap_17[7:0]) +
	( 11'sd 781) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23023) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1367) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28640) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21963) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32202) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12837) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24076) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5167) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10225) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25574) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31312) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10556) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13263) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27523) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25236) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9071) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24311) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18940) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27889) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4901) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6165) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8294) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27088) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24955) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19820) * $signed(input_fmap_44[7:0]) +
	( 16'sd 32341) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13121) * $signed(input_fmap_46[7:0]) +
	( 10'sd 459) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8553) * $signed(input_fmap_49[7:0]) +
	( 11'sd 854) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2628) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19878) * $signed(input_fmap_52[7:0]) +
	( 14'sd 8134) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17616) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12020) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7745) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4496) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23710) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3515) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26140) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1716) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25244) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5234) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19575) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27525) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2955) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25519) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23596) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27226) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10979) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2484) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19339) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27382) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32205) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28901) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29006) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14479) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18445) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1247) * $signed(input_fmap_83[7:0]) +
	( 16'sd 16575) * $signed(input_fmap_84[7:0]) +
	( 15'sd 8743) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9047) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29342) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21380) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3937) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30024) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30201) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24325) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7175) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8213) * $signed(input_fmap_96[7:0]) +
	( 11'sd 794) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24211) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20638) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17397) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26070) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30586) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8539) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9034) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2416) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1124) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3719) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22656) * $signed(input_fmap_108[7:0]) +
	( 13'sd 4089) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28313) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28791) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24975) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31920) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3452) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1387) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31689) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13611) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7576) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10882) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5676) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26898) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14705) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6890) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10795) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18933) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30522) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4980) * $signed(input_fmap_127[7:0]) +
	( 16'sd 32323) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31667) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27841) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19686) * $signed(input_fmap_131[7:0]) +
	( 15'sd 9971) * $signed(input_fmap_132[7:0]) +
	( 16'sd 19588) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4160) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19686) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8382) * $signed(input_fmap_136[7:0]) +
	( 11'sd 955) * $signed(input_fmap_137[7:0]) +
	( 15'sd 12046) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28769) * $signed(input_fmap_139[7:0]) +
	( 16'sd 20623) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29305) * $signed(input_fmap_141[7:0]) +
	( 14'sd 4117) * $signed(input_fmap_142[7:0]) +
	( 15'sd 16117) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9748) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7874) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29074) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8447) * $signed(input_fmap_147[7:0]) +
	( 16'sd 29726) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18642) * $signed(input_fmap_149[7:0]) +
	( 14'sd 6413) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3108) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22882) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27021) * $signed(input_fmap_153[7:0]) +
	( 14'sd 8141) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5042) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13340) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18536) * $signed(input_fmap_157[7:0]) +
	( 15'sd 12363) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5780) * $signed(input_fmap_159[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_160[7:0]) +
	( 15'sd 8391) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26453) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27974) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25457) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2226) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18449) * $signed(input_fmap_166[7:0]) +
	( 16'sd 32727) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6226) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_169[7:0]) +
	( 15'sd 10431) * $signed(input_fmap_170[7:0]) +
	( 16'sd 29387) * $signed(input_fmap_171[7:0]) +
	( 16'sd 21368) * $signed(input_fmap_172[7:0]) +
	( 9'sd 218) * $signed(input_fmap_173[7:0]) +
	( 15'sd 12106) * $signed(input_fmap_174[7:0]) +
	( 16'sd 26092) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18130) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7648) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_178[7:0]) +
	( 16'sd 31945) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29226) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6927) * $signed(input_fmap_181[7:0]) +
	( 11'sd 549) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25503) * $signed(input_fmap_183[7:0]) +
	( 13'sd 2657) * $signed(input_fmap_184[7:0]) +
	( 15'sd 9780) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_186[7:0]) +
	( 14'sd 6426) * $signed(input_fmap_187[7:0]) +
	( 15'sd 11479) * $signed(input_fmap_188[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_189[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_190[7:0]) +
	( 16'sd 27225) * $signed(input_fmap_191[7:0]) +
	( 14'sd 5256) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12135) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21778) * $signed(input_fmap_194[7:0]) +
	( 16'sd 28739) * $signed(input_fmap_195[7:0]) +
	( 16'sd 21731) * $signed(input_fmap_196[7:0]) +
	( 16'sd 32696) * $signed(input_fmap_197[7:0]) +
	( 14'sd 7971) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31925) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6291) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7568) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19101) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11842) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20552) * $signed(input_fmap_206[7:0]) +
	( 16'sd 16583) * $signed(input_fmap_207[7:0]) +
	( 13'sd 2994) * $signed(input_fmap_208[7:0]) +
	( 15'sd 8704) * $signed(input_fmap_209[7:0]) +
	( 16'sd 28533) * $signed(input_fmap_210[7:0]) +
	( 13'sd 2818) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24006) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3221) * $signed(input_fmap_213[7:0]) +
	( 16'sd 19889) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25146) * $signed(input_fmap_215[7:0]) +
	( 15'sd 12109) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19176) * $signed(input_fmap_217[7:0]) +
	( 11'sd 651) * $signed(input_fmap_218[7:0]) +
	( 12'sd 1917) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14730) * $signed(input_fmap_220[7:0]) +
	( 16'sd 30015) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18536) * $signed(input_fmap_222[7:0]) +
	( 16'sd 32043) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30805) * $signed(input_fmap_224[7:0]) +
	( 16'sd 21876) * $signed(input_fmap_225[7:0]) +
	( 16'sd 19807) * $signed(input_fmap_226[7:0]) +
	( 12'sd 1288) * $signed(input_fmap_227[7:0]) +
	( 14'sd 5044) * $signed(input_fmap_228[7:0]) +
	( 13'sd 2448) * $signed(input_fmap_229[7:0]) +
	( 10'sd 375) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3463) * $signed(input_fmap_231[7:0]) +
	( 16'sd 26031) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5355) * $signed(input_fmap_233[7:0]) +
	( 16'sd 16941) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12095) * $signed(input_fmap_235[7:0]) +
	( 16'sd 29748) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10620) * $signed(input_fmap_237[7:0]) +
	( 15'sd 9513) * $signed(input_fmap_238[7:0]) +
	( 16'sd 17643) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18910) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20738) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22436) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20824) * $signed(input_fmap_244[7:0]) +
	( 16'sd 31836) * $signed(input_fmap_245[7:0]) +
	( 14'sd 4694) * $signed(input_fmap_246[7:0]) +
	( 16'sd 29828) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4653) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3003) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3153) * $signed(input_fmap_250[7:0]) +
	( 16'sd 17773) * $signed(input_fmap_251[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5004) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23011) * $signed(input_fmap_254[7:0]) +
	( 12'sd 1306) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_142;
assign conv_mac_142 = 
	( 14'sd 6676) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21204) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21896) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21882) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21049) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2656) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22534) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8398) * $signed(input_fmap_7[7:0]) +
	( 10'sd 343) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25749) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23062) * $signed(input_fmap_10[7:0]) +
	( 9'sd 208) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2952) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20815) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32279) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5346) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16133) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2795) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8409) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20649) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6779) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21023) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24571) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16785) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2085) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23022) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17876) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16983) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27994) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13534) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12004) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8245) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21805) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11387) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29771) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4263) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15304) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26733) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8196) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29865) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32565) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11005) * $signed(input_fmap_43[7:0]) +
	( 15'sd 8983) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1607) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28254) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15159) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13431) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22559) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31078) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32468) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27450) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2848) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17388) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12388) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17577) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11107) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17340) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29188) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21982) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12688) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22003) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18685) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27895) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22660) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17167) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27065) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32623) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4194) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23288) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2200) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2251) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2630) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24482) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3866) * $signed(input_fmap_78[7:0]) +
	( 13'sd 2546) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24925) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27210) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24471) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12723) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28505) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32709) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17584) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32492) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26527) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30011) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24700) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6800) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30510) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10970) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5507) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26741) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28974) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18993) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3570) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21636) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30894) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13273) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5025) * $signed(input_fmap_104[7:0]) +
	( 16'sd 19271) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27862) * $signed(input_fmap_106[7:0]) +
	( 11'sd 809) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15545) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29282) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27706) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13126) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16283) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21751) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13197) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9196) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8690) * $signed(input_fmap_117[7:0]) +
	( 15'sd 8715) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3529) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24485) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18534) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17077) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15665) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22540) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16399) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30735) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28436) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31689) * $signed(input_fmap_130[7:0]) +
	( 15'sd 10381) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5288) * $signed(input_fmap_132[7:0]) +
	( 16'sd 23144) * $signed(input_fmap_133[7:0]) +
	( 16'sd 30573) * $signed(input_fmap_134[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31600) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24241) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31427) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31151) * $signed(input_fmap_139[7:0]) +
	( 14'sd 7290) * $signed(input_fmap_140[7:0]) +
	( 13'sd 2872) * $signed(input_fmap_141[7:0]) +
	( 15'sd 13490) * $signed(input_fmap_142[7:0]) +
	( 16'sd 25497) * $signed(input_fmap_143[7:0]) +
	( 14'sd 8121) * $signed(input_fmap_144[7:0]) +
	( 15'sd 15789) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14416) * $signed(input_fmap_146[7:0]) +
	( 13'sd 2809) * $signed(input_fmap_147[7:0]) +
	( 15'sd 10133) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12888) * $signed(input_fmap_149[7:0]) +
	( 16'sd 26820) * $signed(input_fmap_150[7:0]) +
	( 15'sd 15237) * $signed(input_fmap_151[7:0]) +
	( 16'sd 32693) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12027) * $signed(input_fmap_153[7:0]) +
	( 16'sd 27188) * $signed(input_fmap_154[7:0]) +
	( 13'sd 3490) * $signed(input_fmap_155[7:0]) +
	( 16'sd 28922) * $signed(input_fmap_156[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_157[7:0]) +
	( 16'sd 24304) * $signed(input_fmap_158[7:0]) +
	( 16'sd 23724) * $signed(input_fmap_159[7:0]) +
	( 16'sd 19713) * $signed(input_fmap_160[7:0]) +
	( 16'sd 29844) * $signed(input_fmap_161[7:0]) +
	( 16'sd 31504) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30766) * $signed(input_fmap_163[7:0]) +
	( 16'sd 31755) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_165[7:0]) +
	( 16'sd 29981) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13691) * $signed(input_fmap_167[7:0]) +
	( 15'sd 13438) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10250) * $signed(input_fmap_169[7:0]) +
	( 16'sd 21165) * $signed(input_fmap_170[7:0]) +
	( 15'sd 8772) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14898) * $signed(input_fmap_172[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_173[7:0]) +
	( 15'sd 13441) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1227) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3407) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2483) * $signed(input_fmap_177[7:0]) +
	( 16'sd 16549) * $signed(input_fmap_178[7:0]) +
	( 16'sd 26823) * $signed(input_fmap_179[7:0]) +
	( 12'sd 1340) * $signed(input_fmap_180[7:0]) +
	( 16'sd 20572) * $signed(input_fmap_181[7:0]) +
	( 16'sd 27150) * $signed(input_fmap_182[7:0]) +
	( 15'sd 8196) * $signed(input_fmap_183[7:0]) +
	( 16'sd 32329) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5885) * $signed(input_fmap_185[7:0]) +
	( 15'sd 14281) * $signed(input_fmap_186[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_187[7:0]) +
	( 16'sd 25951) * $signed(input_fmap_188[7:0]) +
	( 12'sd 1611) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31290) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17031) * $signed(input_fmap_191[7:0]) +
	( 16'sd 25109) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9278) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13737) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24906) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19620) * $signed(input_fmap_197[7:0]) +
	( 14'sd 6266) * $signed(input_fmap_198[7:0]) +
	( 15'sd 11322) * $signed(input_fmap_199[7:0]) +
	( 16'sd 21217) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22959) * $signed(input_fmap_201[7:0]) +
	( 16'sd 29636) * $signed(input_fmap_202[7:0]) +
	( 12'sd 1559) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4775) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28155) * $signed(input_fmap_205[7:0]) +
	( 15'sd 14943) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21348) * $signed(input_fmap_207[7:0]) +
	( 13'sd 3167) * $signed(input_fmap_208[7:0]) +
	( 16'sd 17983) * $signed(input_fmap_209[7:0]) +
	( 16'sd 24153) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11789) * $signed(input_fmap_212[7:0]) +
	( 16'sd 22301) * $signed(input_fmap_213[7:0]) +
	( 13'sd 3839) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5988) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17429) * $signed(input_fmap_216[7:0]) +
	( 13'sd 2641) * $signed(input_fmap_217[7:0]) +
	( 15'sd 12574) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20069) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_220[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28444) * $signed(input_fmap_222[7:0]) +
	( 16'sd 16863) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7428) * $signed(input_fmap_224[7:0]) +
	( 15'sd 10389) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29857) * $signed(input_fmap_226[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_227[7:0]) +
	( 14'sd 7706) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3565) * $signed(input_fmap_229[7:0]) +
	( 16'sd 22658) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25677) * $signed(input_fmap_231[7:0]) +
	( 12'sd 1243) * $signed(input_fmap_232[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_233[7:0]) +
	( 15'sd 10732) * $signed(input_fmap_234[7:0]) +
	( 16'sd 20668) * $signed(input_fmap_235[7:0]) +
	( 16'sd 26150) * $signed(input_fmap_236[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3284) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26247) * $signed(input_fmap_239[7:0]) +
	( 16'sd 27544) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15064) * $signed(input_fmap_242[7:0]) +
	( 15'sd 8540) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18743) * $signed(input_fmap_244[7:0]) +
	( 16'sd 18580) * $signed(input_fmap_245[7:0]) +
	( 15'sd 12976) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18473) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13612) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30133) * $signed(input_fmap_249[7:0]) +
	( 14'sd 4872) * $signed(input_fmap_250[7:0]) +
	( 16'sd 16779) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4931) * $signed(input_fmap_252[7:0]) +
	( 16'sd 30913) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1311) * $signed(input_fmap_254[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_143;
assign conv_mac_143 = 
	( 16'sd 31476) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23004) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32071) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13439) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25117) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27476) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16376) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12821) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24028) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12473) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8705) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32288) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29634) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2283) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13779) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16188) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30237) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18354) * $signed(input_fmap_18[7:0]) +
	( 13'sd 3878) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30903) * $signed(input_fmap_20[7:0]) +
	( 15'sd 8465) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5990) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13904) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31182) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22620) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5900) * $signed(input_fmap_26[7:0]) +
	( 15'sd 12424) * $signed(input_fmap_27[7:0]) +
	( 15'sd 16007) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3075) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2603) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9689) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23065) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8778) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7751) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2117) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30076) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16738) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17095) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22054) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6797) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21379) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14091) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9061) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27164) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21585) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13257) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6537) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7950) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5281) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4382) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7685) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14397) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20018) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5742) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12294) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26657) * $signed(input_fmap_59[7:0]) +
	( 13'sd 4025) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32304) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25194) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6776) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15149) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21695) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15587) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22030) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30598) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11092) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21578) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32436) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14751) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28787) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6928) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27206) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7522) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7603) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7535) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28459) * $signed(input_fmap_79[7:0]) +
	( 10'sd 300) * $signed(input_fmap_80[7:0]) +
	( 16'sd 32312) * $signed(input_fmap_81[7:0]) +
	( 13'sd 4065) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29897) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20416) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14940) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24628) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18715) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5100) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29122) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26441) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27557) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17249) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15861) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31022) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10146) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32045) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26381) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4473) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29293) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6873) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12601) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7810) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25992) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5731) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13437) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5025) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15598) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27397) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18203) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6711) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12223) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12580) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22933) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18461) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1454) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13809) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28761) * $signed(input_fmap_119[7:0]) +
	( 15'sd 14195) * $signed(input_fmap_120[7:0]) +
	( 13'sd 4003) * $signed(input_fmap_121[7:0]) +
	( 14'sd 8131) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13037) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12152) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2762) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5716) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23224) * $signed(input_fmap_128[7:0]) +
	( 14'sd 4878) * $signed(input_fmap_129[7:0]) +
	( 15'sd 11590) * $signed(input_fmap_130[7:0]) +
	( 12'sd 1240) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10409) * $signed(input_fmap_132[7:0]) +
	( 14'sd 4168) * $signed(input_fmap_133[7:0]) +
	( 9'sd 138) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23910) * $signed(input_fmap_135[7:0]) +
	( 16'sd 24394) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15965) * $signed(input_fmap_137[7:0]) +
	( 11'sd 562) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8259) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24404) * $signed(input_fmap_140[7:0]) +
	( 16'sd 23740) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22031) * $signed(input_fmap_142[7:0]) +
	( 15'sd 13108) * $signed(input_fmap_143[7:0]) +
	( 16'sd 16483) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25855) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_146[7:0]) +
	( 16'sd 16735) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4422) * $signed(input_fmap_148[7:0]) +
	( 15'sd 16057) * $signed(input_fmap_149[7:0]) +
	( 15'sd 11708) * $signed(input_fmap_150[7:0]) +
	( 12'sd 1932) * $signed(input_fmap_151[7:0]) +
	( 12'sd 1831) * $signed(input_fmap_152[7:0]) +
	( 16'sd 28792) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6765) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19553) * $signed(input_fmap_155[7:0]) +
	( 15'sd 9974) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_157[7:0]) +
	( 16'sd 30525) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3087) * $signed(input_fmap_159[7:0]) +
	( 16'sd 28432) * $signed(input_fmap_160[7:0]) +
	( 13'sd 3442) * $signed(input_fmap_161[7:0]) +
	( 14'sd 7510) * $signed(input_fmap_162[7:0]) +
	( 15'sd 9846) * $signed(input_fmap_163[7:0]) +
	( 16'sd 32523) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22608) * $signed(input_fmap_165[7:0]) +
	( 11'sd 905) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20199) * $signed(input_fmap_167[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18893) * $signed(input_fmap_169[7:0]) +
	( 12'sd 1895) * $signed(input_fmap_170[7:0]) +
	( 16'sd 27786) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31115) * $signed(input_fmap_172[7:0]) +
	( 11'sd 621) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27398) * $signed(input_fmap_174[7:0]) +
	( 15'sd 10424) * $signed(input_fmap_175[7:0]) +
	( 16'sd 28459) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5208) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2438) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15526) * $signed(input_fmap_179[7:0]) +
	( 8'sd 84) * $signed(input_fmap_180[7:0]) +
	( 16'sd 27237) * $signed(input_fmap_181[7:0]) +
	( 16'sd 18606) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12928) * $signed(input_fmap_183[7:0]) +
	( 16'sd 25293) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7837) * $signed(input_fmap_185[7:0]) +
	( 15'sd 14010) * $signed(input_fmap_186[7:0]) +
	( 15'sd 10355) * $signed(input_fmap_187[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_188[7:0]) +
	( 15'sd 16268) * $signed(input_fmap_189[7:0]) +
	( 15'sd 14416) * $signed(input_fmap_190[7:0]) +
	( 14'sd 4879) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31945) * $signed(input_fmap_192[7:0]) +
	( 16'sd 25643) * $signed(input_fmap_193[7:0]) +
	( 12'sd 1397) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_195[7:0]) +
	( 16'sd 21202) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15386) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29767) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25954) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11797) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17294) * $signed(input_fmap_202[7:0]) +
	( 16'sd 23482) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12418) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1131) * $signed(input_fmap_205[7:0]) +
	( 14'sd 7159) * $signed(input_fmap_206[7:0]) +
	( 16'sd 16740) * $signed(input_fmap_207[7:0]) +
	( 13'sd 3384) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7060) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3413) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20699) * $signed(input_fmap_211[7:0]) +
	( 15'sd 8277) * $signed(input_fmap_212[7:0]) +
	( 16'sd 25382) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_214[7:0]) +
	( 16'sd 27154) * $signed(input_fmap_215[7:0]) +
	( 16'sd 29388) * $signed(input_fmap_216[7:0]) +
	( 13'sd 2222) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5332) * $signed(input_fmap_218[7:0]) +
	( 16'sd 32379) * $signed(input_fmap_219[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_220[7:0]) +
	( 16'sd 17936) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28971) * $signed(input_fmap_223[7:0]) +
	( 14'sd 5853) * $signed(input_fmap_224[7:0]) +
	( 16'sd 19706) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11438) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22628) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_228[7:0]) +
	( 15'sd 15857) * $signed(input_fmap_229[7:0]) +
	( 15'sd 10817) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_231[7:0]) +
	( 12'sd 1756) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24994) * $signed(input_fmap_233[7:0]) +
	( 16'sd 17532) * $signed(input_fmap_234[7:0]) +
	( 8'sd 124) * $signed(input_fmap_235[7:0]) +
	( 16'sd 21286) * $signed(input_fmap_236[7:0]) +
	( 15'sd 9368) * $signed(input_fmap_237[7:0]) +
	( 16'sd 30175) * $signed(input_fmap_238[7:0]) +
	( 16'sd 18973) * $signed(input_fmap_239[7:0]) +
	( 13'sd 3892) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7669) * $signed(input_fmap_241[7:0]) +
	( 13'sd 3347) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7026) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13223) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19138) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23767) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_247[7:0]) +
	( 16'sd 31598) * $signed(input_fmap_248[7:0]) +
	( 14'sd 6810) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24666) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2650) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20416) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6557) * $signed(input_fmap_253[7:0]) +
	( 15'sd 12457) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26142) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_144;
assign conv_mac_144 = 
	( 16'sd 22598) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8834) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11393) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19890) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23829) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3942) * $signed(input_fmap_6[7:0]) +
	( 9'sd 142) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24866) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3005) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27470) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12178) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28922) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17940) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10966) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6575) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9374) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26644) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24269) * $signed(input_fmap_21[7:0]) +
	( 11'sd 953) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22991) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11127) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20320) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_26[7:0]) +
	( 11'sd 997) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19390) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20421) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1150) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17277) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2356) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12824) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14812) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9732) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6086) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32496) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21470) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26833) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29073) * $signed(input_fmap_40[7:0]) +
	( 5'sd 14) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24496) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26025) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6289) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29872) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9610) * $signed(input_fmap_46[7:0]) +
	( 11'sd 839) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22156) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22078) * $signed(input_fmap_49[7:0]) +
	( 16'sd 31298) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18760) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10391) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31405) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19531) * $signed(input_fmap_54[7:0]) +
	( 14'sd 8117) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12402) * $signed(input_fmap_56[7:0]) +
	( 13'sd 3375) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3765) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10524) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2935) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12258) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_62[7:0]) +
	( 10'sd 304) * $signed(input_fmap_63[7:0]) +
	( 16'sd 26872) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21859) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8796) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6981) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8876) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29039) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27388) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_74[7:0]) +
	( 9'sd 224) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20777) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23592) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25941) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13925) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18875) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4343) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21238) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30205) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28554) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11721) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10471) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10961) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3714) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11111) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29854) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23492) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5986) * $signed(input_fmap_93[7:0]) +
	( 16'sd 19818) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7884) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26076) * $signed(input_fmap_96[7:0]) +
	( 16'sd 21171) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21278) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24733) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12079) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15761) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30352) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24839) * $signed(input_fmap_104[7:0]) +
	( 11'sd 748) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21789) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6322) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22945) * $signed(input_fmap_108[7:0]) +
	( 10'sd 323) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29801) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25377) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24499) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27023) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4883) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12269) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19873) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18733) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8321) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8363) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24215) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13783) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17025) * $signed(input_fmap_124[7:0]) +
	( 14'sd 8149) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10060) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27213) * $signed(input_fmap_127[7:0]) +
	( 16'sd 25525) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17941) * $signed(input_fmap_129[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20559) * $signed(input_fmap_131[7:0]) +
	( 16'sd 24050) * $signed(input_fmap_132[7:0]) +
	( 14'sd 4861) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24996) * $signed(input_fmap_134[7:0]) +
	( 16'sd 29240) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7752) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24062) * $signed(input_fmap_137[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27043) * $signed(input_fmap_139[7:0]) +
	( 16'sd 32072) * $signed(input_fmap_140[7:0]) +
	( 14'sd 6949) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28804) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23346) * $signed(input_fmap_143[7:0]) +
	( 12'sd 2023) * $signed(input_fmap_144[7:0]) +
	( 15'sd 15580) * $signed(input_fmap_145[7:0]) +
	( 15'sd 16017) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3824) * $signed(input_fmap_147[7:0]) +
	( 15'sd 13049) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18744) * $signed(input_fmap_150[7:0]) +
	( 16'sd 25907) * $signed(input_fmap_151[7:0]) +
	( 16'sd 17231) * $signed(input_fmap_152[7:0]) +
	( 15'sd 8796) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4215) * $signed(input_fmap_154[7:0]) +
	( 15'sd 14729) * $signed(input_fmap_155[7:0]) +
	( 16'sd 23903) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27116) * $signed(input_fmap_157[7:0]) +
	( 13'sd 2533) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21510) * $signed(input_fmap_159[7:0]) +
	( 14'sd 8050) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13038) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32495) * $signed(input_fmap_163[7:0]) +
	( 16'sd 20477) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28702) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18619) * $signed(input_fmap_166[7:0]) +
	( 16'sd 18440) * $signed(input_fmap_167[7:0]) +
	( 15'sd 11512) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6361) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28124) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30774) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4685) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18488) * $signed(input_fmap_173[7:0]) +
	( 15'sd 9892) * $signed(input_fmap_174[7:0]) +
	( 16'sd 30986) * $signed(input_fmap_175[7:0]) +
	( 16'sd 32014) * $signed(input_fmap_176[7:0]) +
	( 16'sd 32695) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22496) * $signed(input_fmap_178[7:0]) +
	( 14'sd 7265) * $signed(input_fmap_179[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_180[7:0]) +
	( 12'sd 1939) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30117) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29099) * $signed(input_fmap_183[7:0]) +
	( 16'sd 29882) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7836) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23778) * $signed(input_fmap_186[7:0]) +
	( 16'sd 24830) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4299) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7815) * $signed(input_fmap_189[7:0]) +
	( 12'sd 1256) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23498) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22504) * $signed(input_fmap_192[7:0]) +
	( 16'sd 17137) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3487) * $signed(input_fmap_194[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14982) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22459) * $signed(input_fmap_197[7:0]) +
	( 15'sd 13574) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1795) * $signed(input_fmap_199[7:0]) +
	( 16'sd 19621) * $signed(input_fmap_200[7:0]) +
	( 16'sd 19542) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14667) * $signed(input_fmap_202[7:0]) +
	( 16'sd 31490) * $signed(input_fmap_203[7:0]) +
	( 16'sd 22140) * $signed(input_fmap_204[7:0]) +
	( 16'sd 22767) * $signed(input_fmap_205[7:0]) +
	( 16'sd 25680) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17854) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8837) * $signed(input_fmap_208[7:0]) +
	( 15'sd 9643) * $signed(input_fmap_209[7:0]) +
	( 11'sd 1001) * $signed(input_fmap_210[7:0]) +
	( 16'sd 24383) * $signed(input_fmap_211[7:0]) +
	( 14'sd 8149) * $signed(input_fmap_212[7:0]) +
	( 16'sd 32266) * $signed(input_fmap_213[7:0]) +
	( 14'sd 5481) * $signed(input_fmap_214[7:0]) +
	( 16'sd 28680) * $signed(input_fmap_215[7:0]) +
	( 15'sd 10615) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32358) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7729) * $signed(input_fmap_218[7:0]) +
	( 12'sd 1890) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4884) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5421) * $signed(input_fmap_221[7:0]) +
	( 16'sd 23601) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25250) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25640) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5224) * $signed(input_fmap_225[7:0]) +
	( 16'sd 25067) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5111) * $signed(input_fmap_227[7:0]) +
	( 15'sd 9180) * $signed(input_fmap_228[7:0]) +
	( 12'sd 1827) * $signed(input_fmap_229[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_230[7:0]) +
	( 15'sd 12367) * $signed(input_fmap_231[7:0]) +
	( 14'sd 6137) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21398) * $signed(input_fmap_233[7:0]) +
	( 16'sd 32218) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19143) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31161) * $signed(input_fmap_236[7:0]) +
	( 13'sd 3644) * $signed(input_fmap_237[7:0]) +
	( 16'sd 24956) * $signed(input_fmap_238[7:0]) +
	( 14'sd 4806) * $signed(input_fmap_239[7:0]) +
	( 14'sd 4325) * $signed(input_fmap_240[7:0]) +
	( 16'sd 27351) * $signed(input_fmap_241[7:0]) +
	( 16'sd 32497) * $signed(input_fmap_242[7:0]) +
	( 15'sd 8805) * $signed(input_fmap_243[7:0]) +
	( 16'sd 31498) * $signed(input_fmap_244[7:0]) +
	( 16'sd 29339) * $signed(input_fmap_245[7:0]) +
	( 14'sd 7969) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17465) * $signed(input_fmap_247[7:0]) +
	( 16'sd 23868) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30039) * $signed(input_fmap_249[7:0]) +
	( 16'sd 27804) * $signed(input_fmap_250[7:0]) +
	( 16'sd 32385) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4921) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24717) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2214) * $signed(input_fmap_254[7:0]) +
	( 14'sd 6485) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_145;
assign conv_mac_145 = 
	( 16'sd 19253) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19687) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25595) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25983) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3300) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15488) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2474) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18242) * $signed(input_fmap_7[7:0]) +
	( 16'sd 21711) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12729) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18629) * $signed(input_fmap_10[7:0]) +
	( 11'sd 580) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17694) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20807) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28420) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5422) * $signed(input_fmap_16[7:0]) +
	( 15'sd 16359) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13611) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14464) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22110) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19779) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9767) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22311) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31157) * $signed(input_fmap_24[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19320) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15249) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12918) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26844) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4163) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3840) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2682) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30644) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10082) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31702) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17423) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1079) * $signed(input_fmap_37[7:0]) +
	( 14'sd 8178) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17099) * $signed(input_fmap_39[7:0]) +
	( 11'sd 623) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6642) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16940) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11089) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21077) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12017) * $signed(input_fmap_45[7:0]) +
	( 10'sd 283) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24762) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13049) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24268) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18727) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26223) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4800) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10553) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21934) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28726) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32265) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28864) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24250) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23049) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10585) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17857) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18598) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10377) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12817) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10863) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14976) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31795) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15257) * $signed(input_fmap_72[7:0]) +
	( 11'sd 956) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14198) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7170) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12938) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21515) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3519) * $signed(input_fmap_79[7:0]) +
	( 16'sd 18560) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31941) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5605) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2662) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3546) * $signed(input_fmap_84[7:0]) +
	( 11'sd 829) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2142) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17946) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3855) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21646) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26366) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26052) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25145) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23760) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4539) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3466) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30531) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7631) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28510) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25043) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16626) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11799) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26827) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25437) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_104[7:0]) +
	( 16'sd 22224) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23315) * $signed(input_fmap_106[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5309) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5992) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15599) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31953) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3928) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3141) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6393) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17189) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19988) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13122) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3916) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27822) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26863) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20062) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30031) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24782) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24598) * $signed(input_fmap_127[7:0]) +
	( 13'sd 3843) * $signed(input_fmap_128[7:0]) +
	( 13'sd 2570) * $signed(input_fmap_129[7:0]) +
	( 14'sd 7293) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11831) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16454) * $signed(input_fmap_133[7:0]) +
	( 16'sd 23146) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27724) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_136[7:0]) +
	( 16'sd 21942) * $signed(input_fmap_137[7:0]) +
	( 16'sd 20589) * $signed(input_fmap_138[7:0]) +
	( 16'sd 17846) * $signed(input_fmap_139[7:0]) +
	( 15'sd 10924) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5213) * $signed(input_fmap_141[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_142[7:0]) +
	( 16'sd 16781) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13031) * $signed(input_fmap_144[7:0]) +
	( 14'sd 4292) * $signed(input_fmap_145[7:0]) +
	( 14'sd 8110) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3765) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28027) * $signed(input_fmap_148[7:0]) +
	( 16'sd 29073) * $signed(input_fmap_149[7:0]) +
	( 13'sd 2726) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19433) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6739) * $signed(input_fmap_152[7:0]) +
	( 16'sd 29827) * $signed(input_fmap_153[7:0]) +
	( 13'sd 3716) * $signed(input_fmap_154[7:0]) +
	( 16'sd 26521) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24518) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30233) * $signed(input_fmap_157[7:0]) +
	( 14'sd 5287) * $signed(input_fmap_158[7:0]) +
	( 16'sd 25959) * $signed(input_fmap_159[7:0]) +
	( 16'sd 28409) * $signed(input_fmap_160[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14427) * $signed(input_fmap_162[7:0]) +
	( 12'sd 1410) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6167) * $signed(input_fmap_164[7:0]) +
	( 16'sd 17994) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2486) * $signed(input_fmap_166[7:0]) +
	( 14'sd 4211) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14325) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17150) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7923) * $signed(input_fmap_170[7:0]) +
	( 16'sd 27342) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19384) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5245) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14370) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5761) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1153) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22728) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22807) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22758) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3277) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23741) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19239) * $signed(input_fmap_182[7:0]) +
	( 15'sd 9557) * $signed(input_fmap_183[7:0]) +
	( 16'sd 29088) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15341) * $signed(input_fmap_185[7:0]) +
	( 15'sd 11089) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28293) * $signed(input_fmap_187[7:0]) +
	( 15'sd 10147) * $signed(input_fmap_188[7:0]) +
	( 15'sd 14034) * $signed(input_fmap_189[7:0]) +
	( 15'sd 11460) * $signed(input_fmap_190[7:0]) +
	( 16'sd 28679) * $signed(input_fmap_191[7:0]) +
	( 16'sd 25582) * $signed(input_fmap_192[7:0]) +
	( 16'sd 25527) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3663) * $signed(input_fmap_194[7:0]) +
	( 14'sd 4867) * $signed(input_fmap_195[7:0]) +
	( 16'sd 21235) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19272) * $signed(input_fmap_197[7:0]) +
	( 11'sd 782) * $signed(input_fmap_198[7:0]) +
	( 14'sd 4927) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6979) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13209) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18681) * $signed(input_fmap_202[7:0]) +
	( 16'sd 16830) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15136) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31609) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9817) * $signed(input_fmap_206[7:0]) +
	( 16'sd 24162) * $signed(input_fmap_207[7:0]) +
	( 16'sd 29662) * $signed(input_fmap_208[7:0]) +
	( 16'sd 27976) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17233) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24000) * $signed(input_fmap_212[7:0]) +
	( 16'sd 22644) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30394) * $signed(input_fmap_214[7:0]) +
	( 16'sd 21979) * $signed(input_fmap_215[7:0]) +
	( 13'sd 3661) * $signed(input_fmap_216[7:0]) +
	( 16'sd 21573) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22815) * $signed(input_fmap_218[7:0]) +
	( 16'sd 29042) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19439) * $signed(input_fmap_220[7:0]) +
	( 14'sd 4619) * $signed(input_fmap_221[7:0]) +
	( 16'sd 17059) * $signed(input_fmap_222[7:0]) +
	( 14'sd 6661) * $signed(input_fmap_223[7:0]) +
	( 16'sd 22997) * $signed(input_fmap_224[7:0]) +
	( 16'sd 32002) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27116) * $signed(input_fmap_226[7:0]) +
	( 16'sd 23262) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22026) * $signed(input_fmap_228[7:0]) +
	( 16'sd 30323) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15898) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17155) * $signed(input_fmap_231[7:0]) +
	( 13'sd 3871) * $signed(input_fmap_232[7:0]) +
	( 15'sd 8922) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4135) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5710) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11100) * $signed(input_fmap_236[7:0]) +
	( 16'sd 17386) * $signed(input_fmap_237[7:0]) +
	( 12'sd 1884) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9362) * $signed(input_fmap_239[7:0]) +
	( 13'sd 3175) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15929) * $signed(input_fmap_241[7:0]) +
	( 13'sd 2100) * $signed(input_fmap_242[7:0]) +
	( 14'sd 4910) * $signed(input_fmap_243[7:0]) +
	( 16'sd 17726) * $signed(input_fmap_244[7:0]) +
	( 16'sd 26268) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11557) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30928) * $signed(input_fmap_247[7:0]) +
	( 16'sd 24654) * $signed(input_fmap_248[7:0]) +
	( 11'sd 567) * $signed(input_fmap_249[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20032) * $signed(input_fmap_252[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_253[7:0]) +
	( 16'sd 21201) * $signed(input_fmap_254[7:0]) +
	( 16'sd 25266) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_146;
assign conv_mac_146 = 
	( 16'sd 19978) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18706) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14170) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20728) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30135) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11782) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4174) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32741) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9610) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16749) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6936) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19284) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1723) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2947) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14482) * $signed(input_fmap_16[7:0]) +
	( 11'sd 741) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32564) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13156) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14111) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13428) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25855) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31283) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6554) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16158) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22247) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13410) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20849) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10183) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30651) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1626) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18068) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1317) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2603) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15109) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27554) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18990) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32206) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29775) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25568) * $signed(input_fmap_41[7:0]) +
	( 14'sd 7133) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16658) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3346) * $signed(input_fmap_44[7:0]) +
	( 16'sd 19573) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3902) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5326) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4536) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17702) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4563) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5384) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26559) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29707) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8905) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20208) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10143) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15708) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28360) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19982) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17525) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28270) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1231) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28533) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27652) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30179) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_68[7:0]) +
	( 15'sd 12498) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20020) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26335) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25847) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30512) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15611) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16092) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19742) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17071) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24658) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16781) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20593) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27021) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18568) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4161) * $signed(input_fmap_89[7:0]) +
	( 9'sd 190) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5728) * $signed(input_fmap_91[7:0]) +
	( 11'sd 881) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7331) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1359) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22455) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19214) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27314) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4274) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5847) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22272) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5940) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4110) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10475) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26794) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25934) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16400) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14778) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5773) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14826) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31387) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8462) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18087) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28959) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5309) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24020) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12053) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18447) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13166) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18931) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20117) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2134) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13813) * $signed(input_fmap_123[7:0]) +
	( 4'sd 6) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25146) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25571) * $signed(input_fmap_127[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_128[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_129[7:0]) +
	( 13'sd 3222) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14318) * $signed(input_fmap_131[7:0]) +
	( 13'sd 3943) * $signed(input_fmap_132[7:0]) +
	( 16'sd 26289) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31936) * $signed(input_fmap_135[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_136[7:0]) +
	( 16'sd 31159) * $signed(input_fmap_137[7:0]) +
	( 14'sd 4883) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_139[7:0]) +
	( 16'sd 16909) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22361) * $signed(input_fmap_141[7:0]) +
	( 15'sd 16028) * $signed(input_fmap_142[7:0]) +
	( 15'sd 9388) * $signed(input_fmap_143[7:0]) +
	( 15'sd 8288) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3786) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29847) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23694) * $signed(input_fmap_148[7:0]) +
	( 14'sd 8091) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5628) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17703) * $signed(input_fmap_151[7:0]) +
	( 12'sd 1498) * $signed(input_fmap_152[7:0]) +
	( 15'sd 9981) * $signed(input_fmap_153[7:0]) +
	( 16'sd 27937) * $signed(input_fmap_154[7:0]) +
	( 13'sd 3641) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24606) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14529) * $signed(input_fmap_157[7:0]) +
	( 16'sd 21983) * $signed(input_fmap_158[7:0]) +
	( 16'sd 23444) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17004) * $signed(input_fmap_160[7:0]) +
	( 15'sd 10680) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29908) * $signed(input_fmap_162[7:0]) +
	( 15'sd 12293) * $signed(input_fmap_163[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28567) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18876) * $signed(input_fmap_166[7:0]) +
	( 16'sd 32149) * $signed(input_fmap_167[7:0]) +
	( 13'sd 3684) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25612) * $signed(input_fmap_169[7:0]) +
	( 15'sd 12685) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11831) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_173[7:0]) +
	( 13'sd 2610) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3646) * $signed(input_fmap_175[7:0]) +
	( 16'sd 24268) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30717) * $signed(input_fmap_177[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_178[7:0]) +
	( 15'sd 9463) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23003) * $signed(input_fmap_180[7:0]) +
	( 14'sd 5686) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30771) * $signed(input_fmap_182[7:0]) +
	( 16'sd 22286) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26225) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11744) * $signed(input_fmap_185[7:0]) +
	( 15'sd 15373) * $signed(input_fmap_186[7:0]) +
	( 16'sd 21444) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1054) * $signed(input_fmap_188[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_189[7:0]) +
	( 15'sd 10848) * $signed(input_fmap_190[7:0]) +
	( 15'sd 10462) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20906) * $signed(input_fmap_192[7:0]) +
	( 16'sd 17016) * $signed(input_fmap_193[7:0]) +
	( 16'sd 28072) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1877) * $signed(input_fmap_195[7:0]) +
	( 16'sd 31858) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31021) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18313) * $signed(input_fmap_198[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_199[7:0]) +
	( 15'sd 9687) * $signed(input_fmap_200[7:0]) +
	( 14'sd 7683) * $signed(input_fmap_201[7:0]) +
	( 13'sd 3658) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12280) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2393) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2078) * $signed(input_fmap_205[7:0]) +
	( 16'sd 17076) * $signed(input_fmap_206[7:0]) +
	( 11'sd 589) * $signed(input_fmap_207[7:0]) +
	( 14'sd 5231) * $signed(input_fmap_208[7:0]) +
	( 15'sd 10703) * $signed(input_fmap_209[7:0]) +
	( 15'sd 13024) * $signed(input_fmap_210[7:0]) +
	( 16'sd 25301) * $signed(input_fmap_211[7:0]) +
	( 16'sd 16683) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3540) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20343) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29877) * $signed(input_fmap_215[7:0]) +
	( 16'sd 16942) * $signed(input_fmap_216[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_217[7:0]) +
	( 15'sd 9431) * $signed(input_fmap_218[7:0]) +
	( 16'sd 23023) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31320) * $signed(input_fmap_220[7:0]) +
	( 15'sd 10440) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25132) * $signed(input_fmap_222[7:0]) +
	( 10'sd 286) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5030) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30675) * $signed(input_fmap_226[7:0]) +
	( 12'sd 2016) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22596) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20864) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14977) * $signed(input_fmap_230[7:0]) +
	( 16'sd 30497) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14444) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10934) * $signed(input_fmap_233[7:0]) +
	( 16'sd 17266) * $signed(input_fmap_234[7:0]) +
	( 16'sd 25418) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23075) * $signed(input_fmap_236[7:0]) +
	( 9'sd 190) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5530) * $signed(input_fmap_238[7:0]) +
	( 14'sd 6774) * $signed(input_fmap_239[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3664) * $signed(input_fmap_241[7:0]) +
	( 16'sd 18861) * $signed(input_fmap_242[7:0]) +
	( 10'sd 376) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19635) * $signed(input_fmap_244[7:0]) +
	( 15'sd 9993) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9568) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13343) * $signed(input_fmap_247[7:0]) +
	( 11'sd 784) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14832) * $signed(input_fmap_249[7:0]) +
	( 16'sd 27134) * $signed(input_fmap_250[7:0]) +
	( 16'sd 25486) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_253[7:0]) +
	( 13'sd 3369) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14717) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_147;
assign conv_mac_147 = 
	( 16'sd 20804) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21589) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6685) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5098) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9027) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1582) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16093) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14686) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12872) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25722) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2547) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23768) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25390) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5301) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14449) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16702) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31504) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4478) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4109) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10268) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12800) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27199) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4555) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18642) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20215) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5284) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16590) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9829) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28689) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3818) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16720) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27384) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26559) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27963) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1173) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14022) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2543) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15281) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16569) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14069) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24390) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25389) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13249) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22677) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19719) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4694) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24012) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30159) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6831) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_51[7:0]) +
	( 16'sd 31360) * $signed(input_fmap_52[7:0]) +
	( 16'sd 26368) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19518) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22114) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16854) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32505) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22500) * $signed(input_fmap_62[7:0]) +
	( 16'sd 31235) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5945) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10281) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7476) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30167) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3543) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2508) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6160) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32295) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8624) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27598) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3872) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1458) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20776) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21608) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28225) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3400) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25985) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25753) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11781) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13816) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25879) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31702) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10671) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21156) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11830) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8577) * $signed(input_fmap_91[7:0]) +
	( 15'sd 8460) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3548) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12346) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_95[7:0]) +
	( 16'sd 26130) * $signed(input_fmap_96[7:0]) +
	( 11'sd 726) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13807) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12806) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10209) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10254) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28154) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19888) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28244) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4836) * $signed(input_fmap_106[7:0]) +
	( 11'sd 713) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25416) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15368) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15617) * $signed(input_fmap_110[7:0]) +
	( 11'sd 899) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13059) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13647) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11743) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5029) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9973) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31071) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12893) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12583) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5637) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1753) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22789) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13182) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28105) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18218) * $signed(input_fmap_127[7:0]) +
	( 16'sd 20788) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31619) * $signed(input_fmap_129[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23977) * $signed(input_fmap_131[7:0]) +
	( 16'sd 23128) * $signed(input_fmap_132[7:0]) +
	( 15'sd 13786) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32444) * $signed(input_fmap_134[7:0]) +
	( 16'sd 24527) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30833) * $signed(input_fmap_136[7:0]) +
	( 16'sd 21659) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_139[7:0]) +
	( 14'sd 5454) * $signed(input_fmap_140[7:0]) +
	( 15'sd 14268) * $signed(input_fmap_141[7:0]) +
	( 16'sd 24251) * $signed(input_fmap_142[7:0]) +
	( 16'sd 19211) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22682) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22896) * $signed(input_fmap_145[7:0]) +
	( 15'sd 13070) * $signed(input_fmap_146[7:0]) +
	( 16'sd 16763) * $signed(input_fmap_147[7:0]) +
	( 16'sd 16498) * $signed(input_fmap_148[7:0]) +
	( 16'sd 19515) * $signed(input_fmap_149[7:0]) +
	( 16'sd 29506) * $signed(input_fmap_150[7:0]) +
	( 15'sd 10676) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_152[7:0]) +
	( 15'sd 13179) * $signed(input_fmap_153[7:0]) +
	( 12'sd 1766) * $signed(input_fmap_154[7:0]) +
	( 13'sd 2283) * $signed(input_fmap_155[7:0]) +
	( 16'sd 26882) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6022) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28653) * $signed(input_fmap_158[7:0]) +
	( 16'sd 16811) * $signed(input_fmap_159[7:0]) +
	( 16'sd 29323) * $signed(input_fmap_160[7:0]) +
	( 14'sd 8144) * $signed(input_fmap_161[7:0]) +
	( 16'sd 25999) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2346) * $signed(input_fmap_163[7:0]) +
	( 16'sd 17413) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4902) * $signed(input_fmap_165[7:0]) +
	( 14'sd 6302) * $signed(input_fmap_166[7:0]) +
	( 15'sd 8308) * $signed(input_fmap_167[7:0]) +
	( 16'sd 30514) * $signed(input_fmap_168[7:0]) +
	( 9'sd 129) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14176) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3836) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15854) * $signed(input_fmap_172[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_173[7:0]) +
	( 16'sd 28119) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21736) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10390) * $signed(input_fmap_176[7:0]) +
	( 15'sd 9656) * $signed(input_fmap_177[7:0]) +
	( 15'sd 12187) * $signed(input_fmap_178[7:0]) +
	( 16'sd 26581) * $signed(input_fmap_179[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_180[7:0]) +
	( 9'sd 194) * $signed(input_fmap_181[7:0]) +
	( 16'sd 25450) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30006) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26866) * $signed(input_fmap_184[7:0]) +
	( 16'sd 16603) * $signed(input_fmap_185[7:0]) +
	( 16'sd 16793) * $signed(input_fmap_186[7:0]) +
	( 16'sd 26901) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32456) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5047) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20297) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20496) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12342) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23425) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22164) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7918) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21214) * $signed(input_fmap_197[7:0]) +
	( 16'sd 23391) * $signed(input_fmap_198[7:0]) +
	( 15'sd 15310) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15164) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27276) * $signed(input_fmap_201[7:0]) +
	( 15'sd 13735) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19439) * $signed(input_fmap_203[7:0]) +
	( 16'sd 26985) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6098) * $signed(input_fmap_205[7:0]) +
	( 15'sd 10838) * $signed(input_fmap_206[7:0]) +
	( 14'sd 6069) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28311) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13176) * $signed(input_fmap_209[7:0]) +
	( 16'sd 32325) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15074) * $signed(input_fmap_211[7:0]) +
	( 14'sd 5699) * $signed(input_fmap_212[7:0]) +
	( 16'sd 30446) * $signed(input_fmap_213[7:0]) +
	( 16'sd 22459) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11625) * $signed(input_fmap_215[7:0]) +
	( 15'sd 13493) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10045) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7455) * $signed(input_fmap_218[7:0]) +
	( 16'sd 29577) * $signed(input_fmap_219[7:0]) +
	( 13'sd 2706) * $signed(input_fmap_220[7:0]) +
	( 13'sd 3199) * $signed(input_fmap_221[7:0]) +
	( 14'sd 6867) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8726) * $signed(input_fmap_223[7:0]) +
	( 16'sd 26533) * $signed(input_fmap_224[7:0]) +
	( 16'sd 23568) * $signed(input_fmap_225[7:0]) +
	( 15'sd 13875) * $signed(input_fmap_226[7:0]) +
	( 16'sd 30232) * $signed(input_fmap_227[7:0]) +
	( 16'sd 28775) * $signed(input_fmap_228[7:0]) +
	( 11'sd 764) * $signed(input_fmap_229[7:0]) +
	( 16'sd 26640) * $signed(input_fmap_230[7:0]) +
	( 13'sd 2706) * $signed(input_fmap_231[7:0]) +
	( 16'sd 22900) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21638) * $signed(input_fmap_233[7:0]) +
	( 13'sd 4094) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22138) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23896) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6008) * $signed(input_fmap_237[7:0]) +
	( 15'sd 10417) * $signed(input_fmap_238[7:0]) +
	( 15'sd 14557) * $signed(input_fmap_239[7:0]) +
	( 15'sd 16153) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26011) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11971) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13445) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24837) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28582) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1857) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12871) * $signed(input_fmap_247[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_248[7:0]) +
	( 14'sd 7379) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25757) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13203) * $signed(input_fmap_251[7:0]) +
	( 16'sd 29051) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28108) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10103) * $signed(input_fmap_254[7:0]) +
	( 13'sd 3098) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_148;
assign conv_mac_148 = 
	( 11'sd 515) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2511) * $signed(input_fmap_1[7:0]) +
	( 14'sd 8054) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14319) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23885) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4382) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3553) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6227) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12108) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11129) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24908) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10595) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18305) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12590) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27843) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18385) * $signed(input_fmap_15[7:0]) +
	( 11'sd 842) * $signed(input_fmap_16[7:0]) +
	( 16'sd 32400) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13988) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30303) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27502) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13876) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26067) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32046) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13722) * $signed(input_fmap_25[7:0]) +
	( 14'sd 6054) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17823) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22123) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14987) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7682) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12343) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3880) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15021) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31020) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2988) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2049) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6553) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25538) * $signed(input_fmap_40[7:0]) +
	( 10'sd 502) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29537) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_44[7:0]) +
	( 11'sd 879) * $signed(input_fmap_45[7:0]) +
	( 7'sd 41) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17612) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29994) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2203) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24305) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13893) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24689) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21278) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21436) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10949) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6037) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20174) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16331) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2379) * $signed(input_fmap_60[7:0]) +
	( 12'sd 1394) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21245) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28073) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23037) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22174) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22693) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12362) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1430) * $signed(input_fmap_69[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1637) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14286) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18784) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19847) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30303) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20530) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11356) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6573) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25705) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27294) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5894) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12246) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27685) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3334) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16066) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32520) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19815) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28692) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28386) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15884) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23478) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_94[7:0]) +
	( 16'sd 17841) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3995) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13107) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4820) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15492) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9643) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21069) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11294) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2583) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12392) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23105) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17293) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17328) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1966) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7312) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8340) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13569) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18138) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21685) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24032) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8971) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20080) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26326) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12677) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28081) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14139) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5359) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2220) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19482) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23048) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2740) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14640) * $signed(input_fmap_130[7:0]) +
	( 16'sd 21333) * $signed(input_fmap_131[7:0]) +
	( 16'sd 32602) * $signed(input_fmap_132[7:0]) +
	( 16'sd 17152) * $signed(input_fmap_133[7:0]) +
	( 16'sd 23105) * $signed(input_fmap_134[7:0]) +
	( 15'sd 13693) * $signed(input_fmap_135[7:0]) +
	( 15'sd 11328) * $signed(input_fmap_136[7:0]) +
	( 16'sd 16532) * $signed(input_fmap_137[7:0]) +
	( 16'sd 24759) * $signed(input_fmap_138[7:0]) +
	( 15'sd 13642) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24094) * $signed(input_fmap_140[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_141[7:0]) +
	( 16'sd 24554) * $signed(input_fmap_142[7:0]) +
	( 15'sd 13136) * $signed(input_fmap_143[7:0]) +
	( 16'sd 32416) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7970) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24132) * $signed(input_fmap_147[7:0]) +
	( 12'sd 1653) * $signed(input_fmap_148[7:0]) +
	( 16'sd 32028) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23285) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28288) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23039) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22984) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27463) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20201) * $signed(input_fmap_156[7:0]) +
	( 16'sd 28274) * $signed(input_fmap_157[7:0]) +
	( 16'sd 32335) * $signed(input_fmap_158[7:0]) +
	( 12'sd 1770) * $signed(input_fmap_159[7:0]) +
	( 15'sd 8621) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31025) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4951) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20405) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6646) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19714) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31152) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30776) * $signed(input_fmap_167[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_168[7:0]) +
	( 14'sd 7460) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_170[7:0]) +
	( 16'sd 25825) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_172[7:0]) +
	( 16'sd 32000) * $signed(input_fmap_173[7:0]) +
	( 14'sd 8076) * $signed(input_fmap_174[7:0]) +
	( 16'sd 22442) * $signed(input_fmap_175[7:0]) +
	( 15'sd 12141) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2878) * $signed(input_fmap_177[7:0]) +
	( 16'sd 21234) * $signed(input_fmap_178[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_179[7:0]) +
	( 16'sd 17645) * $signed(input_fmap_180[7:0]) +
	( 13'sd 2119) * $signed(input_fmap_181[7:0]) +
	( 15'sd 8784) * $signed(input_fmap_182[7:0]) +
	( 16'sd 23754) * $signed(input_fmap_183[7:0]) +
	( 16'sd 17202) * $signed(input_fmap_184[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_185[7:0]) +
	( 16'sd 21717) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28269) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13675) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19074) * $signed(input_fmap_189[7:0]) +
	( 16'sd 21559) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3724) * $signed(input_fmap_191[7:0]) +
	( 15'sd 13889) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27522) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24251) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6840) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10984) * $signed(input_fmap_197[7:0]) +
	( 16'sd 16460) * $signed(input_fmap_198[7:0]) +
	( 16'sd 21107) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26837) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11129) * $signed(input_fmap_201[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_202[7:0]) +
	( 14'sd 7933) * $signed(input_fmap_203[7:0]) +
	( 14'sd 7033) * $signed(input_fmap_204[7:0]) +
	( 16'sd 22296) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28299) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1753) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8834) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11022) * $signed(input_fmap_209[7:0]) +
	( 16'sd 20168) * $signed(input_fmap_210[7:0]) +
	( 16'sd 31123) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29540) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3771) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15057) * $signed(input_fmap_214[7:0]) +
	( 16'sd 21682) * $signed(input_fmap_215[7:0]) +
	( 13'sd 2146) * $signed(input_fmap_216[7:0]) +
	( 15'sd 11073) * $signed(input_fmap_217[7:0]) +
	( 15'sd 11043) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5379) * $signed(input_fmap_219[7:0]) +
	( 16'sd 23836) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19962) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18291) * $signed(input_fmap_222[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_223[7:0]) +
	( 16'sd 24306) * $signed(input_fmap_224[7:0]) +
	( 16'sd 30658) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29112) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22943) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10048) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23273) * $signed(input_fmap_229[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24073) * $signed(input_fmap_231[7:0]) +
	( 15'sd 11205) * $signed(input_fmap_232[7:0]) +
	( 16'sd 19183) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23241) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12562) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2881) * $signed(input_fmap_236[7:0]) +
	( 10'sd 306) * $signed(input_fmap_237[7:0]) +
	( 16'sd 21572) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23816) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10352) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30198) * $signed(input_fmap_241[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23942) * $signed(input_fmap_243[7:0]) +
	( 16'sd 21656) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3957) * $signed(input_fmap_245[7:0]) +
	( 14'sd 6713) * $signed(input_fmap_246[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32424) * $signed(input_fmap_248[7:0]) +
	( 14'sd 6111) * $signed(input_fmap_249[7:0]) +
	( 16'sd 27752) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19563) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4834) * $signed(input_fmap_252[7:0]) +
	( 15'sd 12708) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10910) * $signed(input_fmap_254[7:0]) +
	( 15'sd 13964) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_149;
assign conv_mac_149 = 
	( 16'sd 19013) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31022) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29646) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7409) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28466) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24465) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12950) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10869) * $signed(input_fmap_7[7:0]) +
	( 13'sd 2276) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27019) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15231) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22468) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12730) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31414) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16420) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28840) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7653) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27141) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11389) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27839) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12664) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14271) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7741) * $signed(input_fmap_24[7:0]) +
	( 13'sd 4064) * $signed(input_fmap_25[7:0]) +
	( 16'sd 19837) * $signed(input_fmap_26[7:0]) +
	( 15'sd 16209) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17210) * $signed(input_fmap_28[7:0]) +
	( 14'sd 8063) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19606) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20551) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29451) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28073) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23386) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4342) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11274) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17327) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19367) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21520) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15284) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6157) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24680) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2458) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17876) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22304) * $signed(input_fmap_47[7:0]) +
	( 15'sd 16312) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21889) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28930) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1247) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25801) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2088) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27885) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13154) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1349) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14115) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3693) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19941) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31616) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9051) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14813) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6506) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20009) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12243) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12693) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12210) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10603) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30959) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32582) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25693) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25274) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31393) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29166) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16473) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14039) * $signed(input_fmap_78[7:0]) +
	( 13'sd 4095) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20829) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8422) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14507) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3721) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19436) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3164) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26260) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14157) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3141) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2355) * $signed(input_fmap_90[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_92[7:0]) +
	( 13'sd 2832) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10104) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19631) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24417) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1650) * $signed(input_fmap_98[7:0]) +
	( 14'sd 6262) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25721) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31013) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10544) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12911) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9822) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9467) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17836) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30898) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26713) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20219) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10367) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2522) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7126) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24702) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2624) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13955) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1037) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8308) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19460) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18479) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_120[7:0]) +
	( 16'sd 26468) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14500) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23536) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16925) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9151) * $signed(input_fmap_125[7:0]) +
	( 10'sd 420) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12472) * $signed(input_fmap_127[7:0]) +
	( 15'sd 16219) * $signed(input_fmap_128[7:0]) +
	( 16'sd 18735) * $signed(input_fmap_129[7:0]) +
	( 14'sd 5320) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24147) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25811) * $signed(input_fmap_132[7:0]) +
	( 16'sd 24371) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11284) * $signed(input_fmap_134[7:0]) +
	( 16'sd 17634) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30741) * $signed(input_fmap_136[7:0]) +
	( 16'sd 18381) * $signed(input_fmap_137[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8891) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18433) * $signed(input_fmap_141[7:0]) +
	( 13'sd 2912) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20167) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_144[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_145[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_146[7:0]) +
	( 16'sd 26693) * $signed(input_fmap_147[7:0]) +
	( 15'sd 12484) * $signed(input_fmap_148[7:0]) +
	( 16'sd 22093) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25256) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_151[7:0]) +
	( 15'sd 12768) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4760) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25336) * $signed(input_fmap_154[7:0]) +
	( 16'sd 25378) * $signed(input_fmap_155[7:0]) +
	( 14'sd 5428) * $signed(input_fmap_156[7:0]) +
	( 16'sd 26921) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17770) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14630) * $signed(input_fmap_159[7:0]) +
	( 15'sd 13327) * $signed(input_fmap_160[7:0]) +
	( 16'sd 27013) * $signed(input_fmap_161[7:0]) +
	( 12'sd 1267) * $signed(input_fmap_162[7:0]) +
	( 15'sd 9965) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25705) * $signed(input_fmap_164[7:0]) +
	( 16'sd 21821) * $signed(input_fmap_165[7:0]) +
	( 16'sd 16812) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20890) * $signed(input_fmap_167[7:0]) +
	( 15'sd 10960) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27773) * $signed(input_fmap_169[7:0]) +
	( 15'sd 15784) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19203) * $signed(input_fmap_171[7:0]) +
	( 16'sd 29636) * $signed(input_fmap_172[7:0]) +
	( 11'sd 1023) * $signed(input_fmap_173[7:0]) +
	( 15'sd 15859) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15695) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3309) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2368) * $signed(input_fmap_177[7:0]) +
	( 15'sd 16145) * $signed(input_fmap_178[7:0]) +
	( 15'sd 10805) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_180[7:0]) +
	( 14'sd 7153) * $signed(input_fmap_181[7:0]) +
	( 16'sd 32702) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30293) * $signed(input_fmap_183[7:0]) +
	( 11'sd 753) * $signed(input_fmap_184[7:0]) +
	( 16'sd 16437) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4386) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28543) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1819) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5148) * $signed(input_fmap_189[7:0]) +
	( 13'sd 2997) * $signed(input_fmap_190[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20179) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5908) * $signed(input_fmap_193[7:0]) +
	( 6'sd 23) * $signed(input_fmap_194[7:0]) +
	( 14'sd 4226) * $signed(input_fmap_195[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22052) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5739) * $signed(input_fmap_198[7:0]) +
	( 15'sd 9186) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5978) * $signed(input_fmap_202[7:0]) +
	( 15'sd 11347) * $signed(input_fmap_203[7:0]) +
	( 16'sd 28792) * $signed(input_fmap_204[7:0]) +
	( 15'sd 13410) * $signed(input_fmap_205[7:0]) +
	( 15'sd 10003) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1818) * $signed(input_fmap_207[7:0]) +
	( 13'sd 2503) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3905) * $signed(input_fmap_209[7:0]) +
	( 16'sd 17394) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20553) * $signed(input_fmap_211[7:0]) +
	( 16'sd 25889) * $signed(input_fmap_212[7:0]) +
	( 16'sd 25811) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18700) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6767) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23088) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32608) * $signed(input_fmap_217[7:0]) +
	( 10'sd 460) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21650) * $signed(input_fmap_219[7:0]) +
	( 16'sd 20638) * $signed(input_fmap_220[7:0]) +
	( 16'sd 29370) * $signed(input_fmap_221[7:0]) +
	( 15'sd 8835) * $signed(input_fmap_222[7:0]) +
	( 14'sd 6411) * $signed(input_fmap_223[7:0]) +
	( 15'sd 9204) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18261) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30585) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6154) * $signed(input_fmap_227[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_228[7:0]) +
	( 16'sd 25423) * $signed(input_fmap_229[7:0]) +
	( 16'sd 26678) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3037) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7929) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3190) * $signed(input_fmap_233[7:0]) +
	( 12'sd 1363) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14683) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12865) * $signed(input_fmap_236[7:0]) +
	( 16'sd 25088) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22478) * $signed(input_fmap_238[7:0]) +
	( 14'sd 7829) * $signed(input_fmap_239[7:0]) +
	( 15'sd 16337) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18879) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5657) * $signed(input_fmap_242[7:0]) +
	( 16'sd 27384) * $signed(input_fmap_243[7:0]) +
	( 16'sd 32533) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14624) * $signed(input_fmap_245[7:0]) +
	( 13'sd 2403) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9422) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1918) * $signed(input_fmap_248[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_249[7:0]) +
	( 16'sd 18491) * $signed(input_fmap_250[7:0]) +
	( 13'sd 4080) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17370) * $signed(input_fmap_252[7:0]) +
	( 15'sd 8508) * $signed(input_fmap_253[7:0]) +
	( 16'sd 21971) * $signed(input_fmap_254[7:0]) +
	( 14'sd 4833) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_150;
assign conv_mac_150 = 
	( 16'sd 30870) * $signed(input_fmap_0[7:0]) +
	( 10'sd 256) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5467) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13781) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14539) * $signed(input_fmap_4[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14782) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5542) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11149) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13697) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19109) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2543) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27470) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29058) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6725) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16745) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6456) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19686) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19172) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15648) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18315) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4162) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11013) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17235) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22871) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15263) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25603) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2642) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25086) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1044) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27534) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3148) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28308) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2472) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18156) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17735) * $signed(input_fmap_39[7:0]) +
	( 9'sd 154) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2165) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5031) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9862) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25036) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31436) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4614) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26594) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29869) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17330) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25115) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29324) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3433) * $signed(input_fmap_56[7:0]) +
	( 10'sd 484) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18591) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18361) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4526) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30836) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5521) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24796) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23794) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24029) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25843) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9040) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1701) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20733) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14068) * $signed(input_fmap_72[7:0]) +
	( 16'sd 22895) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11228) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19358) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8078) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1663) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5166) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10404) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20867) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7736) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25400) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1723) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15323) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2265) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8628) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31962) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16609) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13444) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27334) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12159) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3575) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6475) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16820) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25502) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30946) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14366) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18092) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6830) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3141) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4106) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29157) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25466) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7599) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15472) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13892) * $signed(input_fmap_107[7:0]) +
	( 16'sd 31828) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19632) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4677) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18245) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19001) * $signed(input_fmap_112[7:0]) +
	( 11'sd 645) * $signed(input_fmap_113[7:0]) +
	( 8'sd 87) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6728) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10369) * $signed(input_fmap_116[7:0]) +
	( 15'sd 9434) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25263) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2598) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3380) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32623) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1309) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2106) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26517) * $signed(input_fmap_125[7:0]) +
	( 15'sd 16340) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29610) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_128[7:0]) +
	( 16'sd 18096) * $signed(input_fmap_129[7:0]) +
	( 16'sd 26187) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14497) * $signed(input_fmap_131[7:0]) +
	( 16'sd 29589) * $signed(input_fmap_132[7:0]) +
	( 15'sd 8274) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21450) * $signed(input_fmap_134[7:0]) +
	( 16'sd 22354) * $signed(input_fmap_135[7:0]) +
	( 16'sd 32435) * $signed(input_fmap_136[7:0]) +
	( 16'sd 17178) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10905) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28040) * $signed(input_fmap_139[7:0]) +
	( 16'sd 22217) * $signed(input_fmap_140[7:0]) +
	( 16'sd 28137) * $signed(input_fmap_141[7:0]) +
	( 16'sd 29368) * $signed(input_fmap_142[7:0]) +
	( 16'sd 27198) * $signed(input_fmap_143[7:0]) +
	( 16'sd 25808) * $signed(input_fmap_144[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9482) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11926) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3562) * $signed(input_fmap_148[7:0]) +
	( 16'sd 31158) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25512) * $signed(input_fmap_150[7:0]) +
	( 14'sd 8022) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23632) * $signed(input_fmap_152[7:0]) +
	( 16'sd 26221) * $signed(input_fmap_153[7:0]) +
	( 16'sd 21534) * $signed(input_fmap_154[7:0]) +
	( 13'sd 2746) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18320) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22282) * $signed(input_fmap_157[7:0]) +
	( 16'sd 19549) * $signed(input_fmap_158[7:0]) +
	( 14'sd 7289) * $signed(input_fmap_159[7:0]) +
	( 14'sd 4642) * $signed(input_fmap_160[7:0]) +
	( 13'sd 3357) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10807) * $signed(input_fmap_162[7:0]) +
	( 15'sd 13181) * $signed(input_fmap_163[7:0]) +
	( 16'sd 18891) * $signed(input_fmap_164[7:0]) +
	( 11'sd 541) * $signed(input_fmap_165[7:0]) +
	( 13'sd 4054) * $signed(input_fmap_166[7:0]) +
	( 16'sd 22693) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26903) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6099) * $signed(input_fmap_169[7:0]) +
	( 13'sd 3896) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16431) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6843) * $signed(input_fmap_172[7:0]) +
	( 9'sd 157) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16828) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1054) * $signed(input_fmap_175[7:0]) +
	( 16'sd 24655) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_177[7:0]) +
	( 16'sd 18161) * $signed(input_fmap_178[7:0]) +
	( 16'sd 17468) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28800) * $signed(input_fmap_180[7:0]) +
	( 15'sd 12282) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5803) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29132) * $signed(input_fmap_183[7:0]) +
	( 15'sd 12979) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7226) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4245) * $signed(input_fmap_186[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_187[7:0]) +
	( 16'sd 18740) * $signed(input_fmap_188[7:0]) +
	( 16'sd 18968) * $signed(input_fmap_189[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23768) * $signed(input_fmap_191[7:0]) +
	( 13'sd 2998) * $signed(input_fmap_192[7:0]) +
	( 16'sd 23604) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27967) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14911) * $signed(input_fmap_195[7:0]) +
	( 16'sd 32031) * $signed(input_fmap_196[7:0]) +
	( 16'sd 27203) * $signed(input_fmap_197[7:0]) +
	( 16'sd 32177) * $signed(input_fmap_198[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_199[7:0]) +
	( 16'sd 21438) * $signed(input_fmap_200[7:0]) +
	( 16'sd 20237) * $signed(input_fmap_201[7:0]) +
	( 12'sd 1887) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2642) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19290) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18762) * $signed(input_fmap_205[7:0]) +
	( 14'sd 5264) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12315) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24735) * $signed(input_fmap_209[7:0]) +
	( 15'sd 14382) * $signed(input_fmap_210[7:0]) +
	( 16'sd 24153) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17887) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1846) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14263) * $signed(input_fmap_214[7:0]) +
	( 16'sd 31646) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5316) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_217[7:0]) +
	( 11'sd 674) * $signed(input_fmap_218[7:0]) +
	( 14'sd 4598) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19185) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23077) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28325) * $signed(input_fmap_222[7:0]) +
	( 14'sd 7331) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14803) * $signed(input_fmap_224[7:0]) +
	( 16'sd 32739) * $signed(input_fmap_225[7:0]) +
	( 16'sd 24361) * $signed(input_fmap_226[7:0]) +
	( 16'sd 18304) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24517) * $signed(input_fmap_228[7:0]) +
	( 16'sd 22929) * $signed(input_fmap_229[7:0]) +
	( 16'sd 21946) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20930) * $signed(input_fmap_231[7:0]) +
	( 13'sd 2981) * $signed(input_fmap_232[7:0]) +
	( 13'sd 4070) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15792) * $signed(input_fmap_234[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_235[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_236[7:0]) +
	( 16'sd 26041) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14291) * $signed(input_fmap_238[7:0]) +
	( 16'sd 17007) * $signed(input_fmap_239[7:0]) +
	( 13'sd 3219) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25201) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23019) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31321) * $signed(input_fmap_243[7:0]) +
	( 16'sd 31532) * $signed(input_fmap_244[7:0]) +
	( 16'sd 32404) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15936) * $signed(input_fmap_246[7:0]) +
	( 14'sd 6746) * $signed(input_fmap_247[7:0]) +
	( 16'sd 22024) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3084) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9352) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_251[7:0]) +
	( 16'sd 31859) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11143) * $signed(input_fmap_253[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_254[7:0]) +
	( 16'sd 29748) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_151;
assign conv_mac_151 = 
	( 16'sd 20074) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19672) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32582) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29470) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5981) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5953) * $signed(input_fmap_5[7:0]) +
	( 15'sd 16302) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27495) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22276) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11285) * $signed(input_fmap_9[7:0]) +
	( 13'sd 2585) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29964) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15929) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1418) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25176) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22099) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22474) * $signed(input_fmap_18[7:0]) +
	( 10'sd 482) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21456) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23103) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9109) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21940) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20488) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15917) * $signed(input_fmap_25[7:0]) +
	( 15'sd 10715) * $signed(input_fmap_26[7:0]) +
	( 11'sd 932) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20232) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9806) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13229) * $signed(input_fmap_30[7:0]) +
	( 10'sd 427) * $signed(input_fmap_31[7:0]) +
	( 11'sd 609) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29883) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11839) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5425) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13455) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22208) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22989) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3283) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_40[7:0]) +
	( 11'sd 810) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16159) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14361) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6654) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7604) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18281) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24507) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23238) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6793) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32475) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11777) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2378) * $signed(input_fmap_53[7:0]) +
	( 11'sd 835) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10730) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2279) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27586) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7472) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27873) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30135) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3889) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3047) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9275) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23528) * $signed(input_fmap_66[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13712) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24436) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5448) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12385) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6659) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15285) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23973) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22338) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12372) * $signed(input_fmap_76[7:0]) +
	( 16'sd 28987) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27744) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17466) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32049) * $signed(input_fmap_80[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32733) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21625) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19238) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12973) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19583) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32267) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12770) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7680) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29968) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31164) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11237) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15852) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5836) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15086) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11554) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16462) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3612) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27902) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1317) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20454) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1406) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19864) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32681) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12417) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_111[7:0]) +
	( 16'sd 20664) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3742) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17069) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12999) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22329) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21780) * $signed(input_fmap_117[7:0]) +
	( 16'sd 19643) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3832) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_120[7:0]) +
	( 15'sd 11843) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19633) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6160) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22406) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10107) * $signed(input_fmap_127[7:0]) +
	( 12'sd 1523) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_129[7:0]) +
	( 13'sd 3595) * $signed(input_fmap_130[7:0]) +
	( 16'sd 25790) * $signed(input_fmap_131[7:0]) +
	( 16'sd 32224) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19130) * $signed(input_fmap_135[7:0]) +
	( 15'sd 11502) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13718) * $signed(input_fmap_137[7:0]) +
	( 8'sd 120) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31767) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9650) * $signed(input_fmap_140[7:0]) +
	( 16'sd 28910) * $signed(input_fmap_141[7:0]) +
	( 16'sd 16947) * $signed(input_fmap_142[7:0]) +
	( 16'sd 27980) * $signed(input_fmap_143[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_144[7:0]) +
	( 16'sd 30349) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9375) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29355) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21501) * $signed(input_fmap_148[7:0]) +
	( 16'sd 29384) * $signed(input_fmap_149[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_150[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_151[7:0]) +
	( 16'sd 17889) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14949) * $signed(input_fmap_153[7:0]) +
	( 12'sd 1391) * $signed(input_fmap_154[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_155[7:0]) +
	( 16'sd 26740) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22154) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18593) * $signed(input_fmap_158[7:0]) +
	( 12'sd 1670) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11199) * $signed(input_fmap_160[7:0]) +
	( 15'sd 12604) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26418) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26137) * $signed(input_fmap_163[7:0]) +
	( 16'sd 28122) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9163) * $signed(input_fmap_166[7:0]) +
	( 15'sd 15697) * $signed(input_fmap_167[7:0]) +
	( 16'sd 30800) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20553) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30073) * $signed(input_fmap_171[7:0]) +
	( 16'sd 29663) * $signed(input_fmap_172[7:0]) +
	( 16'sd 16523) * $signed(input_fmap_173[7:0]) +
	( 14'sd 5262) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4633) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10829) * $signed(input_fmap_176[7:0]) +
	( 16'sd 20367) * $signed(input_fmap_177[7:0]) +
	( 16'sd 20976) * $signed(input_fmap_178[7:0]) +
	( 14'sd 8184) * $signed(input_fmap_179[7:0]) +
	( 12'sd 1104) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3959) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4261) * $signed(input_fmap_182[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11174) * $signed(input_fmap_184[7:0]) +
	( 15'sd 9092) * $signed(input_fmap_185[7:0]) +
	( 15'sd 15132) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30555) * $signed(input_fmap_189[7:0]) +
	( 13'sd 3708) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29790) * $signed(input_fmap_191[7:0]) +
	( 16'sd 18470) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26195) * $signed(input_fmap_193[7:0]) +
	( 16'sd 19928) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14469) * $signed(input_fmap_195[7:0]) +
	( 13'sd 4049) * $signed(input_fmap_196[7:0]) +
	( 16'sd 27618) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19036) * $signed(input_fmap_198[7:0]) +
	( 11'sd 521) * $signed(input_fmap_199[7:0]) +
	( 13'sd 2312) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22978) * $signed(input_fmap_201[7:0]) +
	( 15'sd 15196) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24638) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15562) * $signed(input_fmap_204[7:0]) +
	( 15'sd 10505) * $signed(input_fmap_205[7:0]) +
	( 16'sd 19494) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5630) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22805) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22761) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10375) * $signed(input_fmap_210[7:0]) +
	( 16'sd 18709) * $signed(input_fmap_211[7:0]) +
	( 13'sd 3827) * $signed(input_fmap_212[7:0]) +
	( 16'sd 16802) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23193) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_215[7:0]) +
	( 15'sd 12955) * $signed(input_fmap_216[7:0]) +
	( 14'sd 6065) * $signed(input_fmap_217[7:0]) +
	( 16'sd 27151) * $signed(input_fmap_218[7:0]) +
	( 16'sd 25692) * $signed(input_fmap_219[7:0]) +
	( 15'sd 16070) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5069) * $signed(input_fmap_221[7:0]) +
	( 16'sd 26133) * $signed(input_fmap_222[7:0]) +
	( 14'sd 5839) * $signed(input_fmap_223[7:0]) +
	( 16'sd 31098) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18542) * $signed(input_fmap_225[7:0]) +
	( 16'sd 25880) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_227[7:0]) +
	( 15'sd 11654) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8538) * $signed(input_fmap_229[7:0]) +
	( 14'sd 5187) * $signed(input_fmap_230[7:0]) +
	( 16'sd 22020) * $signed(input_fmap_231[7:0]) +
	( 14'sd 5901) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_233[7:0]) +
	( 16'sd 32559) * $signed(input_fmap_234[7:0]) +
	( 15'sd 10633) * $signed(input_fmap_235[7:0]) +
	( 15'sd 14076) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6759) * $signed(input_fmap_237[7:0]) +
	( 14'sd 6735) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5462) * $signed(input_fmap_239[7:0]) +
	( 16'sd 27941) * $signed(input_fmap_240[7:0]) +
	( 15'sd 9953) * $signed(input_fmap_241[7:0]) +
	( 16'sd 22586) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13102) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28957) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28515) * $signed(input_fmap_245[7:0]) +
	( 14'sd 6037) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20013) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1538) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2704) * $signed(input_fmap_249[7:0]) +
	( 16'sd 19833) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12720) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17242) * $signed(input_fmap_252[7:0]) +
	( 14'sd 4226) * $signed(input_fmap_253[7:0]) +
	( 15'sd 11802) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23700) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_152;
assign conv_mac_152 = 
	( 16'sd 16635) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28690) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6636) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32414) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12068) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23495) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25280) * $signed(input_fmap_7[7:0]) +
	( 6'sd 18) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12038) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19426) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21426) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25599) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28062) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3612) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18596) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11651) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21065) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21475) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15448) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26936) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13750) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20015) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31354) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27432) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27314) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16638) * $signed(input_fmap_29[7:0]) +
	( 15'sd 11219) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23324) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16551) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13333) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24538) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2492) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30222) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2204) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17338) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12358) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3159) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29603) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27965) * $signed(input_fmap_43[7:0]) +
	( 15'sd 14318) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27179) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3288) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9415) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21729) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21417) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2187) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25027) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27725) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19859) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9477) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1643) * $signed(input_fmap_57[7:0]) +
	( 14'sd 8039) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26598) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14319) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8384) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23655) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23633) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17583) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25611) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29331) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18730) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13197) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_70[7:0]) +
	( 14'sd 8037) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21959) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6020) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30638) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5818) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23705) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12046) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12420) * $signed(input_fmap_78[7:0]) +
	( 16'sd 32256) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19558) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27036) * $signed(input_fmap_81[7:0]) +
	( 13'sd 4036) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10485) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4992) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9251) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31888) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21524) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14440) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15331) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16401) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12698) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16711) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28417) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23866) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11520) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25050) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9797) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3082) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21892) * $signed(input_fmap_104[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30084) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32090) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6742) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30576) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22996) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25196) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7196) * $signed(input_fmap_113[7:0]) +
	( 11'sd 803) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15346) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26707) * $signed(input_fmap_116[7:0]) +
	( 12'sd 2008) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14272) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20559) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30812) * $signed(input_fmap_120[7:0]) +
	( 13'sd 2386) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29326) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8317) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10379) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27644) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18743) * $signed(input_fmap_126[7:0]) +
	( 11'sd 709) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13034) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24787) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10470) * $signed(input_fmap_130[7:0]) +
	( 12'sd 1721) * $signed(input_fmap_131[7:0]) +
	( 16'sd 21296) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10060) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2649) * $signed(input_fmap_134[7:0]) +
	( 15'sd 8580) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1612) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25248) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11533) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28326) * $signed(input_fmap_139[7:0]) +
	( 16'sd 20226) * $signed(input_fmap_140[7:0]) +
	( 15'sd 8405) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21880) * $signed(input_fmap_142[7:0]) +
	( 16'sd 19668) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31815) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2085) * $signed(input_fmap_145[7:0]) +
	( 16'sd 17517) * $signed(input_fmap_146[7:0]) +
	( 12'sd 1721) * $signed(input_fmap_147[7:0]) +
	( 16'sd 16883) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23018) * $signed(input_fmap_149[7:0]) +
	( 16'sd 28207) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14835) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23043) * $signed(input_fmap_152[7:0]) +
	( 16'sd 30916) * $signed(input_fmap_153[7:0]) +
	( 15'sd 9851) * $signed(input_fmap_154[7:0]) +
	( 16'sd 24790) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14871) * $signed(input_fmap_156[7:0]) +
	( 16'sd 32208) * $signed(input_fmap_157[7:0]) +
	( 13'sd 2435) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_159[7:0]) +
	( 12'sd 1998) * $signed(input_fmap_160[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_161[7:0]) +
	( 12'sd 1730) * $signed(input_fmap_162[7:0]) +
	( 15'sd 14228) * $signed(input_fmap_163[7:0]) +
	( 8'sd 91) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14646) * $signed(input_fmap_165[7:0]) +
	( 16'sd 21225) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13561) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6031) * $signed(input_fmap_168[7:0]) +
	( 16'sd 23461) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24183) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7214) * $signed(input_fmap_171[7:0]) +
	( 16'sd 24605) * $signed(input_fmap_172[7:0]) +
	( 16'sd 25846) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32320) * $signed(input_fmap_174[7:0]) +
	( 16'sd 27558) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27737) * $signed(input_fmap_176[7:0]) +
	( 16'sd 17584) * $signed(input_fmap_177[7:0]) +
	( 15'sd 13307) * $signed(input_fmap_178[7:0]) +
	( 15'sd 13003) * $signed(input_fmap_179[7:0]) +
	( 15'sd 10870) * $signed(input_fmap_180[7:0]) +
	( 14'sd 7757) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5097) * $signed(input_fmap_182[7:0]) +
	( 15'sd 8537) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22567) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27895) * $signed(input_fmap_185[7:0]) +
	( 16'sd 30996) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25192) * $signed(input_fmap_187[7:0]) +
	( 15'sd 10429) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26166) * $signed(input_fmap_189[7:0]) +
	( 15'sd 15878) * $signed(input_fmap_190[7:0]) +
	( 15'sd 12205) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22394) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30789) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12788) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15592) * $signed(input_fmap_196[7:0]) +
	( 15'sd 8212) * $signed(input_fmap_197[7:0]) +
	( 16'sd 16619) * $signed(input_fmap_198[7:0]) +
	( 16'sd 31803) * $signed(input_fmap_199[7:0]) +
	( 16'sd 16432) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1396) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21465) * $signed(input_fmap_202[7:0]) +
	( 15'sd 8448) * $signed(input_fmap_203[7:0]) +
	( 7'sd 57) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15789) * $signed(input_fmap_205[7:0]) +
	( 14'sd 7291) * $signed(input_fmap_206[7:0]) +
	( 16'sd 22331) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6779) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24656) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23473) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23738) * $signed(input_fmap_211[7:0]) +
	( 15'sd 15189) * $signed(input_fmap_212[7:0]) +
	( 16'sd 20989) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28604) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1449) * $signed(input_fmap_215[7:0]) +
	( 16'sd 29311) * $signed(input_fmap_216[7:0]) +
	( 16'sd 27079) * $signed(input_fmap_217[7:0]) +
	( 13'sd 3649) * $signed(input_fmap_218[7:0]) +
	( 16'sd 18607) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25836) * $signed(input_fmap_220[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_221[7:0]) +
	( 8'sd 106) * $signed(input_fmap_222[7:0]) +
	( 16'sd 21193) * $signed(input_fmap_223[7:0]) +
	( 15'sd 10146) * $signed(input_fmap_224[7:0]) +
	( 15'sd 12816) * $signed(input_fmap_225[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_226[7:0]) +
	( 16'sd 19139) * $signed(input_fmap_227[7:0]) +
	( 16'sd 21496) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_229[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31880) * $signed(input_fmap_231[7:0]) +
	( 16'sd 23152) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23991) * $signed(input_fmap_233[7:0]) +
	( 14'sd 6593) * $signed(input_fmap_234[7:0]) +
	( 15'sd 9084) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30918) * $signed(input_fmap_236[7:0]) +
	( 15'sd 13017) * $signed(input_fmap_237[7:0]) +
	( 15'sd 9570) * $signed(input_fmap_238[7:0]) +
	( 11'sd 1006) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1953) * $signed(input_fmap_240[7:0]) +
	( 15'sd 16305) * $signed(input_fmap_241[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_242[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_243[7:0]) +
	( 15'sd 8500) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22889) * $signed(input_fmap_245[7:0]) +
	( 16'sd 25792) * $signed(input_fmap_246[7:0]) +
	( 12'sd 1578) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21101) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21623) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26828) * $signed(input_fmap_250[7:0]) +
	( 15'sd 9024) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29078) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_254[7:0]) +
	( 11'sd 916) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_153;
assign conv_mac_153 = 
	( 16'sd 20258) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29647) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2118) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16948) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26848) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32106) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6552) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17726) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11974) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14047) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5720) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21054) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29743) * $signed(input_fmap_12[7:0]) +
	( 15'sd 16298) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10399) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10823) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2840) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28278) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22591) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18332) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32695) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14471) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23133) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_23[7:0]) +
	( 16'sd 19228) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30024) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12549) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24218) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30547) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32712) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21480) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20946) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29058) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16947) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16995) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6687) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7423) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30559) * $signed(input_fmap_38[7:0]) +
	( 12'sd 2033) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23964) * $signed(input_fmap_40[7:0]) +
	( 16'sd 29187) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12631) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3076) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27925) * $signed(input_fmap_44[7:0]) +
	( 14'sd 5349) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19941) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22339) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29940) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6106) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27045) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22179) * $signed(input_fmap_53[7:0]) +
	( 16'sd 20264) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18274) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22127) * $signed(input_fmap_56[7:0]) +
	( 10'sd 352) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24364) * $signed(input_fmap_58[7:0]) +
	( 11'sd 868) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6710) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27607) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_62[7:0]) +
	( 11'sd 1005) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24363) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6053) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11762) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5931) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3003) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2372) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29622) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29273) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29017) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8479) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21426) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1956) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29375) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30750) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25780) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10047) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3332) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20802) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21661) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26899) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4426) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2591) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24959) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19305) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2666) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11777) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22015) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30540) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5511) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18134) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19267) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22989) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30682) * $signed(input_fmap_99[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24105) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29059) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16823) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31527) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4929) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10686) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21615) * $signed(input_fmap_107[7:0]) +
	( 15'sd 11855) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17935) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18891) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4644) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17384) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30072) * $signed(input_fmap_114[7:0]) +
	( 16'sd 22176) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3264) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18106) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31608) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12792) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17461) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26857) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30415) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9360) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7967) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2519) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18463) * $signed(input_fmap_128[7:0]) +
	( 16'sd 26101) * $signed(input_fmap_129[7:0]) +
	( 15'sd 13592) * $signed(input_fmap_130[7:0]) +
	( 16'sd 18695) * $signed(input_fmap_131[7:0]) +
	( 16'sd 28825) * $signed(input_fmap_132[7:0]) +
	( 12'sd 1949) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18874) * $signed(input_fmap_134[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12618) * $signed(input_fmap_136[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19232) * $signed(input_fmap_138[7:0]) +
	( 14'sd 4733) * $signed(input_fmap_139[7:0]) +
	( 16'sd 22994) * $signed(input_fmap_140[7:0]) +
	( 16'sd 28213) * $signed(input_fmap_141[7:0]) +
	( 15'sd 13322) * $signed(input_fmap_142[7:0]) +
	( 15'sd 14995) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19738) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17846) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14139) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9018) * $signed(input_fmap_147[7:0]) +
	( 15'sd 9311) * $signed(input_fmap_148[7:0]) +
	( 12'sd 1801) * $signed(input_fmap_149[7:0]) +
	( 15'sd 8738) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30993) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20153) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25244) * $signed(input_fmap_153[7:0]) +
	( 13'sd 2838) * $signed(input_fmap_154[7:0]) +
	( 16'sd 17876) * $signed(input_fmap_155[7:0]) +
	( 16'sd 23803) * $signed(input_fmap_156[7:0]) +
	( 15'sd 16130) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1133) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2484) * $signed(input_fmap_159[7:0]) +
	( 13'sd 2816) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31804) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27603) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26567) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3619) * $signed(input_fmap_164[7:0]) +
	( 16'sd 27843) * $signed(input_fmap_165[7:0]) +
	( 15'sd 15145) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30940) * $signed(input_fmap_167[7:0]) +
	( 13'sd 3716) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26876) * $signed(input_fmap_169[7:0]) +
	( 16'sd 32585) * $signed(input_fmap_170[7:0]) +
	( 16'sd 22044) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7538) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12858) * $signed(input_fmap_173[7:0]) +
	( 15'sd 16058) * $signed(input_fmap_174[7:0]) +
	( 16'sd 19144) * $signed(input_fmap_175[7:0]) +
	( 16'sd 30859) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5403) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2445) * $signed(input_fmap_179[7:0]) +
	( 14'sd 7508) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11370) * $signed(input_fmap_181[7:0]) +
	( 15'sd 8480) * $signed(input_fmap_182[7:0]) +
	( 16'sd 31637) * $signed(input_fmap_183[7:0]) +
	( 16'sd 16711) * $signed(input_fmap_184[7:0]) +
	( 10'sd 386) * $signed(input_fmap_185[7:0]) +
	( 16'sd 29227) * $signed(input_fmap_186[7:0]) +
	( 16'sd 23207) * $signed(input_fmap_187[7:0]) +
	( 16'sd 27149) * $signed(input_fmap_188[7:0]) +
	( 15'sd 14065) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13551) * $signed(input_fmap_190[7:0]) +
	( 11'sd 682) * $signed(input_fmap_191[7:0]) +
	( 16'sd 30687) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28118) * $signed(input_fmap_193[7:0]) +
	( 16'sd 17588) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17115) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17257) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21171) * $signed(input_fmap_197[7:0]) +
	( 7'sd 53) * $signed(input_fmap_198[7:0]) +
	( 10'sd 267) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6180) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18660) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12979) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4571) * $signed(input_fmap_204[7:0]) +
	( 15'sd 8752) * $signed(input_fmap_205[7:0]) +
	( 16'sd 26926) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5292) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11283) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19534) * $signed(input_fmap_210[7:0]) +
	( 16'sd 22624) * $signed(input_fmap_211[7:0]) +
	( 13'sd 3565) * $signed(input_fmap_212[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_213[7:0]) +
	( 13'sd 3649) * $signed(input_fmap_214[7:0]) +
	( 16'sd 21269) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4440) * $signed(input_fmap_216[7:0]) +
	( 16'sd 20637) * $signed(input_fmap_217[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_218[7:0]) +
	( 14'sd 7932) * $signed(input_fmap_219[7:0]) +
	( 16'sd 29630) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13533) * $signed(input_fmap_221[7:0]) +
	( 16'sd 17326) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2940) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30503) * $signed(input_fmap_224[7:0]) +
	( 15'sd 11739) * $signed(input_fmap_225[7:0]) +
	( 16'sd 20244) * $signed(input_fmap_226[7:0]) +
	( 16'sd 19463) * $signed(input_fmap_227[7:0]) +
	( 16'sd 32132) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10549) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18729) * $signed(input_fmap_230[7:0]) +
	( 15'sd 9099) * $signed(input_fmap_231[7:0]) +
	( 13'sd 3233) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15208) * $signed(input_fmap_233[7:0]) +
	( 11'sd 582) * $signed(input_fmap_234[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5726) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29610) * $signed(input_fmap_237[7:0]) +
	( 12'sd 1245) * $signed(input_fmap_238[7:0]) +
	( 16'sd 25140) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19496) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21416) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15633) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2563) * $signed(input_fmap_243[7:0]) +
	( 16'sd 25598) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3421) * $signed(input_fmap_245[7:0]) +
	( 14'sd 7493) * $signed(input_fmap_246[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_247[7:0]) +
	( 11'sd 966) * $signed(input_fmap_248[7:0]) +
	( 16'sd 29278) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30692) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19713) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26987) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_253[7:0]) +
	( 16'sd 29238) * $signed(input_fmap_254[7:0]) +
	( 16'sd 22950) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_154;
assign conv_mac_154 = 
	( 15'sd 9197) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32439) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21985) * $signed(input_fmap_2[7:0]) +
	( 11'sd 512) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21045) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22144) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31461) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8678) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_8[7:0]) +
	( 16'sd 19748) * $signed(input_fmap_9[7:0]) +
	( 16'sd 22324) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13480) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23247) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7352) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5349) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20447) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32125) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22512) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7728) * $signed(input_fmap_19[7:0]) +
	( 16'sd 21133) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24852) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24819) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22523) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7686) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3682) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27957) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1212) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19485) * $signed(input_fmap_28[7:0]) +
	( 16'sd 20050) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23524) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10366) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8942) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32012) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13698) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24237) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27040) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18302) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9548) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7000) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9491) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27481) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11580) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6576) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19326) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25335) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24779) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31540) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4141) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22201) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23525) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31000) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11269) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15538) * $signed(input_fmap_58[7:0]) +
	( 14'sd 8059) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7394) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13878) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31728) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26822) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24585) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27573) * $signed(input_fmap_65[7:0]) +
	( 11'sd 904) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12411) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25220) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32331) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11056) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21144) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27932) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24335) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11440) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3081) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20306) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2555) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4557) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8786) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7462) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29193) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14406) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12758) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27141) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25423) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27522) * $signed(input_fmap_87[7:0]) +
	( 16'sd 29130) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23459) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22557) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13779) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15334) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24058) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14033) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15632) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8503) * $signed(input_fmap_97[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23937) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10275) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12271) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23326) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29170) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23534) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12242) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11828) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10920) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30621) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6937) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4903) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_112[7:0]) +
	( 14'sd 6438) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21677) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17459) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26297) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4334) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3755) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14834) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20940) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5815) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12016) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26257) * $signed(input_fmap_123[7:0]) +
	( 8'sd 85) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12873) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14772) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_127[7:0]) +
	( 16'sd 25412) * $signed(input_fmap_128[7:0]) +
	( 16'sd 21047) * $signed(input_fmap_129[7:0]) +
	( 13'sd 2613) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31240) * $signed(input_fmap_131[7:0]) +
	( 11'sd 856) * $signed(input_fmap_132[7:0]) +
	( 14'sd 7078) * $signed(input_fmap_133[7:0]) +
	( 16'sd 21531) * $signed(input_fmap_134[7:0]) +
	( 15'sd 12782) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17138) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6700) * $signed(input_fmap_137[7:0]) +
	( 14'sd 8061) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11940) * $signed(input_fmap_139[7:0]) +
	( 16'sd 16737) * $signed(input_fmap_140[7:0]) +
	( 14'sd 6993) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1385) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11327) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28194) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14046) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23839) * $signed(input_fmap_148[7:0]) +
	( 11'sd 665) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15658) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14380) * $signed(input_fmap_151[7:0]) +
	( 16'sd 26202) * $signed(input_fmap_152[7:0]) +
	( 16'sd 22381) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22060) * $signed(input_fmap_154[7:0]) +
	( 16'sd 16534) * $signed(input_fmap_155[7:0]) +
	( 15'sd 12392) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18616) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1855) * $signed(input_fmap_158[7:0]) +
	( 16'sd 22651) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26950) * $signed(input_fmap_160[7:0]) +
	( 16'sd 27162) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21148) * $signed(input_fmap_162[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_163[7:0]) +
	( 15'sd 14398) * $signed(input_fmap_164[7:0]) +
	( 10'sd 470) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19971) * $signed(input_fmap_166[7:0]) +
	( 9'sd 194) * $signed(input_fmap_167[7:0]) +
	( 16'sd 30331) * $signed(input_fmap_168[7:0]) +
	( 15'sd 13808) * $signed(input_fmap_169[7:0]) +
	( 16'sd 21984) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11186) * $signed(input_fmap_171[7:0]) +
	( 9'sd 157) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27301) * $signed(input_fmap_173[7:0]) +
	( 16'sd 20908) * $signed(input_fmap_174[7:0]) +
	( 16'sd 20581) * $signed(input_fmap_175[7:0]) +
	( 9'sd 217) * $signed(input_fmap_176[7:0]) +
	( 16'sd 23289) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9090) * $signed(input_fmap_178[7:0]) +
	( 14'sd 4446) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29887) * $signed(input_fmap_180[7:0]) +
	( 12'sd 1076) * $signed(input_fmap_181[7:0]) +
	( 15'sd 13510) * $signed(input_fmap_182[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9364) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_185[7:0]) +
	( 14'sd 7291) * $signed(input_fmap_186[7:0]) +
	( 16'sd 17380) * $signed(input_fmap_187[7:0]) +
	( 16'sd 24687) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7004) * $signed(input_fmap_189[7:0]) +
	( 16'sd 18045) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17915) * $signed(input_fmap_191[7:0]) +
	( 15'sd 9007) * $signed(input_fmap_192[7:0]) +
	( 16'sd 31647) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26643) * $signed(input_fmap_194[7:0]) +
	( 16'sd 30911) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11469) * $signed(input_fmap_196[7:0]) +
	( 16'sd 29658) * $signed(input_fmap_197[7:0]) +
	( 16'sd 28862) * $signed(input_fmap_198[7:0]) +
	( 15'sd 9239) * $signed(input_fmap_199[7:0]) +
	( 14'sd 4802) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6641) * $signed(input_fmap_201[7:0]) +
	( 15'sd 13416) * $signed(input_fmap_202[7:0]) +
	( 12'sd 1043) * $signed(input_fmap_203[7:0]) +
	( 16'sd 29850) * $signed(input_fmap_204[7:0]) +
	( 14'sd 4856) * $signed(input_fmap_205[7:0]) +
	( 16'sd 23112) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17132) * $signed(input_fmap_207[7:0]) +
	( 16'sd 31268) * $signed(input_fmap_208[7:0]) +
	( 16'sd 29440) * $signed(input_fmap_209[7:0]) +
	( 14'sd 8031) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3975) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14029) * $signed(input_fmap_212[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_214[7:0]) +
	( 16'sd 24128) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5554) * $signed(input_fmap_216[7:0]) +
	( 11'sd 766) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30316) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3953) * $signed(input_fmap_219[7:0]) +
	( 15'sd 16096) * $signed(input_fmap_220[7:0]) +
	( 16'sd 24549) * $signed(input_fmap_221[7:0]) +
	( 10'sd 373) * $signed(input_fmap_222[7:0]) +
	( 14'sd 4307) * $signed(input_fmap_223[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27975) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7063) * $signed(input_fmap_226[7:0]) +
	( 16'sd 21462) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19637) * $signed(input_fmap_228[7:0]) +
	( 16'sd 27761) * $signed(input_fmap_229[7:0]) +
	( 15'sd 11849) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28100) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18170) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28794) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5121) * $signed(input_fmap_234[7:0]) +
	( 16'sd 28228) * $signed(input_fmap_235[7:0]) +
	( 15'sd 9138) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29468) * $signed(input_fmap_237[7:0]) +
	( 14'sd 6102) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_239[7:0]) +
	( 15'sd 12781) * $signed(input_fmap_240[7:0]) +
	( 15'sd 12182) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29224) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22313) * $signed(input_fmap_243[7:0]) +
	( 14'sd 4454) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6235) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9053) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30288) * $signed(input_fmap_247[7:0]) +
	( 14'sd 6829) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21427) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22916) * $signed(input_fmap_250[7:0]) +
	( 16'sd 28254) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6510) * $signed(input_fmap_252[7:0]) +
	( 16'sd 16663) * $signed(input_fmap_253[7:0]) +
	( 15'sd 16193) * $signed(input_fmap_254[7:0]) +
	( 12'sd 1095) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_155;
assign conv_mac_155 = 
	( 16'sd 27921) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9135) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6892) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3270) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30040) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2729) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27067) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16249) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27526) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18579) * $signed(input_fmap_10[7:0]) +
	( 15'sd 13986) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13440) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6005) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13502) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13944) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23846) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13681) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6398) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4496) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20949) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1348) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5279) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25783) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11195) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21265) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9164) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25115) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7764) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29295) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16504) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31624) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28435) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30176) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15549) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25990) * $signed(input_fmap_36[7:0]) +
	( 11'sd 864) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21753) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8426) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17294) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6558) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23289) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19167) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27043) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7862) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17744) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5311) * $signed(input_fmap_48[7:0]) +
	( 14'sd 4779) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25666) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12307) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27829) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7117) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30679) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11955) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4496) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16896) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25461) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3349) * $signed(input_fmap_60[7:0]) +
	( 14'sd 5868) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32477) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4978) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20009) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32493) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12427) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5482) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25603) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28337) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27202) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19866) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30531) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29727) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16847) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1150) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17546) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29080) * $signed(input_fmap_78[7:0]) +
	( 11'sd 522) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9686) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29325) * $signed(input_fmap_81[7:0]) +
	( 16'sd 31848) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1266) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19110) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1710) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21892) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4217) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32517) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4349) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28467) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6766) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19375) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19691) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4112) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23854) * $signed(input_fmap_95[7:0]) +
	( 10'sd 372) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13539) * $signed(input_fmap_97[7:0]) +
	( 15'sd 16259) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21694) * $signed(input_fmap_99[7:0]) +
	( 16'sd 25220) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10138) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23534) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22999) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7947) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1483) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7734) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7749) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25346) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5895) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25365) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8280) * $signed(input_fmap_112[7:0]) +
	( 16'sd 16823) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_114[7:0]) +
	( 14'sd 7494) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26549) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18900) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29964) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4728) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14249) * $signed(input_fmap_122[7:0]) +
	( 16'sd 31331) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29897) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20338) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19768) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2449) * $signed(input_fmap_127[7:0]) +
	( 12'sd 1553) * $signed(input_fmap_128[7:0]) +
	( 15'sd 8857) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27079) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13925) * $signed(input_fmap_131[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_132[7:0]) +
	( 16'sd 26030) * $signed(input_fmap_133[7:0]) +
	( 15'sd 8945) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10557) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4146) * $signed(input_fmap_136[7:0]) +
	( 15'sd 8279) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_138[7:0]) +
	( 14'sd 4513) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1323) * $signed(input_fmap_140[7:0]) +
	( 11'sd 717) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12274) * $signed(input_fmap_143[7:0]) +
	( 16'sd 27576) * $signed(input_fmap_144[7:0]) +
	( 16'sd 16444) * $signed(input_fmap_145[7:0]) +
	( 16'sd 17009) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24355) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_148[7:0]) +
	( 15'sd 8866) * $signed(input_fmap_149[7:0]) +
	( 15'sd 14241) * $signed(input_fmap_150[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_151[7:0]) +
	( 16'sd 25179) * $signed(input_fmap_152[7:0]) +
	( 14'sd 7316) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31647) * $signed(input_fmap_154[7:0]) +
	( 14'sd 6017) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14123) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5737) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32155) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22729) * $signed(input_fmap_160[7:0]) +
	( 11'sd 862) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10085) * $signed(input_fmap_162[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9673) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23606) * $signed(input_fmap_165[7:0]) +
	( 14'sd 7127) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23043) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4285) * $signed(input_fmap_168[7:0]) +
	( 14'sd 4953) * $signed(input_fmap_169[7:0]) +
	( 16'sd 30016) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12922) * $signed(input_fmap_171[7:0]) +
	( 15'sd 8561) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19504) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14053) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10782) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18427) * $signed(input_fmap_177[7:0]) +
	( 16'sd 20589) * $signed(input_fmap_178[7:0]) +
	( 15'sd 9977) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24058) * $signed(input_fmap_180[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_181[7:0]) +
	( 16'sd 18782) * $signed(input_fmap_182[7:0]) +
	( 14'sd 4269) * $signed(input_fmap_183[7:0]) +
	( 16'sd 23671) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7944) * $signed(input_fmap_185[7:0]) +
	( 16'sd 19973) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2977) * $signed(input_fmap_187[7:0]) +
	( 16'sd 16457) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26348) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9012) * $signed(input_fmap_190[7:0]) +
	( 13'sd 2561) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20375) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5322) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29492) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5229) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19584) * $signed(input_fmap_197[7:0]) +
	( 16'sd 17667) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14393) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26087) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_202[7:0]) +
	( 16'sd 32586) * $signed(input_fmap_203[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_204[7:0]) +
	( 15'sd 16005) * $signed(input_fmap_205[7:0]) +
	( 16'sd 18925) * $signed(input_fmap_206[7:0]) +
	( 16'sd 27097) * $signed(input_fmap_207[7:0]) +
	( 16'sd 19217) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20110) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1165) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12872) * $signed(input_fmap_211[7:0]) +
	( 10'sd 336) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12598) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20923) * $signed(input_fmap_214[7:0]) +
	( 14'sd 8152) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28490) * $signed(input_fmap_216[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5752) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19521) * $signed(input_fmap_220[7:0]) +
	( 15'sd 14262) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_222[7:0]) +
	( 13'sd 3214) * $signed(input_fmap_223[7:0]) +
	( 14'sd 4548) * $signed(input_fmap_224[7:0]) +
	( 15'sd 12838) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_226[7:0]) +
	( 16'sd 23609) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4798) * $signed(input_fmap_228[7:0]) +
	( 15'sd 14165) * $signed(input_fmap_229[7:0]) +
	( 14'sd 5171) * $signed(input_fmap_230[7:0]) +
	( 16'sd 19841) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15979) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24554) * $signed(input_fmap_233[7:0]) +
	( 16'sd 22028) * $signed(input_fmap_234[7:0]) +
	( 15'sd 8533) * $signed(input_fmap_235[7:0]) +
	( 12'sd 2043) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11154) * $signed(input_fmap_237[7:0]) +
	( 15'sd 9001) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23771) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26734) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_241[7:0]) +
	( 16'sd 30813) * $signed(input_fmap_242[7:0]) +
	( 15'sd 14486) * $signed(input_fmap_243[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_244[7:0]) +
	( 15'sd 13754) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30273) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3717) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18356) * $signed(input_fmap_248[7:0]) +
	( 15'sd 8742) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24093) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7845) * $signed(input_fmap_251[7:0]) +
	( 15'sd 14304) * $signed(input_fmap_252[7:0]) +
	( 16'sd 23792) * $signed(input_fmap_253[7:0]) +
	( 16'sd 32605) * $signed(input_fmap_254[7:0]) +
	( 13'sd 2995) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_156;
assign conv_mac_156 = 
	( 14'sd 7453) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32749) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25615) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23409) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26845) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21706) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4131) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25290) * $signed(input_fmap_7[7:0]) +
	( 16'sd 29473) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28733) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9762) * $signed(input_fmap_10[7:0]) +
	( 11'sd 736) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20180) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18810) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9316) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1315) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11673) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28240) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12804) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20240) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6254) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12272) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_25[7:0]) +
	( 11'sd 807) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7804) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26428) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6329) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17149) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17330) * $signed(input_fmap_31[7:0]) +
	( 15'sd 14054) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32487) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26702) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9689) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24558) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14560) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32364) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20192) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23984) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10704) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14232) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21600) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28750) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10709) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17726) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25364) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10349) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23298) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4638) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30163) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4261) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19280) * $signed(input_fmap_53[7:0]) +
	( 15'sd 12627) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9240) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28168) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23214) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30622) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32133) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32092) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18297) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23349) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19633) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5900) * $signed(input_fmap_64[7:0]) +
	( 10'sd 343) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15672) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18693) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23606) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9057) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5407) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32494) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13641) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26687) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25935) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20842) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31404) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27526) * $signed(input_fmap_77[7:0]) +
	( 16'sd 32306) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6814) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10617) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26603) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19440) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9074) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26666) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18808) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28234) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28017) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6054) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13914) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26540) * $signed(input_fmap_92[7:0]) +
	( 10'sd 395) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23585) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23189) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29124) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17057) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19260) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20939) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28432) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7616) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28393) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22440) * $signed(input_fmap_103[7:0]) +
	( 16'sd 29563) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1277) * $signed(input_fmap_105[7:0]) +
	( 11'sd 689) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_108[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20001) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30110) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27273) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4653) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10880) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14695) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23061) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12280) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8420) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30927) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12247) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4228) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27681) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28841) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24224) * $signed(input_fmap_127[7:0]) +
	( 16'sd 20535) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24471) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1459) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3107) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5037) * $signed(input_fmap_132[7:0]) +
	( 13'sd 3076) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31459) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20496) * $signed(input_fmap_135[7:0]) +
	( 16'sd 18694) * $signed(input_fmap_136[7:0]) +
	( 12'sd 1679) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22038) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28526) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17717) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10892) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14226) * $signed(input_fmap_142[7:0]) +
	( 11'sd 956) * $signed(input_fmap_143[7:0]) +
	( 15'sd 10386) * $signed(input_fmap_144[7:0]) +
	( 16'sd 20603) * $signed(input_fmap_145[7:0]) +
	( 16'sd 26999) * $signed(input_fmap_146[7:0]) +
	( 8'sd 92) * $signed(input_fmap_147[7:0]) +
	( 15'sd 10712) * $signed(input_fmap_148[7:0]) +
	( 16'sd 30572) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21114) * $signed(input_fmap_150[7:0]) +
	( 15'sd 10347) * $signed(input_fmap_151[7:0]) +
	( 15'sd 9152) * $signed(input_fmap_152[7:0]) +
	( 16'sd 20647) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_154[7:0]) +
	( 16'sd 21718) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20308) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5918) * $signed(input_fmap_157[7:0]) +
	( 16'sd 21408) * $signed(input_fmap_158[7:0]) +
	( 14'sd 8185) * $signed(input_fmap_159[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_160[7:0]) +
	( 15'sd 15184) * $signed(input_fmap_161[7:0]) +
	( 14'sd 5531) * $signed(input_fmap_162[7:0]) +
	( 15'sd 13847) * $signed(input_fmap_163[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10455) * $signed(input_fmap_165[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_166[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1028) * $signed(input_fmap_168[7:0]) +
	( 16'sd 28261) * $signed(input_fmap_169[7:0]) +
	( 16'sd 21611) * $signed(input_fmap_170[7:0]) +
	( 16'sd 22536) * $signed(input_fmap_171[7:0]) +
	( 9'sd 217) * $signed(input_fmap_172[7:0]) +
	( 16'sd 16492) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6609) * $signed(input_fmap_174[7:0]) +
	( 15'sd 14835) * $signed(input_fmap_175[7:0]) +
	( 16'sd 31423) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_177[7:0]) +
	( 13'sd 3338) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3286) * $signed(input_fmap_179[7:0]) +
	( 16'sd 22672) * $signed(input_fmap_180[7:0]) +
	( 16'sd 20314) * $signed(input_fmap_181[7:0]) +
	( 13'sd 2267) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27915) * $signed(input_fmap_183[7:0]) +
	( 11'sd 945) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26180) * $signed(input_fmap_185[7:0]) +
	( 14'sd 7549) * $signed(input_fmap_186[7:0]) +
	( 16'sd 26999) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23712) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2227) * $signed(input_fmap_189[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_190[7:0]) +
	( 14'sd 6527) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31556) * $signed(input_fmap_192[7:0]) +
	( 10'sd 360) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_194[7:0]) +
	( 16'sd 31035) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25560) * $signed(input_fmap_196[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_197[7:0]) +
	( 16'sd 23458) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23236) * $signed(input_fmap_199[7:0]) +
	( 16'sd 16693) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9651) * $signed(input_fmap_201[7:0]) +
	( 16'sd 24589) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13446) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19703) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11054) * $signed(input_fmap_205[7:0]) +
	( 14'sd 7176) * $signed(input_fmap_206[7:0]) +
	( 15'sd 10696) * $signed(input_fmap_207[7:0]) +
	( 11'sd 785) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3683) * $signed(input_fmap_209[7:0]) +
	( 15'sd 16035) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12918) * $signed(input_fmap_211[7:0]) +
	( 14'sd 7935) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23311) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23900) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23981) * $signed(input_fmap_215[7:0]) +
	( 14'sd 6379) * $signed(input_fmap_216[7:0]) +
	( 14'sd 6155) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19298) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27319) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19801) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24238) * $signed(input_fmap_223[7:0]) +
	( 15'sd 9921) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1705) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29512) * $signed(input_fmap_226[7:0]) +
	( 15'sd 12721) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2388) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23593) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7336) * $signed(input_fmap_230[7:0]) +
	( 12'sd 2019) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12684) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3417) * $signed(input_fmap_233[7:0]) +
	( 16'sd 27083) * $signed(input_fmap_234[7:0]) +
	( 16'sd 31739) * $signed(input_fmap_235[7:0]) +
	( 16'sd 18508) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20361) * $signed(input_fmap_237[7:0]) +
	( 16'sd 29086) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_239[7:0]) +
	( 16'sd 16736) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27491) * $signed(input_fmap_242[7:0]) +
	( 16'sd 17817) * $signed(input_fmap_243[7:0]) +
	( 16'sd 29928) * $signed(input_fmap_244[7:0]) +
	( 16'sd 27184) * $signed(input_fmap_245[7:0]) +
	( 14'sd 7927) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30879) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21534) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17162) * $signed(input_fmap_249[7:0]) +
	( 15'sd 13207) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27375) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30532) * $signed(input_fmap_252[7:0]) +
	( 15'sd 16295) * $signed(input_fmap_253[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_157;
assign conv_mac_157 = 
	( 12'sd 1479) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15810) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11147) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26449) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21337) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12527) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14636) * $signed(input_fmap_6[7:0]) +
	( 15'sd 11119) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3723) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28641) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7242) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31199) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12380) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10900) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3293) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5595) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31404) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26057) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30551) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4556) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31882) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25189) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5952) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21826) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23885) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8712) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28741) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13925) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27069) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29555) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22654) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14222) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9759) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28977) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2262) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2819) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8890) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6410) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21106) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27838) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3775) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16081) * $signed(input_fmap_44[7:0]) +
	( 16'sd 31707) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3273) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12823) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17408) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16648) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29015) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4871) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25812) * $signed(input_fmap_52[7:0]) +
	( 15'sd 9992) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24005) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4706) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14464) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29695) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30928) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14475) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22029) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30030) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4339) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1256) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13737) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20234) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7974) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17300) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13946) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28168) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27481) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25178) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14630) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14231) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14801) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15303) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25280) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21803) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7189) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10478) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6350) * $signed(input_fmap_80[7:0]) +
	( 16'sd 21271) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22739) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18399) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18972) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29060) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_86[7:0]) +
	( 15'sd 9118) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14374) * $signed(input_fmap_88[7:0]) +
	( 11'sd 624) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22910) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3196) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4398) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30178) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1524) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32637) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25827) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4782) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2446) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21265) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5393) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9840) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7893) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27433) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21662) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18324) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11658) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32000) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22673) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23868) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4506) * $signed(input_fmap_114[7:0]) +
	( 16'sd 28681) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29763) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25294) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16638) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29855) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8637) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3084) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32370) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24431) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26107) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5175) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4371) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5989) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12573) * $signed(input_fmap_130[7:0]) +
	( 16'sd 22197) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14234) * $signed(input_fmap_132[7:0]) +
	( 15'sd 16239) * $signed(input_fmap_133[7:0]) +
	( 11'sd 829) * $signed(input_fmap_134[7:0]) +
	( 16'sd 30795) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12468) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9287) * $signed(input_fmap_137[7:0]) +
	( 16'sd 28661) * $signed(input_fmap_138[7:0]) +
	( 15'sd 9941) * $signed(input_fmap_139[7:0]) +
	( 15'sd 12596) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29286) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14667) * $signed(input_fmap_142[7:0]) +
	( 16'sd 18677) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3195) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7256) * $signed(input_fmap_145[7:0]) +
	( 15'sd 16022) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_147[7:0]) +
	( 16'sd 30267) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15535) * $signed(input_fmap_149[7:0]) +
	( 14'sd 4722) * $signed(input_fmap_150[7:0]) +
	( 15'sd 9072) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22534) * $signed(input_fmap_152[7:0]) +
	( 16'sd 32112) * $signed(input_fmap_153[7:0]) +
	( 12'sd 1481) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13334) * $signed(input_fmap_155[7:0]) +
	( 16'sd 27457) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29836) * $signed(input_fmap_157[7:0]) +
	( 16'sd 31456) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27951) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17632) * $signed(input_fmap_160[7:0]) +
	( 16'sd 21443) * $signed(input_fmap_161[7:0]) +
	( 14'sd 7384) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19349) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12441) * $signed(input_fmap_165[7:0]) +
	( 15'sd 15431) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_167[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27000) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23058) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18137) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15289) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19723) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19259) * $signed(input_fmap_174[7:0]) +
	( 10'sd 412) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20412) * $signed(input_fmap_176[7:0]) +
	( 16'sd 25171) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1331) * $signed(input_fmap_178[7:0]) +
	( 16'sd 16621) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27000) * $signed(input_fmap_180[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5193) * $signed(input_fmap_182[7:0]) +
	( 16'sd 19963) * $signed(input_fmap_183[7:0]) +
	( 16'sd 27670) * $signed(input_fmap_184[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_185[7:0]) +
	( 14'sd 7648) * $signed(input_fmap_186[7:0]) +
	( 16'sd 16446) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17874) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17032) * $signed(input_fmap_189[7:0]) +
	( 14'sd 7519) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_191[7:0]) +
	( 15'sd 11288) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20353) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23857) * $signed(input_fmap_194[7:0]) +
	( 14'sd 6684) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20574) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5984) * $signed(input_fmap_197[7:0]) +
	( 15'sd 8599) * $signed(input_fmap_198[7:0]) +
	( 15'sd 11146) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25703) * $signed(input_fmap_200[7:0]) +
	( 16'sd 19851) * $signed(input_fmap_201[7:0]) +
	( 15'sd 12490) * $signed(input_fmap_202[7:0]) +
	( 13'sd 4042) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14297) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29986) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31176) * $signed(input_fmap_206[7:0]) +
	( 15'sd 11921) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13820) * $signed(input_fmap_209[7:0]) +
	( 15'sd 14146) * $signed(input_fmap_210[7:0]) +
	( 15'sd 11034) * $signed(input_fmap_211[7:0]) +
	( 15'sd 9255) * $signed(input_fmap_212[7:0]) +
	( 16'sd 17075) * $signed(input_fmap_213[7:0]) +
	( 16'sd 29100) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10278) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17133) * $signed(input_fmap_216[7:0]) +
	( 15'sd 13549) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13989) * $signed(input_fmap_218[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_219[7:0]) +
	( 10'sd 332) * $signed(input_fmap_220[7:0]) +
	( 16'sd 26049) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10185) * $signed(input_fmap_222[7:0]) +
	( 16'sd 30909) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12608) * $signed(input_fmap_224[7:0]) +
	( 16'sd 25247) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18254) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14525) * $signed(input_fmap_227[7:0]) +
	( 15'sd 15080) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3772) * $signed(input_fmap_229[7:0]) +
	( 15'sd 12552) * $signed(input_fmap_230[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_231[7:0]) +
	( 15'sd 10152) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1078) * $signed(input_fmap_233[7:0]) +
	( 16'sd 21110) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22274) * $signed(input_fmap_235[7:0]) +
	( 14'sd 6552) * $signed(input_fmap_236[7:0]) +
	( 14'sd 5917) * $signed(input_fmap_237[7:0]) +
	( 16'sd 25569) * $signed(input_fmap_238[7:0]) +
	( 15'sd 8324) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_240[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_241[7:0]) +
	( 16'sd 24901) * $signed(input_fmap_242[7:0]) +
	( 16'sd 24772) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6862) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_245[7:0]) +
	( 16'sd 29189) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8869) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3225) * $signed(input_fmap_248[7:0]) +
	( 16'sd 19334) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22907) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_251[7:0]) +
	( 16'sd 22460) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24001) * $signed(input_fmap_253[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14802) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_158;
assign conv_mac_158 = 
	( 16'sd 18126) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5852) * $signed(input_fmap_1[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14974) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17989) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9255) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6285) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4274) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18389) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12044) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8971) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29813) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15368) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26177) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28188) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15885) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20166) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26993) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25801) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16153) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19052) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29741) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12718) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11932) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20555) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19070) * $signed(input_fmap_28[7:0]) +
	( 15'sd 10509) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25873) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_31[7:0]) +
	( 15'sd 11538) * $signed(input_fmap_32[7:0]) +
	( 12'sd 2019) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27171) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17658) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11016) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24938) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23983) * $signed(input_fmap_39[7:0]) +
	( 16'sd 29267) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11973) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28482) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7103) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16272) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30315) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19370) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8700) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3998) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2833) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6827) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9834) * $signed(input_fmap_51[7:0]) +
	( 11'sd 549) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21051) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26153) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25788) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21547) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10445) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23332) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4681) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28489) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30388) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26353) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13422) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20717) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16045) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24023) * $signed(input_fmap_67[7:0]) +
	( 15'sd 8822) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29527) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29143) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27148) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15060) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10958) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19539) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32094) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12809) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4367) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13147) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10281) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19220) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31559) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1559) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11979) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4744) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25460) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18171) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14962) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21030) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17119) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_92[7:0]) +
	( 8'sd 84) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13998) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25062) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15832) * $signed(input_fmap_96[7:0]) +
	( 14'sd 8081) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5979) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8800) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_100[7:0]) +
	( 14'sd 8038) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13868) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_103[7:0]) +
	( 11'sd 914) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17132) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31340) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31550) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24011) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29084) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12793) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1472) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10670) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23041) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32427) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27935) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11687) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4711) * $signed(input_fmap_117[7:0]) +
	( 11'sd 537) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9171) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5724) * $signed(input_fmap_121[7:0]) +
	( 13'sd 4020) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6836) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14771) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22173) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25655) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3056) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18941) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17472) * $signed(input_fmap_129[7:0]) +
	( 14'sd 5127) * $signed(input_fmap_130[7:0]) +
	( 9'sd 236) * $signed(input_fmap_131[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_132[7:0]) +
	( 13'sd 3605) * $signed(input_fmap_133[7:0]) +
	( 15'sd 15965) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27684) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21815) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26981) * $signed(input_fmap_137[7:0]) +
	( 16'sd 26067) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_139[7:0]) +
	( 16'sd 23549) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13988) * $signed(input_fmap_141[7:0]) +
	( 16'sd 24948) * $signed(input_fmap_142[7:0]) +
	( 9'sd 251) * $signed(input_fmap_143[7:0]) +
	( 15'sd 15505) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22947) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3692) * $signed(input_fmap_146[7:0]) +
	( 16'sd 16718) * $signed(input_fmap_147[7:0]) +
	( 10'sd 402) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7312) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25599) * $signed(input_fmap_150[7:0]) +
	( 9'sd 161) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20464) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24319) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_154[7:0]) +
	( 16'sd 21752) * $signed(input_fmap_155[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_156[7:0]) +
	( 15'sd 12217) * $signed(input_fmap_157[7:0]) +
	( 13'sd 3791) * $signed(input_fmap_158[7:0]) +
	( 16'sd 30372) * $signed(input_fmap_159[7:0]) +
	( 15'sd 15237) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_161[7:0]) +
	( 15'sd 15712) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28313) * $signed(input_fmap_163[7:0]) +
	( 14'sd 7650) * $signed(input_fmap_164[7:0]) +
	( 16'sd 25743) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22991) * $signed(input_fmap_166[7:0]) +
	( 16'sd 21273) * $signed(input_fmap_167[7:0]) +
	( 15'sd 8579) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6949) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31151) * $signed(input_fmap_170[7:0]) +
	( 15'sd 15713) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6946) * $signed(input_fmap_172[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6312) * $signed(input_fmap_174[7:0]) +
	( 15'sd 13426) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15943) * $signed(input_fmap_176[7:0]) +
	( 16'sd 32132) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2603) * $signed(input_fmap_178[7:0]) +
	( 16'sd 31597) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4697) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25906) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10792) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_183[7:0]) +
	( 16'sd 16448) * $signed(input_fmap_184[7:0]) +
	( 15'sd 8737) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3120) * $signed(input_fmap_186[7:0]) +
	( 15'sd 13072) * $signed(input_fmap_187[7:0]) +
	( 16'sd 18241) * $signed(input_fmap_188[7:0]) +
	( 16'sd 18108) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31569) * $signed(input_fmap_190[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_191[7:0]) +
	( 16'sd 23170) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11032) * $signed(input_fmap_193[7:0]) +
	( 16'sd 32189) * $signed(input_fmap_194[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_195[7:0]) +
	( 12'sd 1543) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26396) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_198[7:0]) +
	( 13'sd 2134) * $signed(input_fmap_199[7:0]) +
	( 16'sd 17789) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1465) * $signed(input_fmap_201[7:0]) +
	( 16'sd 30507) * $signed(input_fmap_202[7:0]) +
	( 16'sd 27783) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6746) * $signed(input_fmap_204[7:0]) +
	( 14'sd 4514) * $signed(input_fmap_205[7:0]) +
	( 16'sd 30723) * $signed(input_fmap_206[7:0]) +
	( 14'sd 4359) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18012) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24150) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1992) * $signed(input_fmap_210[7:0]) +
	( 16'sd 21540) * $signed(input_fmap_211[7:0]) +
	( 16'sd 21117) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5430) * $signed(input_fmap_213[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_214[7:0]) +
	( 14'sd 4336) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17812) * $signed(input_fmap_216[7:0]) +
	( 16'sd 31979) * $signed(input_fmap_217[7:0]) +
	( 16'sd 19450) * $signed(input_fmap_218[7:0]) +
	( 16'sd 22966) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13286) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1928) * $signed(input_fmap_221[7:0]) +
	( 11'sd 702) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17654) * $signed(input_fmap_223[7:0]) +
	( 16'sd 28461) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26828) * $signed(input_fmap_225[7:0]) +
	( 16'sd 17614) * $signed(input_fmap_226[7:0]) +
	( 11'sd 512) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31287) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17204) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6610) * $signed(input_fmap_230[7:0]) +
	( 16'sd 30046) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14448) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1661) * $signed(input_fmap_233[7:0]) +
	( 16'sd 29214) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26919) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12726) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6007) * $signed(input_fmap_237[7:0]) +
	( 10'sd 384) * $signed(input_fmap_238[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_239[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_240[7:0]) +
	( 16'sd 31391) * $signed(input_fmap_241[7:0]) +
	( 13'sd 3894) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13468) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19068) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14899) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30792) * $signed(input_fmap_246[7:0]) +
	( 14'sd 7379) * $signed(input_fmap_247[7:0]) +
	( 16'sd 29104) * $signed(input_fmap_248[7:0]) +
	( 16'sd 20677) * $signed(input_fmap_249[7:0]) +
	( 16'sd 23171) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6632) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_252[7:0]) +
	( 16'sd 21090) * $signed(input_fmap_253[7:0]) +
	( 16'sd 18478) * $signed(input_fmap_254[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_159;
assign conv_mac_159 = 
	( 10'sd 496) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5923) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3259) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25856) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22091) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27882) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27183) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27700) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19760) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4130) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30381) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8543) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18183) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31092) * $signed(input_fmap_13[7:0]) +
	( 11'sd 589) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20366) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8651) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13990) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9344) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20866) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20299) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13632) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24802) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4097) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13407) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6858) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13902) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18764) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21240) * $signed(input_fmap_30[7:0]) +
	( 15'sd 8881) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17489) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2110) * $signed(input_fmap_33[7:0]) +
	( 15'sd 15950) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24981) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20087) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5462) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11968) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15112) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22480) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32305) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6347) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28719) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27721) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4647) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16670) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21090) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6801) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22803) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7625) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23052) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23161) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3767) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15786) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3213) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30533) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18938) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4555) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31662) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22908) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18025) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7465) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18666) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32516) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24942) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5243) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10560) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19610) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12936) * $signed(input_fmap_71[7:0]) +
	( 16'sd 29036) * $signed(input_fmap_72[7:0]) +
	( 16'sd 23123) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10493) * $signed(input_fmap_74[7:0]) +
	( 14'sd 8147) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13117) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7876) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14514) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8298) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23532) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16053) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3032) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12097) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32475) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5475) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25462) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32247) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19610) * $signed(input_fmap_89[7:0]) +
	( 13'sd 2712) * $signed(input_fmap_90[7:0]) +
	( 11'sd 872) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3054) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8535) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28208) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21106) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10098) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10881) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17336) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17345) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20815) * $signed(input_fmap_101[7:0]) +
	( 15'sd 15024) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13786) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25604) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24982) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22587) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31889) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18814) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15073) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17316) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2496) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11140) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27088) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1084) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15420) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4771) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22907) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12766) * $signed(input_fmap_118[7:0]) +
	( 15'sd 10861) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15562) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4643) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19507) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2422) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21746) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30446) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13701) * $signed(input_fmap_126[7:0]) +
	( 6'sd 26) * $signed(input_fmap_127[7:0]) +
	( 16'sd 19159) * $signed(input_fmap_128[7:0]) +
	( 16'sd 24703) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27755) * $signed(input_fmap_130[7:0]) +
	( 15'sd 11129) * $signed(input_fmap_131[7:0]) +
	( 15'sd 13008) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28411) * $signed(input_fmap_133[7:0]) +
	( 16'sd 28939) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21742) * $signed(input_fmap_135[7:0]) +
	( 16'sd 18815) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25515) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7442) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28717) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_140[7:0]) +
	( 15'sd 9081) * $signed(input_fmap_141[7:0]) +
	( 13'sd 2267) * $signed(input_fmap_142[7:0]) +
	( 16'sd 27921) * $signed(input_fmap_143[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_144[7:0]) +
	( 15'sd 15717) * $signed(input_fmap_145[7:0]) +
	( 16'sd 20701) * $signed(input_fmap_146[7:0]) +
	( 14'sd 7217) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28037) * $signed(input_fmap_148[7:0]) +
	( 12'sd 1783) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25457) * $signed(input_fmap_150[7:0]) +
	( 15'sd 15242) * $signed(input_fmap_151[7:0]) +
	( 16'sd 28787) * $signed(input_fmap_152[7:0]) +
	( 15'sd 15421) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24438) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10607) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14397) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20663) * $signed(input_fmap_157[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_158[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_159[7:0]) +
	( 15'sd 13598) * $signed(input_fmap_160[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_161[7:0]) +
	( 15'sd 15667) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22347) * $signed(input_fmap_163[7:0]) +
	( 16'sd 26385) * $signed(input_fmap_164[7:0]) +
	( 16'sd 26164) * $signed(input_fmap_165[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23850) * $signed(input_fmap_167[7:0]) +
	( 16'sd 24868) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3327) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5334) * $signed(input_fmap_170[7:0]) +
	( 16'sd 17070) * $signed(input_fmap_171[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_172[7:0]) +
	( 16'sd 31613) * $signed(input_fmap_173[7:0]) +
	( 13'sd 3710) * $signed(input_fmap_174[7:0]) +
	( 16'sd 26797) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15770) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5907) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9141) * $signed(input_fmap_178[7:0]) +
	( 16'sd 23909) * $signed(input_fmap_179[7:0]) +
	( 16'sd 18335) * $signed(input_fmap_180[7:0]) +
	( 16'sd 26782) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_182[7:0]) +
	( 14'sd 6109) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30144) * $signed(input_fmap_184[7:0]) +
	( 15'sd 14598) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23104) * $signed(input_fmap_186[7:0]) +
	( 13'sd 3340) * $signed(input_fmap_187[7:0]) +
	( 16'sd 16706) * $signed(input_fmap_188[7:0]) +
	( 12'sd 1180) * $signed(input_fmap_189[7:0]) +
	( 16'sd 19474) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23224) * $signed(input_fmap_191[7:0]) +
	( 15'sd 13643) * $signed(input_fmap_192[7:0]) +
	( 16'sd 23337) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23987) * $signed(input_fmap_194[7:0]) +
	( 16'sd 16731) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12581) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11500) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10435) * $signed(input_fmap_198[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_199[7:0]) +
	( 15'sd 9172) * $signed(input_fmap_200[7:0]) +
	( 16'sd 19745) * $signed(input_fmap_201[7:0]) +
	( 16'sd 20684) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6505) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17486) * $signed(input_fmap_204[7:0]) +
	( 15'sd 14378) * $signed(input_fmap_205[7:0]) +
	( 16'sd 25130) * $signed(input_fmap_206[7:0]) +
	( 16'sd 25518) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12585) * $signed(input_fmap_208[7:0]) +
	( 15'sd 12394) * $signed(input_fmap_209[7:0]) +
	( 16'sd 29437) * $signed(input_fmap_210[7:0]) +
	( 16'sd 18018) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14720) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28105) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30368) * $signed(input_fmap_214[7:0]) +
	( 11'sd 643) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18001) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30952) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30366) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19772) * $signed(input_fmap_219[7:0]) +
	( 16'sd 20658) * $signed(input_fmap_220[7:0]) +
	( 16'sd 17645) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25728) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25802) * $signed(input_fmap_223[7:0]) +
	( 16'sd 29807) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13543) * $signed(input_fmap_225[7:0]) +
	( 16'sd 28177) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_227[7:0]) +
	( 16'sd 20248) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8825) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29949) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31811) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24856) * $signed(input_fmap_233[7:0]) +
	( 14'sd 6178) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21412) * $signed(input_fmap_235[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_236[7:0]) +
	( 14'sd 7263) * $signed(input_fmap_237[7:0]) +
	( 16'sd 25495) * $signed(input_fmap_238[7:0]) +
	( 14'sd 6901) * $signed(input_fmap_239[7:0]) +
	( 16'sd 32229) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_242[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_243[7:0]) +
	( 15'sd 15689) * $signed(input_fmap_244[7:0]) +
	( 16'sd 32625) * $signed(input_fmap_245[7:0]) +
	( 16'sd 27109) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20171) * $signed(input_fmap_247[7:0]) +
	( 14'sd 5251) * $signed(input_fmap_248[7:0]) +
	( 16'sd 23324) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24512) * $signed(input_fmap_250[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_251[7:0]) +
	( 13'sd 3415) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24014) * $signed(input_fmap_253[7:0]) +
	( 13'sd 3598) * $signed(input_fmap_254[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_160;
assign conv_mac_160 = 
	( 14'sd 7545) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29788) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27161) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19304) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11775) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27775) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27427) * $signed(input_fmap_8[7:0]) +
	( 16'sd 28543) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12291) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12530) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31145) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13690) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18203) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16779) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4884) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8245) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21213) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26426) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8819) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14042) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17925) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2929) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2870) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25089) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9628) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3844) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11455) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1592) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12819) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8960) * $signed(input_fmap_32[7:0]) +
	( 16'sd 30173) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29429) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29354) * $signed(input_fmap_35[7:0]) +
	( 15'sd 11005) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29207) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29237) * $signed(input_fmap_39[7:0]) +
	( 11'sd 901) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10955) * $signed(input_fmap_41[7:0]) +
	( 16'sd 27727) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_43[7:0]) +
	( 10'sd 511) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20380) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31504) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19890) * $signed(input_fmap_47[7:0]) +
	( 11'sd 686) * $signed(input_fmap_48[7:0]) +
	( 16'sd 26152) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15302) * $signed(input_fmap_50[7:0]) +
	( 16'sd 16583) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11474) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15625) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17262) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7197) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19863) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15509) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25590) * $signed(input_fmap_58[7:0]) +
	( 16'sd 30759) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29197) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23948) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3229) * $signed(input_fmap_63[7:0]) +
	( 11'sd 790) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10363) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29215) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29207) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4417) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21731) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7135) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24898) * $signed(input_fmap_71[7:0]) +
	( 15'sd 16323) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5008) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4127) * $signed(input_fmap_74[7:0]) +
	( 11'sd 613) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6937) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3968) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26432) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1564) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21936) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17159) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21234) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23490) * $signed(input_fmap_83[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10863) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1374) * $signed(input_fmap_86[7:0]) +
	( 14'sd 6387) * $signed(input_fmap_87[7:0]) +
	( 15'sd 12098) * $signed(input_fmap_88[7:0]) +
	( 8'sd 101) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27978) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27289) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30293) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25056) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27432) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8494) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5779) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6293) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7175) * $signed(input_fmap_99[7:0]) +
	( 11'sd 675) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23659) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30919) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20567) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21966) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28593) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17912) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21451) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13767) * $signed(input_fmap_110[7:0]) +
	( 15'sd 16157) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28718) * $signed(input_fmap_112[7:0]) +
	( 16'sd 27451) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27244) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27691) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5331) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7919) * $signed(input_fmap_118[7:0]) +
	( 9'sd 188) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25861) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17005) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4841) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26382) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24640) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31924) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18994) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10382) * $signed(input_fmap_127[7:0]) +
	( 12'sd 2045) * $signed(input_fmap_128[7:0]) +
	( 9'sd 167) * $signed(input_fmap_129[7:0]) +
	( 15'sd 15921) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13595) * $signed(input_fmap_131[7:0]) +
	( 16'sd 24719) * $signed(input_fmap_132[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_133[7:0]) +
	( 15'sd 13599) * $signed(input_fmap_134[7:0]) +
	( 14'sd 6165) * $signed(input_fmap_135[7:0]) +
	( 15'sd 16040) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25664) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27397) * $signed(input_fmap_138[7:0]) +
	( 16'sd 23195) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15866) * $signed(input_fmap_140[7:0]) +
	( 14'sd 8071) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19287) * $signed(input_fmap_142[7:0]) +
	( 15'sd 14357) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18452) * $signed(input_fmap_144[7:0]) +
	( 16'sd 32099) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21386) * $signed(input_fmap_146[7:0]) +
	( 14'sd 8034) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3498) * $signed(input_fmap_148[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_149[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_150[7:0]) +
	( 16'sd 27168) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22672) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25963) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22625) * $signed(input_fmap_154[7:0]) +
	( 15'sd 11388) * $signed(input_fmap_155[7:0]) +
	( 16'sd 19548) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20494) * $signed(input_fmap_157[7:0]) +
	( 14'sd 7786) * $signed(input_fmap_158[7:0]) +
	( 16'sd 16998) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22451) * $signed(input_fmap_160[7:0]) +
	( 16'sd 18095) * $signed(input_fmap_161[7:0]) +
	( 16'sd 23244) * $signed(input_fmap_162[7:0]) +
	( 15'sd 12948) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11460) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3382) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17135) * $signed(input_fmap_167[7:0]) +
	( 15'sd 11796) * $signed(input_fmap_168[7:0]) +
	( 16'sd 19807) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7893) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11736) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6035) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18524) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11701) * $signed(input_fmap_174[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_175[7:0]) +
	( 11'sd 514) * $signed(input_fmap_176[7:0]) +
	( 15'sd 8922) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27326) * $signed(input_fmap_178[7:0]) +
	( 15'sd 13231) * $signed(input_fmap_179[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_180[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_181[7:0]) +
	( 16'sd 22937) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2319) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26181) * $signed(input_fmap_184[7:0]) +
	( 16'sd 20079) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2074) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_188[7:0]) +
	( 14'sd 8110) * $signed(input_fmap_189[7:0]) +
	( 15'sd 12914) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15475) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21174) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24118) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24444) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14853) * $signed(input_fmap_197[7:0]) +
	( 12'sd 1734) * $signed(input_fmap_198[7:0]) +
	( 16'sd 30388) * $signed(input_fmap_199[7:0]) +
	( 15'sd 14229) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22374) * $signed(input_fmap_201[7:0]) +
	( 16'sd 25982) * $signed(input_fmap_202[7:0]) +
	( 16'sd 18135) * $signed(input_fmap_203[7:0]) +
	( 8'sd 68) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18974) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20110) * $signed(input_fmap_206[7:0]) +
	( 16'sd 16888) * $signed(input_fmap_207[7:0]) +
	( 16'sd 19813) * $signed(input_fmap_208[7:0]) +
	( 16'sd 31128) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9140) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23491) * $signed(input_fmap_211[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_212[7:0]) +
	( 16'sd 22987) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23604) * $signed(input_fmap_214[7:0]) +
	( 11'sd 904) * $signed(input_fmap_215[7:0]) +
	( 16'sd 21123) * $signed(input_fmap_216[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31460) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3780) * $signed(input_fmap_219[7:0]) +
	( 14'sd 7265) * $signed(input_fmap_220[7:0]) +
	( 16'sd 18037) * $signed(input_fmap_221[7:0]) +
	( 16'sd 22098) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19511) * $signed(input_fmap_223[7:0]) +
	( 13'sd 3652) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26920) * $signed(input_fmap_225[7:0]) +
	( 16'sd 21756) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2518) * $signed(input_fmap_227[7:0]) +
	( 13'sd 4054) * $signed(input_fmap_228[7:0]) +
	( 16'sd 16855) * $signed(input_fmap_229[7:0]) +
	( 10'sd 449) * $signed(input_fmap_230[7:0]) +
	( 11'sd 624) * $signed(input_fmap_231[7:0]) +
	( 16'sd 28830) * $signed(input_fmap_232[7:0]) +
	( 13'sd 2381) * $signed(input_fmap_233[7:0]) +
	( 14'sd 6589) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26022) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28043) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19754) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14232) * $signed(input_fmap_238[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_239[7:0]) +
	( 16'sd 20661) * $signed(input_fmap_240[7:0]) +
	( 16'sd 16444) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1513) * $signed(input_fmap_242[7:0]) +
	( 14'sd 4473) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14135) * $signed(input_fmap_245[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21386) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9361) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12023) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4335) * $signed(input_fmap_251[7:0]) +
	( 15'sd 15401) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_253[7:0]) +
	( 16'sd 24292) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10234) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_161;
assign conv_mac_161 = 
	( 13'sd 3253) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1813) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13957) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8785) * $signed(input_fmap_3[7:0]) +
	( 11'sd 706) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23709) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31413) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12621) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23730) * $signed(input_fmap_8[7:0]) +
	( 14'sd 8099) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17404) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5406) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24787) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26430) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2759) * $signed(input_fmap_15[7:0]) +
	( 15'sd 13463) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2503) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14075) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22033) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17225) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10364) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4750) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25289) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32696) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26770) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8280) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6093) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8840) * $signed(input_fmap_29[7:0]) +
	( 15'sd 14683) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28625) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8850) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4851) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9630) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2943) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27948) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30672) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11116) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19592) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12927) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15237) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7700) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18636) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24084) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3223) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11076) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15544) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32046) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5551) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25613) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22728) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3242) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8107) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12367) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22281) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18565) * $signed(input_fmap_60[7:0]) +
	( 11'sd 969) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24507) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9737) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31389) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20085) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25230) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29366) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2897) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3703) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7601) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23872) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15525) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2830) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23936) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16326) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4319) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28933) * $signed(input_fmap_78[7:0]) +
	( 14'sd 6952) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5984) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16399) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1888) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16374) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26979) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18071) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9488) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14173) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23681) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25061) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17818) * $signed(input_fmap_91[7:0]) +
	( 16'sd 32240) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3841) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22172) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20981) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24732) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26407) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3815) * $signed(input_fmap_98[7:0]) +
	( 14'sd 8153) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10336) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17877) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13570) * $signed(input_fmap_102[7:0]) +
	( 14'sd 5958) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30420) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18099) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7920) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17199) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13732) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22730) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14540) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15200) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31256) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7968) * $signed(input_fmap_113[7:0]) +
	( 7'sd 56) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4944) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5240) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18458) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2108) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28488) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18638) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6961) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10894) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4496) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23207) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19101) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28796) * $signed(input_fmap_127[7:0]) +
	( 12'sd 1827) * $signed(input_fmap_128[7:0]) +
	( 16'sd 32655) * $signed(input_fmap_129[7:0]) +
	( 10'sd 322) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13549) * $signed(input_fmap_131[7:0]) +
	( 16'sd 22820) * $signed(input_fmap_132[7:0]) +
	( 15'sd 9239) * $signed(input_fmap_133[7:0]) +
	( 15'sd 10110) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18242) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4635) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32325) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20075) * $signed(input_fmap_139[7:0]) +
	( 16'sd 19792) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18776) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14363) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26728) * $signed(input_fmap_143[7:0]) +
	( 16'sd 29560) * $signed(input_fmap_144[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1760) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17854) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20673) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18171) * $signed(input_fmap_149[7:0]) +
	( 15'sd 10906) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3031) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2879) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22676) * $signed(input_fmap_154[7:0]) +
	( 16'sd 24323) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25317) * $signed(input_fmap_156[7:0]) +
	( 15'sd 16363) * $signed(input_fmap_157[7:0]) +
	( 15'sd 15543) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_159[7:0]) +
	( 15'sd 12270) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_161[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3984) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1788) * $signed(input_fmap_164[7:0]) +
	( 10'sd 493) * $signed(input_fmap_165[7:0]) +
	( 14'sd 5482) * $signed(input_fmap_166[7:0]) +
	( 16'sd 18901) * $signed(input_fmap_167[7:0]) +
	( 15'sd 15550) * $signed(input_fmap_168[7:0]) +
	( 16'sd 24603) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16480) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31253) * $signed(input_fmap_172[7:0]) +
	( 15'sd 15356) * $signed(input_fmap_173[7:0]) +
	( 16'sd 28574) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7279) * $signed(input_fmap_175[7:0]) +
	( 16'sd 22077) * $signed(input_fmap_176[7:0]) +
	( 10'sd 368) * $signed(input_fmap_177[7:0]) +
	( 15'sd 11975) * $signed(input_fmap_178[7:0]) +
	( 16'sd 21611) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27337) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3762) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5261) * $signed(input_fmap_182[7:0]) +
	( 16'sd 31555) * $signed(input_fmap_183[7:0]) +
	( 16'sd 18950) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_185[7:0]) +
	( 14'sd 5436) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5918) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2666) * $signed(input_fmap_188[7:0]) +
	( 15'sd 8885) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9609) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20083) * $signed(input_fmap_191[7:0]) +
	( 16'sd 26151) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28766) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30871) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27631) * $signed(input_fmap_195[7:0]) +
	( 16'sd 29024) * $signed(input_fmap_196[7:0]) +
	( 16'sd 30466) * $signed(input_fmap_197[7:0]) +
	( 16'sd 23835) * $signed(input_fmap_198[7:0]) +
	( 16'sd 16671) * $signed(input_fmap_199[7:0]) +
	( 13'sd 2495) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13678) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_202[7:0]) +
	( 16'sd 22285) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15333) * $signed(input_fmap_204[7:0]) +
	( 16'sd 23603) * $signed(input_fmap_205[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_206[7:0]) +
	( 11'sd 833) * $signed(input_fmap_207[7:0]) +
	( 15'sd 16342) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7006) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5699) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10431) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26200) * $signed(input_fmap_212[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_213[7:0]) +
	( 15'sd 8875) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17579) * $signed(input_fmap_215[7:0]) +
	( 16'sd 31972) * $signed(input_fmap_216[7:0]) +
	( 14'sd 5130) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26982) * $signed(input_fmap_218[7:0]) +
	( 16'sd 29907) * $signed(input_fmap_219[7:0]) +
	( 16'sd 16614) * $signed(input_fmap_220[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_221[7:0]) +
	( 14'sd 4647) * $signed(input_fmap_222[7:0]) +
	( 14'sd 7864) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6717) * $signed(input_fmap_224[7:0]) +
	( 15'sd 8511) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7055) * $signed(input_fmap_226[7:0]) +
	( 13'sd 4066) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8467) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17717) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6994) * $signed(input_fmap_230[7:0]) +
	( 15'sd 12700) * $signed(input_fmap_231[7:0]) +
	( 10'sd 392) * $signed(input_fmap_232[7:0]) +
	( 14'sd 8054) * $signed(input_fmap_233[7:0]) +
	( 16'sd 30224) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7260) * $signed(input_fmap_235[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6159) * $signed(input_fmap_237[7:0]) +
	( 15'sd 10019) * $signed(input_fmap_238[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_239[7:0]) +
	( 16'sd 21907) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15417) * $signed(input_fmap_241[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_242[7:0]) +
	( 16'sd 27189) * $signed(input_fmap_243[7:0]) +
	( 15'sd 15071) * $signed(input_fmap_244[7:0]) +
	( 9'sd 154) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30613) * $signed(input_fmap_246[7:0]) +
	( 14'sd 6881) * $signed(input_fmap_247[7:0]) +
	( 16'sd 30983) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2184) * $signed(input_fmap_249[7:0]) +
	( 15'sd 8836) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15840) * $signed(input_fmap_251[7:0]) +
	( 13'sd 3198) * $signed(input_fmap_252[7:0]) +
	( 16'sd 16721) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23979) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20719) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_162;
assign conv_mac_162 = 
	( 15'sd 11675) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7676) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7725) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21341) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31091) * $signed(input_fmap_4[7:0]) +
	( 16'sd 29890) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22901) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12437) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26292) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27760) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27307) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21334) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12707) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32092) * $signed(input_fmap_14[7:0]) +
	( 15'sd 12890) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7338) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1260) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28133) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2352) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25332) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24373) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12360) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21517) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8554) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13571) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32508) * $signed(input_fmap_26[7:0]) +
	( 16'sd 24586) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11055) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27968) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15080) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14963) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19517) * $signed(input_fmap_32[7:0]) +
	( 14'sd 6290) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7833) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24259) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8207) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29250) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_38[7:0]) +
	( 15'sd 16327) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12737) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10630) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24961) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1962) * $signed(input_fmap_44[7:0]) +
	( 15'sd 10567) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25238) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29790) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5893) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6699) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1678) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27832) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14537) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28166) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6462) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4705) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24387) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11694) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27262) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6828) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4981) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1833) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28025) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7165) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17780) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14723) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30234) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8481) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9388) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21126) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6016) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21295) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9434) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19323) * $signed(input_fmap_75[7:0]) +
	( 15'sd 14065) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32062) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12808) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24006) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1175) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1793) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31808) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22116) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29127) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31616) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13343) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12609) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9716) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29706) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12862) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13845) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29798) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6742) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10978) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30714) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24359) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1646) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19530) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1415) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26006) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15546) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14836) * $signed(input_fmap_106[7:0]) +
	( 16'sd 17790) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32649) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28520) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7449) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25540) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30916) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18942) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3037) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6486) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28571) * $signed(input_fmap_119[7:0]) +
	( 16'sd 30313) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31024) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14533) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9145) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20383) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9136) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26402) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23629) * $signed(input_fmap_127[7:0]) +
	( 15'sd 11070) * $signed(input_fmap_128[7:0]) +
	( 16'sd 32485) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5553) * $signed(input_fmap_131[7:0]) +
	( 14'sd 7175) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10838) * $signed(input_fmap_133[7:0]) +
	( 15'sd 14538) * $signed(input_fmap_134[7:0]) +
	( 16'sd 25076) * $signed(input_fmap_135[7:0]) +
	( 16'sd 20807) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4681) * $signed(input_fmap_137[7:0]) +
	( 16'sd 23872) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31452) * $signed(input_fmap_139[7:0]) +
	( 14'sd 7851) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12713) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25383) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5273) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19463) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22068) * $signed(input_fmap_145[7:0]) +
	( 16'sd 23448) * $signed(input_fmap_146[7:0]) +
	( 16'sd 29486) * $signed(input_fmap_147[7:0]) +
	( 16'sd 32418) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15490) * $signed(input_fmap_149[7:0]) +
	( 16'sd 32265) * $signed(input_fmap_150[7:0]) +
	( 16'sd 27677) * $signed(input_fmap_151[7:0]) +
	( 13'sd 3004) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31205) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11831) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18365) * $signed(input_fmap_156[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28461) * $signed(input_fmap_158[7:0]) +
	( 16'sd 24743) * $signed(input_fmap_159[7:0]) +
	( 16'sd 19813) * $signed(input_fmap_160[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13260) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30602) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24157) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10416) * $signed(input_fmap_165[7:0]) +
	( 15'sd 11558) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17451) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1271) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27534) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31429) * $signed(input_fmap_170[7:0]) +
	( 16'sd 23104) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_172[7:0]) +
	( 15'sd 10280) * $signed(input_fmap_173[7:0]) +
	( 16'sd 22473) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15767) * $signed(input_fmap_175[7:0]) +
	( 11'sd 544) * $signed(input_fmap_176[7:0]) +
	( 16'sd 25155) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2708) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3729) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15516) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25676) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6498) * $signed(input_fmap_182[7:0]) +
	( 12'sd 1060) * $signed(input_fmap_183[7:0]) +
	( 16'sd 32269) * $signed(input_fmap_184[7:0]) +
	( 13'sd 2087) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4695) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22295) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31088) * $signed(input_fmap_188[7:0]) +
	( 16'sd 29787) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9402) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20958) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19231) * $signed(input_fmap_192[7:0]) +
	( 13'sd 3629) * $signed(input_fmap_193[7:0]) +
	( 16'sd 17584) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5059) * $signed(input_fmap_195[7:0]) +
	( 16'sd 18274) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15441) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27885) * $signed(input_fmap_198[7:0]) +
	( 11'sd 567) * $signed(input_fmap_199[7:0]) +
	( 12'sd 1540) * $signed(input_fmap_200[7:0]) +
	( 16'sd 25042) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7460) * $signed(input_fmap_202[7:0]) +
	( 16'sd 23358) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2738) * $signed(input_fmap_204[7:0]) +
	( 16'sd 17316) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27040) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22918) * $signed(input_fmap_208[7:0]) +
	( 15'sd 15801) * $signed(input_fmap_209[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26374) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26609) * $signed(input_fmap_212[7:0]) +
	( 15'sd 13574) * $signed(input_fmap_213[7:0]) +
	( 16'sd 29968) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7588) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5854) * $signed(input_fmap_216[7:0]) +
	( 15'sd 16017) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10269) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12265) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19175) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12216) * $signed(input_fmap_221[7:0]) +
	( 16'sd 30090) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19138) * $signed(input_fmap_223[7:0]) +
	( 14'sd 5239) * $signed(input_fmap_224[7:0]) +
	( 16'sd 22622) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32048) * $signed(input_fmap_226[7:0]) +
	( 16'sd 21890) * $signed(input_fmap_227[7:0]) +
	( 15'sd 9455) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3496) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15104) * $signed(input_fmap_230[7:0]) +
	( 16'sd 22882) * $signed(input_fmap_231[7:0]) +
	( 15'sd 11301) * $signed(input_fmap_232[7:0]) +
	( 16'sd 30900) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5252) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12803) * $signed(input_fmap_236[7:0]) +
	( 16'sd 16964) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19891) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6360) * $signed(input_fmap_240[7:0]) +
	( 14'sd 4400) * $signed(input_fmap_241[7:0]) +
	( 15'sd 16344) * $signed(input_fmap_242[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_243[7:0]) +
	( 15'sd 8862) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2294) * $signed(input_fmap_245[7:0]) +
	( 16'sd 29626) * $signed(input_fmap_246[7:0]) +
	( 16'sd 22148) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10102) * $signed(input_fmap_248[7:0]) +
	( 10'sd 422) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22801) * $signed(input_fmap_250[7:0]) +
	( 16'sd 20853) * $signed(input_fmap_251[7:0]) +
	( 15'sd 15296) * $signed(input_fmap_252[7:0]) +
	( 15'sd 15017) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20859) * $signed(input_fmap_254[7:0]) +
	( 16'sd 29387) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_163;
assign conv_mac_163 = 
	( 13'sd 2864) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24935) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9898) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14542) * $signed(input_fmap_4[7:0]) +
	( 16'sd 24645) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19700) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12170) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31536) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22064) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28203) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8885) * $signed(input_fmap_12[7:0]) +
	( 16'sd 21259) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24211) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8289) * $signed(input_fmap_15[7:0]) +
	( 16'sd 16825) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26766) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9263) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18307) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6604) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24560) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26631) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17602) * $signed(input_fmap_23[7:0]) +
	( 16'sd 16586) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1724) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26639) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4163) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13183) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1938) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29805) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20314) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19717) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7035) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27336) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12096) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4503) * $signed(input_fmap_37[7:0]) +
	( 14'sd 5763) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14484) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5626) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28968) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14729) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26572) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1656) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30717) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31019) * $signed(input_fmap_47[7:0]) +
	( 16'sd 17915) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17016) * $signed(input_fmap_49[7:0]) +
	( 15'sd 16173) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6091) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32122) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2847) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5856) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11430) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6653) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25828) * $signed(input_fmap_57[7:0]) +
	( 15'sd 16164) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17596) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4685) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23156) * $signed(input_fmap_63[7:0]) +
	( 15'sd 9336) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7290) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1435) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28758) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17775) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11214) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16332) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18130) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12205) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30297) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25874) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1830) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30848) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3996) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13462) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24602) * $signed(input_fmap_81[7:0]) +
	( 14'sd 8067) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20164) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27745) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9354) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31914) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15635) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10902) * $signed(input_fmap_88[7:0]) +
	( 16'sd 22198) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20140) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20929) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12949) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20417) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18338) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19545) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30922) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26563) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5931) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1659) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21699) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10248) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7372) * $signed(input_fmap_103[7:0]) +
	( 6'sd 21) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32070) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21689) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2145) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6270) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12636) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32349) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32752) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24296) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1913) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14546) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16668) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2372) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8933) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29575) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2277) * $signed(input_fmap_119[7:0]) +
	( 14'sd 8085) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30059) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1974) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18854) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30602) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29018) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27085) * $signed(input_fmap_127[7:0]) +
	( 16'sd 21437) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14747) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27219) * $signed(input_fmap_130[7:0]) +
	( 16'sd 16942) * $signed(input_fmap_131[7:0]) +
	( 11'sd 683) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29251) * $signed(input_fmap_133[7:0]) +
	( 16'sd 23371) * $signed(input_fmap_134[7:0]) +
	( 16'sd 29559) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15147) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6311) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11008) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_139[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_140[7:0]) +
	( 16'sd 30369) * $signed(input_fmap_141[7:0]) +
	( 12'sd 1373) * $signed(input_fmap_142[7:0]) +
	( 15'sd 11968) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31088) * $signed(input_fmap_144[7:0]) +
	( 16'sd 18888) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14424) * $signed(input_fmap_146[7:0]) +
	( 15'sd 10162) * $signed(input_fmap_147[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_148[7:0]) +
	( 16'sd 28997) * $signed(input_fmap_149[7:0]) +
	( 15'sd 12809) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17341) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7497) * $signed(input_fmap_152[7:0]) +
	( 16'sd 26911) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4415) * $signed(input_fmap_154[7:0]) +
	( 14'sd 6380) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18503) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18885) * $signed(input_fmap_157[7:0]) +
	( 15'sd 15008) * $signed(input_fmap_158[7:0]) +
	( 16'sd 18968) * $signed(input_fmap_159[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_160[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_162[7:0]) +
	( 15'sd 10669) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19630) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4701) * $signed(input_fmap_165[7:0]) +
	( 16'sd 26910) * $signed(input_fmap_166[7:0]) +
	( 16'sd 32440) * $signed(input_fmap_167[7:0]) +
	( 14'sd 4512) * $signed(input_fmap_168[7:0]) +
	( 13'sd 2597) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17824) * $signed(input_fmap_170[7:0]) +
	( 13'sd 2745) * $signed(input_fmap_171[7:0]) +
	( 16'sd 25005) * $signed(input_fmap_172[7:0]) +
	( 15'sd 13400) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14505) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25666) * $signed(input_fmap_175[7:0]) +
	( 16'sd 23573) * $signed(input_fmap_176[7:0]) +
	( 16'sd 32689) * $signed(input_fmap_177[7:0]) +
	( 16'sd 16621) * $signed(input_fmap_178[7:0]) +
	( 16'sd 31350) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15079) * $signed(input_fmap_180[7:0]) +
	( 15'sd 8818) * $signed(input_fmap_181[7:0]) +
	( 16'sd 23300) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17189) * $signed(input_fmap_183[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_184[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_185[7:0]) +
	( 12'sd 1873) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11870) * $signed(input_fmap_187[7:0]) +
	( 16'sd 18296) * $signed(input_fmap_188[7:0]) +
	( 15'sd 13308) * $signed(input_fmap_189[7:0]) +
	( 16'sd 26961) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29835) * $signed(input_fmap_191[7:0]) +
	( 16'sd 21760) * $signed(input_fmap_192[7:0]) +
	( 13'sd 4026) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23413) * $signed(input_fmap_194[7:0]) +
	( 13'sd 2612) * $signed(input_fmap_195[7:0]) +
	( 16'sd 26598) * $signed(input_fmap_196[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_197[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_198[7:0]) +
	( 16'sd 30689) * $signed(input_fmap_199[7:0]) +
	( 16'sd 24916) * $signed(input_fmap_200[7:0]) +
	( 16'sd 28807) * $signed(input_fmap_201[7:0]) +
	( 15'sd 10096) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2386) * $signed(input_fmap_203[7:0]) +
	( 16'sd 25603) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12286) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3880) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21668) * $signed(input_fmap_207[7:0]) +
	( 15'sd 9160) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_209[7:0]) +
	( 16'sd 29842) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6636) * $signed(input_fmap_211[7:0]) +
	( 16'sd 27982) * $signed(input_fmap_212[7:0]) +
	( 16'sd 26407) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23020) * $signed(input_fmap_214[7:0]) +
	( 16'sd 30799) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20139) * $signed(input_fmap_216[7:0]) +
	( 14'sd 7172) * $signed(input_fmap_217[7:0]) +
	( 16'sd 17358) * $signed(input_fmap_218[7:0]) +
	( 15'sd 11216) * $signed(input_fmap_219[7:0]) +
	( 16'sd 23011) * $signed(input_fmap_220[7:0]) +
	( 14'sd 4600) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15260) * $signed(input_fmap_222[7:0]) +
	( 16'sd 20732) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13382) * $signed(input_fmap_224[7:0]) +
	( 14'sd 6374) * $signed(input_fmap_225[7:0]) +
	( 16'sd 29506) * $signed(input_fmap_226[7:0]) +
	( 16'sd 17079) * $signed(input_fmap_227[7:0]) +
	( 9'sd 196) * $signed(input_fmap_228[7:0]) +
	( 12'sd 1895) * $signed(input_fmap_229[7:0]) +
	( 16'sd 25271) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18350) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9356) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15127) * $signed(input_fmap_233[7:0]) +
	( 16'sd 25490) * $signed(input_fmap_234[7:0]) +
	( 14'sd 6923) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27709) * $signed(input_fmap_236[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_237[7:0]) +
	( 14'sd 7277) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12794) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10907) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26368) * $signed(input_fmap_241[7:0]) +
	( 15'sd 9083) * $signed(input_fmap_242[7:0]) +
	( 16'sd 21651) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19781) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10873) * $signed(input_fmap_245[7:0]) +
	( 14'sd 6606) * $signed(input_fmap_246[7:0]) +
	( 16'sd 19068) * $signed(input_fmap_247[7:0]) +
	( 15'sd 13767) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17155) * $signed(input_fmap_249[7:0]) +
	( 14'sd 4197) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2380) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4843) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28202) * $signed(input_fmap_253[7:0]) +
	( 15'sd 14308) * $signed(input_fmap_254[7:0]) +
	( 16'sd 22476) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_164;
assign conv_mac_164 = 
	( 16'sd 27909) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32476) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31307) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7548) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2605) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12902) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9709) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9487) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7496) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15563) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29204) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2321) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14848) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17851) * $signed(input_fmap_17[7:0]) +
	( 15'sd 13066) * $signed(input_fmap_18[7:0]) +
	( 16'sd 16869) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20855) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8984) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26981) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26145) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3941) * $signed(input_fmap_26[7:0]) +
	( 11'sd 568) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20993) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30084) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4803) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2612) * $signed(input_fmap_31[7:0]) +
	( 16'sd 21865) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14432) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9739) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9031) * $signed(input_fmap_35[7:0]) +
	( 15'sd 13758) * $signed(input_fmap_36[7:0]) +
	( 16'sd 16856) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20416) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28800) * $signed(input_fmap_39[7:0]) +
	( 16'sd 16811) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28932) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_42[7:0]) +
	( 15'sd 11542) * $signed(input_fmap_43[7:0]) +
	( 16'sd 28499) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7313) * $signed(input_fmap_45[7:0]) +
	( 15'sd 12713) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25297) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2822) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5923) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5337) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26903) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22753) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3905) * $signed(input_fmap_54[7:0]) +
	( 14'sd 6875) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4450) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32409) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19774) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4681) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27793) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29204) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11342) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17367) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22053) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11225) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16027) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9795) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4401) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27412) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25710) * $signed(input_fmap_72[7:0]) +
	( 14'sd 5788) * $signed(input_fmap_73[7:0]) +
	( 10'sd 359) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13363) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_77[7:0]) +
	( 15'sd 14573) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10638) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26453) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14126) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14755) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3510) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24862) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25887) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8868) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30088) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13057) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32621) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15853) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2352) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12208) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5638) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31488) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22750) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3810) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14444) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18148) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19499) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16356) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4685) * $signed(input_fmap_102[7:0]) +
	( 13'sd 4093) * $signed(input_fmap_103[7:0]) +
	( 11'sd 890) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1860) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10054) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1750) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7987) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22502) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8981) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2189) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21247) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11677) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16528) * $signed(input_fmap_114[7:0]) +
	( 16'sd 18470) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23313) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14125) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14795) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14052) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7545) * $signed(input_fmap_121[7:0]) +
	( 11'sd 822) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25225) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26504) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12991) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1072) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23667) * $signed(input_fmap_127[7:0]) +
	( 16'sd 28419) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17124) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25748) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3730) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5319) * $signed(input_fmap_132[7:0]) +
	( 16'sd 19487) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18398) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18656) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_136[7:0]) +
	( 16'sd 21839) * $signed(input_fmap_137[7:0]) +
	( 15'sd 15796) * $signed(input_fmap_138[7:0]) +
	( 16'sd 19204) * $signed(input_fmap_139[7:0]) +
	( 15'sd 12429) * $signed(input_fmap_140[7:0]) +
	( 14'sd 6051) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27194) * $signed(input_fmap_142[7:0]) +
	( 13'sd 3918) * $signed(input_fmap_143[7:0]) +
	( 16'sd 27349) * $signed(input_fmap_144[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_145[7:0]) +
	( 15'sd 10872) * $signed(input_fmap_146[7:0]) +
	( 15'sd 15550) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20849) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12874) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15288) * $signed(input_fmap_150[7:0]) +
	( 14'sd 5811) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31809) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10226) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7883) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30607) * $signed(input_fmap_155[7:0]) +
	( 16'sd 30083) * $signed(input_fmap_156[7:0]) +
	( 16'sd 17336) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1214) * $signed(input_fmap_158[7:0]) +
	( 15'sd 9567) * $signed(input_fmap_159[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_160[7:0]) +
	( 13'sd 2718) * $signed(input_fmap_161[7:0]) +
	( 13'sd 3097) * $signed(input_fmap_162[7:0]) +
	( 16'sd 25924) * $signed(input_fmap_163[7:0]) +
	( 16'sd 17339) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2514) * $signed(input_fmap_165[7:0]) +
	( 16'sd 23977) * $signed(input_fmap_166[7:0]) +
	( 13'sd 2511) * $signed(input_fmap_167[7:0]) +
	( 15'sd 15589) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12703) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20634) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11033) * $signed(input_fmap_171[7:0]) +
	( 15'sd 8539) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5563) * $signed(input_fmap_173[7:0]) +
	( 14'sd 5642) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5094) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18032) * $signed(input_fmap_176[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_177[7:0]) +
	( 15'sd 8726) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25358) * $signed(input_fmap_179[7:0]) +
	( 15'sd 13301) * $signed(input_fmap_180[7:0]) +
	( 14'sd 7362) * $signed(input_fmap_181[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_182[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24733) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22389) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2727) * $signed(input_fmap_186[7:0]) +
	( 16'sd 20626) * $signed(input_fmap_187[7:0]) +
	( 16'sd 25007) * $signed(input_fmap_188[7:0]) +
	( 15'sd 9660) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28574) * $signed(input_fmap_190[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_191[7:0]) +
	( 15'sd 11497) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12012) * $signed(input_fmap_193[7:0]) +
	( 16'sd 31116) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14337) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17480) * $signed(input_fmap_196[7:0]) +
	( 14'sd 4957) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2072) * $signed(input_fmap_198[7:0]) +
	( 16'sd 19112) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3757) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9898) * $signed(input_fmap_201[7:0]) +
	( 14'sd 4435) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25393) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4693) * $signed(input_fmap_204[7:0]) +
	( 16'sd 20691) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20534) * $signed(input_fmap_206[7:0]) +
	( 15'sd 11804) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30072) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3211) * $signed(input_fmap_209[7:0]) +
	( 15'sd 16094) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17740) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18055) * $signed(input_fmap_212[7:0]) +
	( 15'sd 14606) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30611) * $signed(input_fmap_214[7:0]) +
	( 11'sd 663) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1510) * $signed(input_fmap_216[7:0]) +
	( 14'sd 8012) * $signed(input_fmap_217[7:0]) +
	( 6'sd 28) * $signed(input_fmap_218[7:0]) +
	( 16'sd 18224) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25908) * $signed(input_fmap_220[7:0]) +
	( 16'sd 21050) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2303) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22937) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30132) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3656) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7384) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5231) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18940) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29715) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_230[7:0]) +
	( 15'sd 9405) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20412) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10847) * $signed(input_fmap_233[7:0]) +
	( 16'sd 29643) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21659) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11670) * $signed(input_fmap_236[7:0]) +
	( 16'sd 16723) * $signed(input_fmap_237[7:0]) +
	( 14'sd 4237) * $signed(input_fmap_238[7:0]) +
	( 16'sd 24155) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_240[7:0]) +
	( 15'sd 14830) * $signed(input_fmap_241[7:0]) +
	( 13'sd 2854) * $signed(input_fmap_242[7:0]) +
	( 13'sd 3146) * $signed(input_fmap_243[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_244[7:0]) +
	( 16'sd 16551) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28535) * $signed(input_fmap_246[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_247[7:0]) +
	( 15'sd 16138) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4138) * $signed(input_fmap_249[7:0]) +
	( 14'sd 6781) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19742) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30336) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11889) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10092) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14490) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_165;
assign conv_mac_165 = 
	( 15'sd 9348) * $signed(input_fmap_0[7:0]) +
	( 13'sd 4086) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15754) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5059) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27419) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6454) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10905) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16959) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27375) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3374) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25663) * $signed(input_fmap_11[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11567) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9138) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21705) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11888) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1452) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25680) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15766) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6845) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9617) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_22[7:0]) +
	( 12'sd 1123) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11037) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16119) * $signed(input_fmap_26[7:0]) +
	( 15'sd 10400) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17655) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19528) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20634) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2719) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9744) * $signed(input_fmap_32[7:0]) +
	( 14'sd 7154) * $signed(input_fmap_33[7:0]) +
	( 13'sd 4074) * $signed(input_fmap_34[7:0]) +
	( 16'sd 27385) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2391) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21653) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2241) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22571) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28564) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7289) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18033) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25887) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27053) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18373) * $signed(input_fmap_45[7:0]) +
	( 9'sd 222) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3421) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9404) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32660) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24587) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22619) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26560) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21552) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26252) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1126) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6814) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_59[7:0]) +
	( 16'sd 23481) * $signed(input_fmap_60[7:0]) +
	( 11'sd 884) * $signed(input_fmap_61[7:0]) +
	( 16'sd 19149) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26820) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18366) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26492) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3718) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28387) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29008) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1337) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4719) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31838) * $signed(input_fmap_72[7:0]) +
	( 16'sd 16442) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18981) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13022) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12479) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3952) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29337) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13208) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22374) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3129) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28825) * $signed(input_fmap_83[7:0]) +
	( 16'sd 22339) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24376) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17911) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12282) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21056) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7097) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29058) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14269) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26659) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30654) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22490) * $signed(input_fmap_94[7:0]) +
	( 9'sd 244) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32471) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28472) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25594) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28980) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7786) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16141) * $signed(input_fmap_102[7:0]) +
	( 16'sd 24004) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20485) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7046) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30219) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3669) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19286) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15276) * $signed(input_fmap_109[7:0]) +
	( 15'sd 10898) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31556) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24997) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18581) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27042) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12258) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19783) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11878) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11153) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12836) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18028) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13780) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24082) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30485) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21583) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20686) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26925) * $signed(input_fmap_126[7:0]) +
	( 10'sd 326) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4767) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27219) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30159) * $signed(input_fmap_130[7:0]) +
	( 16'sd 27478) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10903) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28752) * $signed(input_fmap_133[7:0]) +
	( 15'sd 16209) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23746) * $signed(input_fmap_135[7:0]) +
	( 14'sd 5115) * $signed(input_fmap_136[7:0]) +
	( 16'sd 19803) * $signed(input_fmap_137[7:0]) +
	( 16'sd 18321) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27453) * $signed(input_fmap_139[7:0]) +
	( 16'sd 20314) * $signed(input_fmap_140[7:0]) +
	( 15'sd 9984) * $signed(input_fmap_141[7:0]) +
	( 15'sd 9210) * $signed(input_fmap_142[7:0]) +
	( 16'sd 25497) * $signed(input_fmap_143[7:0]) +
	( 16'sd 24805) * $signed(input_fmap_144[7:0]) +
	( 11'sd 635) * $signed(input_fmap_145[7:0]) +
	( 16'sd 28119) * $signed(input_fmap_146[7:0]) +
	( 16'sd 22569) * $signed(input_fmap_147[7:0]) +
	( 12'sd 1958) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4321) * $signed(input_fmap_149[7:0]) +
	( 15'sd 12642) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28640) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16791) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1159) * $signed(input_fmap_153[7:0]) +
	( 14'sd 5683) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5460) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14811) * $signed(input_fmap_156[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17136) * $signed(input_fmap_158[7:0]) +
	( 15'sd 10236) * $signed(input_fmap_159[7:0]) +
	( 16'sd 30138) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28156) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14603) * $signed(input_fmap_162[7:0]) +
	( 12'sd 1499) * $signed(input_fmap_163[7:0]) +
	( 16'sd 32159) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11868) * $signed(input_fmap_165[7:0]) +
	( 16'sd 26564) * $signed(input_fmap_166[7:0]) +
	( 16'sd 18243) * $signed(input_fmap_167[7:0]) +
	( 15'sd 10394) * $signed(input_fmap_168[7:0]) +
	( 15'sd 14892) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18234) * $signed(input_fmap_171[7:0]) +
	( 16'sd 29612) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_173[7:0]) +
	( 15'sd 15226) * $signed(input_fmap_174[7:0]) +
	( 13'sd 4060) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13793) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18146) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14076) * $signed(input_fmap_178[7:0]) +
	( 15'sd 8439) * $signed(input_fmap_179[7:0]) +
	( 16'sd 25261) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30202) * $signed(input_fmap_181[7:0]) +
	( 15'sd 8325) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17432) * $signed(input_fmap_183[7:0]) +
	( 15'sd 15997) * $signed(input_fmap_184[7:0]) +
	( 15'sd 14546) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_186[7:0]) +
	( 16'sd 31414) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32063) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7075) * $signed(input_fmap_189[7:0]) +
	( 14'sd 6628) * $signed(input_fmap_190[7:0]) +
	( 13'sd 2074) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22919) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29404) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23600) * $signed(input_fmap_194[7:0]) +
	( 16'sd 18869) * $signed(input_fmap_195[7:0]) +
	( 16'sd 23138) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1683) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18571) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_199[7:0]) +
	( 10'sd 416) * $signed(input_fmap_200[7:0]) +
	( 16'sd 26834) * $signed(input_fmap_201[7:0]) +
	( 16'sd 29770) * $signed(input_fmap_202[7:0]) +
	( 16'sd 31054) * $signed(input_fmap_203[7:0]) +
	( 16'sd 22587) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30695) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29876) * $signed(input_fmap_206[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_207[7:0]) +
	( 13'sd 2799) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18442) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11371) * $signed(input_fmap_210[7:0]) +
	( 16'sd 29839) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11574) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6035) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28889) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10973) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20004) * $signed(input_fmap_216[7:0]) +
	( 14'sd 6397) * $signed(input_fmap_217[7:0]) +
	( 6'sd 20) * $signed(input_fmap_218[7:0]) +
	( 16'sd 25837) * $signed(input_fmap_219[7:0]) +
	( 15'sd 8803) * $signed(input_fmap_220[7:0]) +
	( 16'sd 22563) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_222[7:0]) +
	( 15'sd 10194) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7587) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3838) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_226[7:0]) +
	( 14'sd 4900) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1680) * $signed(input_fmap_228[7:0]) +
	( 16'sd 25618) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15391) * $signed(input_fmap_230[7:0]) +
	( 16'sd 26451) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12726) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15683) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5027) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_235[7:0]) +
	( 12'sd 1471) * $signed(input_fmap_236[7:0]) +
	( 14'sd 5382) * $signed(input_fmap_237[7:0]) +
	( 16'sd 29504) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26173) * $signed(input_fmap_239[7:0]) +
	( 14'sd 7528) * $signed(input_fmap_240[7:0]) +
	( 11'sd 588) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17490) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2932) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28162) * $signed(input_fmap_244[7:0]) +
	( 15'sd 8327) * $signed(input_fmap_245[7:0]) +
	( 16'sd 25350) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1900) * $signed(input_fmap_248[7:0]) +
	( 16'sd 22040) * $signed(input_fmap_249[7:0]) +
	( 16'sd 23923) * $signed(input_fmap_250[7:0]) +
	( 10'sd 292) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26030) * $signed(input_fmap_252[7:0]) +
	( 16'sd 26870) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19636) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_166;
assign conv_mac_166 = 
	( 15'sd 15036) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18889) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16949) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23018) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11080) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19887) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6849) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23130) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5024) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26485) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19835) * $signed(input_fmap_12[7:0]) +
	( 16'sd 16764) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22578) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23397) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6417) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10638) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2061) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22939) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17185) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6334) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18184) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21491) * $signed(input_fmap_25[7:0]) +
	( 15'sd 9208) * $signed(input_fmap_26[7:0]) +
	( 13'sd 2903) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22970) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30367) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21578) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11653) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29186) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19847) * $signed(input_fmap_33[7:0]) +
	( 15'sd 9406) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6010) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30636) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16023) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32293) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26331) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3084) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13827) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21421) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3804) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22829) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15780) * $signed(input_fmap_45[7:0]) +
	( 16'sd 17812) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26312) * $signed(input_fmap_47[7:0]) +
	( 10'sd 482) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19533) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15595) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18810) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4273) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15408) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24569) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14277) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21761) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2954) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17936) * $signed(input_fmap_59[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_60[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10281) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23063) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19928) * $signed(input_fmap_64[7:0]) +
	( 11'sd 539) * $signed(input_fmap_65[7:0]) +
	( 15'sd 15384) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17960) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4186) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30516) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23761) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3129) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10025) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29167) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29214) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9952) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29074) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23481) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17692) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10880) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4491) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29972) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13899) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19418) * $signed(input_fmap_85[7:0]) +
	( 14'sd 5018) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13264) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24918) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17223) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20847) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13276) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17581) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5781) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12502) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4478) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2551) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27842) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7575) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3359) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12217) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11987) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24878) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17047) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31237) * $signed(input_fmap_107[7:0]) +
	( 16'sd 29626) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9703) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32288) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19180) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21063) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7607) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9743) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20292) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9766) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32078) * $signed(input_fmap_118[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6648) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2578) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12996) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9985) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20338) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1415) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19252) * $signed(input_fmap_129[7:0]) +
	( 15'sd 8392) * $signed(input_fmap_130[7:0]) +
	( 16'sd 21604) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11763) * $signed(input_fmap_132[7:0]) +
	( 16'sd 26068) * $signed(input_fmap_133[7:0]) +
	( 16'sd 27296) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21741) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25981) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15681) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32298) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14558) * $signed(input_fmap_139[7:0]) +
	( 16'sd 19328) * $signed(input_fmap_140[7:0]) +
	( 16'sd 27723) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30653) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10592) * $signed(input_fmap_143[7:0]) +
	( 15'sd 15955) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8385) * $signed(input_fmap_145[7:0]) +
	( 16'sd 17559) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27211) * $signed(input_fmap_147[7:0]) +
	( 15'sd 14427) * $signed(input_fmap_148[7:0]) +
	( 16'sd 21873) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23753) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28619) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24600) * $signed(input_fmap_152[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_153[7:0]) +
	( 16'sd 19805) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7126) * $signed(input_fmap_155[7:0]) +
	( 15'sd 9551) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13849) * $signed(input_fmap_157[7:0]) +
	( 11'sd 535) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5615) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23206) * $signed(input_fmap_161[7:0]) +
	( 15'sd 9151) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28726) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24020) * $signed(input_fmap_164[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_165[7:0]) +
	( 14'sd 5922) * $signed(input_fmap_166[7:0]) +
	( 14'sd 5660) * $signed(input_fmap_167[7:0]) +
	( 15'sd 10496) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3278) * $signed(input_fmap_169[7:0]) +
	( 16'sd 22365) * $signed(input_fmap_170[7:0]) +
	( 16'sd 23148) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11618) * $signed(input_fmap_172[7:0]) +
	( 13'sd 4017) * $signed(input_fmap_173[7:0]) +
	( 16'sd 29377) * $signed(input_fmap_174[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_176[7:0]) +
	( 14'sd 4235) * $signed(input_fmap_177[7:0]) +
	( 16'sd 20400) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5225) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3090) * $signed(input_fmap_180[7:0]) +
	( 14'sd 7294) * $signed(input_fmap_181[7:0]) +
	( 16'sd 28064) * $signed(input_fmap_182[7:0]) +
	( 15'sd 10909) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8393) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25721) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4770) * $signed(input_fmap_186[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12142) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17999) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29115) * $signed(input_fmap_191[7:0]) +
	( 16'sd 32413) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19610) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_194[7:0]) +
	( 15'sd 9284) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7642) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22954) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29781) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1314) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25357) * $signed(input_fmap_200[7:0]) +
	( 15'sd 10313) * $signed(input_fmap_201[7:0]) +
	( 16'sd 23406) * $signed(input_fmap_202[7:0]) +
	( 11'sd 670) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19499) * $signed(input_fmap_204[7:0]) +
	( 15'sd 10971) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6399) * $signed(input_fmap_206[7:0]) +
	( 14'sd 6491) * $signed(input_fmap_207[7:0]) +
	( 14'sd 5418) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7882) * $signed(input_fmap_209[7:0]) +
	( 13'sd 4038) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10343) * $signed(input_fmap_211[7:0]) +
	( 13'sd 3563) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11154) * $signed(input_fmap_213[7:0]) +
	( 15'sd 13662) * $signed(input_fmap_214[7:0]) +
	( 16'sd 26221) * $signed(input_fmap_215[7:0]) +
	( 16'sd 22082) * $signed(input_fmap_216[7:0]) +
	( 16'sd 16956) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28920) * $signed(input_fmap_218[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_219[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_220[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15686) * $signed(input_fmap_222[7:0]) +
	( 16'sd 32110) * $signed(input_fmap_223[7:0]) +
	( 10'sd 263) * $signed(input_fmap_224[7:0]) +
	( 14'sd 4125) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18521) * $signed(input_fmap_226[7:0]) +
	( 14'sd 4544) * $signed(input_fmap_227[7:0]) +
	( 16'sd 20536) * $signed(input_fmap_228[7:0]) +
	( 16'sd 18042) * $signed(input_fmap_229[7:0]) +
	( 16'sd 26831) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31449) * $signed(input_fmap_231[7:0]) +
	( 16'sd 27131) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_233[7:0]) +
	( 14'sd 8133) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11530) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12006) * $signed(input_fmap_236[7:0]) +
	( 16'sd 20841) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28388) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31297) * $signed(input_fmap_239[7:0]) +
	( 16'sd 17097) * $signed(input_fmap_240[7:0]) +
	( 16'sd 31014) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6162) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12933) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2577) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20296) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3599) * $signed(input_fmap_248[7:0]) +
	( 15'sd 11027) * $signed(input_fmap_249[7:0]) +
	( 11'sd 545) * $signed(input_fmap_250[7:0]) +
	( 15'sd 10383) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5738) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13526) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10814) * $signed(input_fmap_254[7:0]) +
	( 16'sd 32295) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_167;
assign conv_mac_167 = 
	( 16'sd 28520) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10691) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22690) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17071) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6377) * $signed(input_fmap_4[7:0]) +
	( 16'sd 31174) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11043) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23873) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31343) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22618) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5049) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5961) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25338) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27196) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14055) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1889) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13667) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20709) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29843) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25996) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30722) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18460) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20044) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13702) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9569) * $signed(input_fmap_27[7:0]) +
	( 16'sd 32238) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11861) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15608) * $signed(input_fmap_31[7:0]) +
	( 15'sd 12138) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11123) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7035) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2405) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3618) * $signed(input_fmap_36[7:0]) +
	( 16'sd 31894) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21766) * $signed(input_fmap_38[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32568) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28156) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20841) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9953) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18777) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3390) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3461) * $signed(input_fmap_47[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_48[7:0]) +
	( 12'sd 1075) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11821) * $signed(input_fmap_50[7:0]) +
	( 16'sd 18423) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6942) * $signed(input_fmap_52[7:0]) +
	( 16'sd 27495) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29732) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26801) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2395) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19340) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14487) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13828) * $signed(input_fmap_60[7:0]) +
	( 16'sd 20777) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13914) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13180) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8847) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13799) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11845) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13794) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17510) * $signed(input_fmap_68[7:0]) +
	( 15'sd 16120) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28280) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30610) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22431) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14316) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11337) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31496) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22708) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29626) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23997) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9868) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1502) * $signed(input_fmap_81[7:0]) +
	( 16'sd 21093) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11092) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20603) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6753) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9739) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27832) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1135) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24344) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20400) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20750) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13579) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12788) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16093) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22752) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30659) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31103) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9267) * $signed(input_fmap_98[7:0]) +
	( 15'sd 12624) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8542) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15595) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5279) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5260) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15314) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2490) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1912) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22907) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8274) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8537) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19759) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22812) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14847) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14228) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8284) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22125) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1820) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3712) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24205) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6848) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13968) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27476) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2059) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7336) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24082) * $signed(input_fmap_125[7:0]) +
	( 15'sd 9777) * $signed(input_fmap_126[7:0]) +
	( 16'sd 32452) * $signed(input_fmap_127[7:0]) +
	( 16'sd 27003) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28633) * $signed(input_fmap_129[7:0]) +
	( 14'sd 7870) * $signed(input_fmap_130[7:0]) +
	( 16'sd 28616) * $signed(input_fmap_131[7:0]) +
	( 14'sd 8078) * $signed(input_fmap_132[7:0]) +
	( 14'sd 7780) * $signed(input_fmap_133[7:0]) +
	( 16'sd 16903) * $signed(input_fmap_134[7:0]) +
	( 15'sd 11690) * $signed(input_fmap_135[7:0]) +
	( 16'sd 24790) * $signed(input_fmap_136[7:0]) +
	( 16'sd 28381) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22795) * $signed(input_fmap_138[7:0]) +
	( 14'sd 6087) * $signed(input_fmap_139[7:0]) +
	( 14'sd 7642) * $signed(input_fmap_140[7:0]) +
	( 11'sd 515) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30955) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26232) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26032) * $signed(input_fmap_145[7:0]) +
	( 16'sd 32139) * $signed(input_fmap_146[7:0]) +
	( 14'sd 8121) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28067) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2057) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5222) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30622) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21832) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4746) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27089) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17031) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30643) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28451) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27179) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21561) * $signed(input_fmap_160[7:0]) +
	( 13'sd 3903) * $signed(input_fmap_161[7:0]) +
	( 15'sd 8641) * $signed(input_fmap_162[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3917) * $signed(input_fmap_164[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_165[7:0]) +
	( 16'sd 20435) * $signed(input_fmap_166[7:0]) +
	( 16'sd 21031) * $signed(input_fmap_167[7:0]) +
	( 16'sd 32697) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27840) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17910) * $signed(input_fmap_170[7:0]) +
	( 16'sd 32341) * $signed(input_fmap_171[7:0]) +
	( 16'sd 25233) * $signed(input_fmap_172[7:0]) +
	( 16'sd 24870) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27580) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28642) * $signed(input_fmap_175[7:0]) +
	( 11'sd 692) * $signed(input_fmap_176[7:0]) +
	( 16'sd 28767) * $signed(input_fmap_177[7:0]) +
	( 15'sd 12587) * $signed(input_fmap_178[7:0]) +
	( 15'sd 10595) * $signed(input_fmap_179[7:0]) +
	( 16'sd 30604) * $signed(input_fmap_180[7:0]) +
	( 16'sd 32607) * $signed(input_fmap_181[7:0]) +
	( 16'sd 24713) * $signed(input_fmap_182[7:0]) +
	( 16'sd 26071) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31265) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11699) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3591) * $signed(input_fmap_186[7:0]) +
	( 16'sd 32257) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21155) * $signed(input_fmap_188[7:0]) +
	( 16'sd 24986) * $signed(input_fmap_189[7:0]) +
	( 16'sd 25338) * $signed(input_fmap_190[7:0]) +
	( 16'sd 16482) * $signed(input_fmap_191[7:0]) +
	( 15'sd 11284) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29179) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12571) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17826) * $signed(input_fmap_195[7:0]) +
	( 16'sd 29635) * $signed(input_fmap_196[7:0]) +
	( 14'sd 6973) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10075) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29264) * $signed(input_fmap_199[7:0]) +
	( 14'sd 4562) * $signed(input_fmap_200[7:0]) +
	( 16'sd 17657) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19960) * $signed(input_fmap_202[7:0]) +
	( 14'sd 7962) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12983) * $signed(input_fmap_204[7:0]) +
	( 15'sd 8232) * $signed(input_fmap_205[7:0]) +
	( 14'sd 5044) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12716) * $signed(input_fmap_207[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_208[7:0]) +
	( 14'sd 5915) * $signed(input_fmap_209[7:0]) +
	( 16'sd 17828) * $signed(input_fmap_210[7:0]) +
	( 16'sd 16545) * $signed(input_fmap_211[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_212[7:0]) +
	( 15'sd 10506) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28461) * $signed(input_fmap_214[7:0]) +
	( 15'sd 12554) * $signed(input_fmap_215[7:0]) +
	( 15'sd 8823) * $signed(input_fmap_216[7:0]) +
	( 15'sd 8842) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31617) * $signed(input_fmap_218[7:0]) +
	( 15'sd 16036) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12855) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28946) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17504) * $signed(input_fmap_223[7:0]) +
	( 16'sd 23979) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7534) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22023) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2824) * $signed(input_fmap_228[7:0]) +
	( 14'sd 7348) * $signed(input_fmap_229[7:0]) +
	( 14'sd 4730) * $signed(input_fmap_230[7:0]) +
	( 16'sd 28690) * $signed(input_fmap_231[7:0]) +
	( 16'sd 17244) * $signed(input_fmap_232[7:0]) +
	( 16'sd 17978) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18023) * $signed(input_fmap_234[7:0]) +
	( 16'sd 25590) * $signed(input_fmap_235[7:0]) +
	( 12'sd 1940) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14383) * $signed(input_fmap_237[7:0]) +
	( 15'sd 10295) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13030) * $signed(input_fmap_239[7:0]) +
	( 10'sd 295) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29633) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27731) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25703) * $signed(input_fmap_243[7:0]) +
	( 15'sd 10277) * $signed(input_fmap_244[7:0]) +
	( 16'sd 27277) * $signed(input_fmap_245[7:0]) +
	( 16'sd 21597) * $signed(input_fmap_246[7:0]) +
	( 16'sd 31461) * $signed(input_fmap_247[7:0]) +
	( 15'sd 11504) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17095) * $signed(input_fmap_249[7:0]) +
	( 14'sd 6888) * $signed(input_fmap_250[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6697) * $signed(input_fmap_252[7:0]) +
	( 12'sd 1714) * $signed(input_fmap_253[7:0]) +
	( 15'sd 8753) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11375) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_168;
assign conv_mac_168 = 
	( 16'sd 18939) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1166) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14057) * $signed(input_fmap_2[7:0]) +
	( 11'sd 702) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25468) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27089) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26230) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7136) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27059) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31378) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5464) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20088) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19852) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16744) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23982) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20735) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29529) * $signed(input_fmap_20[7:0]) +
	( 16'sd 22916) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1549) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6967) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21290) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28592) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22719) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2060) * $signed(input_fmap_28[7:0]) +
	( 14'sd 8053) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26449) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19378) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18128) * $signed(input_fmap_32[7:0]) +
	( 16'sd 23032) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21851) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12293) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17111) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24972) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12683) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17962) * $signed(input_fmap_41[7:0]) +
	( 15'sd 13062) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15192) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27892) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28818) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27581) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25241) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1736) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10266) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28004) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30852) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30039) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5026) * $signed(input_fmap_53[7:0]) +
	( 11'sd 550) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7203) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17440) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5344) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17008) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24635) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7931) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3793) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24304) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28231) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15680) * $signed(input_fmap_64[7:0]) +
	( 16'sd 25773) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8926) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8549) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17940) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9364) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20071) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32461) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20697) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12583) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11540) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16931) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11926) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13945) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3931) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8843) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26245) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27032) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18397) * $signed(input_fmap_83[7:0]) +
	( 11'sd 610) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4214) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25899) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31628) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7953) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26970) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25437) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6089) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10253) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32006) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28087) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25190) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23947) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28872) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23909) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28971) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23624) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13881) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21381) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26082) * $signed(input_fmap_106[7:0]) +
	( 11'sd 582) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12303) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23327) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30192) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22573) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31133) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29615) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14663) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20910) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30864) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15386) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10993) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27696) * $signed(input_fmap_119[7:0]) +
	( 11'sd 937) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23112) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7671) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28119) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9514) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22464) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20037) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1971) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17631) * $signed(input_fmap_128[7:0]) +
	( 16'sd 27105) * $signed(input_fmap_129[7:0]) +
	( 14'sd 5773) * $signed(input_fmap_130[7:0]) +
	( 15'sd 9415) * $signed(input_fmap_131[7:0]) +
	( 16'sd 27787) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29729) * $signed(input_fmap_133[7:0]) +
	( 14'sd 4874) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28521) * $signed(input_fmap_135[7:0]) +
	( 16'sd 29441) * $signed(input_fmap_136[7:0]) +
	( 12'sd 1717) * $signed(input_fmap_137[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24233) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28308) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3114) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21012) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1370) * $signed(input_fmap_143[7:0]) +
	( 11'sd 724) * $signed(input_fmap_144[7:0]) +
	( 14'sd 5328) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27796) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19754) * $signed(input_fmap_147[7:0]) +
	( 15'sd 15796) * $signed(input_fmap_148[7:0]) +
	( 16'sd 29774) * $signed(input_fmap_149[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_150[7:0]) +
	( 16'sd 29085) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14098) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4102) * $signed(input_fmap_153[7:0]) +
	( 16'sd 18931) * $signed(input_fmap_154[7:0]) +
	( 15'sd 11641) * $signed(input_fmap_155[7:0]) +
	( 14'sd 5011) * $signed(input_fmap_156[7:0]) +
	( 15'sd 12867) * $signed(input_fmap_157[7:0]) +
	( 15'sd 16067) * $signed(input_fmap_158[7:0]) +
	( 16'sd 17521) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5283) * $signed(input_fmap_160[7:0]) +
	( 11'sd 517) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14882) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11776) * $signed(input_fmap_164[7:0]) +
	( 14'sd 5569) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3769) * $signed(input_fmap_166[7:0]) +
	( 12'sd 1735) * $signed(input_fmap_167[7:0]) +
	( 16'sd 32078) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17368) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18255) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20596) * $signed(input_fmap_171[7:0]) +
	( 16'sd 21338) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12734) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6790) * $signed(input_fmap_174[7:0]) +
	( 15'sd 9678) * $signed(input_fmap_175[7:0]) +
	( 16'sd 28513) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17526) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2270) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15991) * $signed(input_fmap_180[7:0]) +
	( 16'sd 32297) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10484) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2151) * $signed(input_fmap_183[7:0]) +
	( 16'sd 21589) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17125) * $signed(input_fmap_185[7:0]) +
	( 15'sd 8426) * $signed(input_fmap_186[7:0]) +
	( 15'sd 8351) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32573) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26558) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9386) * $signed(input_fmap_190[7:0]) +
	( 15'sd 13873) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_192[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_193[7:0]) +
	( 15'sd 15154) * $signed(input_fmap_194[7:0]) +
	( 16'sd 23025) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14572) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24535) * $signed(input_fmap_197[7:0]) +
	( 16'sd 30337) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23254) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15961) * $signed(input_fmap_200[7:0]) +
	( 16'sd 30396) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21268) * $signed(input_fmap_202[7:0]) +
	( 16'sd 29281) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17832) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_205[7:0]) +
	( 16'sd 30403) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21922) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3665) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11700) * $signed(input_fmap_210[7:0]) +
	( 14'sd 7179) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12829) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2341) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23167) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7129) * $signed(input_fmap_215[7:0]) +
	( 15'sd 14832) * $signed(input_fmap_216[7:0]) +
	( 14'sd 5470) * $signed(input_fmap_217[7:0]) +
	( 16'sd 23927) * $signed(input_fmap_218[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13078) * $signed(input_fmap_220[7:0]) +
	( 16'sd 32575) * $signed(input_fmap_221[7:0]) +
	( 15'sd 13356) * $signed(input_fmap_222[7:0]) +
	( 16'sd 23169) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13713) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20496) * $signed(input_fmap_225[7:0]) +
	( 16'sd 20864) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27005) * $signed(input_fmap_227[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17624) * $signed(input_fmap_229[7:0]) +
	( 15'sd 10436) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31866) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14682) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14035) * $signed(input_fmap_233[7:0]) +
	( 11'sd 744) * $signed(input_fmap_234[7:0]) +
	( 15'sd 16123) * $signed(input_fmap_235[7:0]) +
	( 16'sd 21350) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10033) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13185) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20659) * $signed(input_fmap_239[7:0]) +
	( 15'sd 11381) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18541) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6456) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18101) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14325) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20374) * $signed(input_fmap_246[7:0]) +
	( 12'sd 2044) * $signed(input_fmap_247[7:0]) +
	( 15'sd 16162) * $signed(input_fmap_248[7:0]) +
	( 16'sd 20465) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30067) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4149) * $signed(input_fmap_251[7:0]) +
	( 13'sd 2245) * $signed(input_fmap_252[7:0]) +
	( 16'sd 22436) * $signed(input_fmap_253[7:0]) +
	( 15'sd 14423) * $signed(input_fmap_254[7:0]) +
	( 15'sd 8474) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_169;
assign conv_mac_169 = 
	( 16'sd 20498) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8203) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15268) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9654) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18389) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5250) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26140) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3571) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22615) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21943) * $signed(input_fmap_12[7:0]) +
	( 14'sd 4919) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9793) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31161) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6601) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22321) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5488) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14731) * $signed(input_fmap_19[7:0]) +
	( 11'sd 518) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23845) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28132) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7655) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3198) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24236) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31513) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1200) * $signed(input_fmap_28[7:0]) +
	( 7'sd 46) * $signed(input_fmap_29[7:0]) +
	( 15'sd 13480) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14715) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2822) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13604) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21995) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29796) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27428) * $signed(input_fmap_36[7:0]) +
	( 16'sd 23531) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27527) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30210) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9342) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32530) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6596) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2491) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12781) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9134) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26296) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15830) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7480) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15206) * $signed(input_fmap_51[7:0]) +
	( 9'sd 181) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14687) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23303) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31640) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16573) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3437) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8700) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3013) * $signed(input_fmap_61[7:0]) +
	( 16'sd 30896) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21259) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24146) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26352) * $signed(input_fmap_66[7:0]) +
	( 16'sd 29808) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19449) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6855) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20155) * $signed(input_fmap_70[7:0]) +
	( 10'sd 256) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2591) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31118) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28855) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13304) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21926) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29295) * $signed(input_fmap_77[7:0]) +
	( 8'sd 70) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2702) * $signed(input_fmap_80[7:0]) +
	( 14'sd 5552) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18716) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15776) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4388) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25740) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26336) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25988) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4216) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20836) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7802) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13324) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30318) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3570) * $signed(input_fmap_95[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6259) * $signed(input_fmap_97[7:0]) +
	( 14'sd 8131) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15195) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16116) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20732) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27157) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8254) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14568) * $signed(input_fmap_105[7:0]) +
	( 11'sd 908) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15994) * $signed(input_fmap_108[7:0]) +
	( 15'sd 15842) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7552) * $signed(input_fmap_110[7:0]) +
	( 16'sd 27400) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18472) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8650) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25509) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24521) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18784) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27215) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28274) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25888) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29629) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23456) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26559) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28956) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29889) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14817) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19385) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9780) * $signed(input_fmap_128[7:0]) +
	( 14'sd 8064) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19329) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31466) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_132[7:0]) +
	( 16'sd 25063) * $signed(input_fmap_133[7:0]) +
	( 16'sd 26930) * $signed(input_fmap_134[7:0]) +
	( 16'sd 17817) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1567) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25319) * $signed(input_fmap_137[7:0]) +
	( 10'sd 311) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8720) * $signed(input_fmap_139[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29612) * $signed(input_fmap_141[7:0]) +
	( 16'sd 29025) * $signed(input_fmap_142[7:0]) +
	( 16'sd 18524) * $signed(input_fmap_143[7:0]) +
	( 15'sd 8837) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22663) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29435) * $signed(input_fmap_146[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_147[7:0]) +
	( 16'sd 31771) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4199) * $signed(input_fmap_149[7:0]) +
	( 16'sd 24418) * $signed(input_fmap_150[7:0]) +
	( 15'sd 10306) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_153[7:0]) +
	( 16'sd 17167) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28324) * $signed(input_fmap_155[7:0]) +
	( 16'sd 22811) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14120) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28263) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4442) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21576) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20121) * $signed(input_fmap_161[7:0]) +
	( 16'sd 25187) * $signed(input_fmap_162[7:0]) +
	( 12'sd 1706) * $signed(input_fmap_163[7:0]) +
	( 14'sd 4888) * $signed(input_fmap_164[7:0]) +
	( 14'sd 7906) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_166[7:0]) +
	( 14'sd 5650) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_169[7:0]) +
	( 15'sd 8618) * $signed(input_fmap_170[7:0]) +
	( 14'sd 5727) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31371) * $signed(input_fmap_172[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27416) * $signed(input_fmap_174[7:0]) +
	( 10'sd 438) * $signed(input_fmap_175[7:0]) +
	( 15'sd 9611) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1753) * $signed(input_fmap_178[7:0]) +
	( 15'sd 11738) * $signed(input_fmap_179[7:0]) +
	( 16'sd 18078) * $signed(input_fmap_180[7:0]) +
	( 15'sd 14702) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26377) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30659) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22909) * $signed(input_fmap_184[7:0]) +
	( 16'sd 31571) * $signed(input_fmap_185[7:0]) +
	( 16'sd 25304) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22982) * $signed(input_fmap_187[7:0]) +
	( 15'sd 11261) * $signed(input_fmap_188[7:0]) +
	( 12'sd 1193) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13547) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31568) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27258) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18943) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27869) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11367) * $signed(input_fmap_196[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18303) * $signed(input_fmap_198[7:0]) +
	( 14'sd 7346) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6730) * $signed(input_fmap_200[7:0]) +
	( 16'sd 25812) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14258) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25284) * $signed(input_fmap_203[7:0]) +
	( 16'sd 31985) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11315) * $signed(input_fmap_205[7:0]) +
	( 15'sd 14424) * $signed(input_fmap_206[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_207[7:0]) +
	( 13'sd 3842) * $signed(input_fmap_208[7:0]) +
	( 16'sd 31960) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10552) * $signed(input_fmap_210[7:0]) +
	( 15'sd 9866) * $signed(input_fmap_211[7:0]) +
	( 15'sd 16228) * $signed(input_fmap_212[7:0]) +
	( 16'sd 21165) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1164) * $signed(input_fmap_214[7:0]) +
	( 14'sd 4429) * $signed(input_fmap_215[7:0]) +
	( 15'sd 9808) * $signed(input_fmap_216[7:0]) +
	( 16'sd 31478) * $signed(input_fmap_217[7:0]) +
	( 16'sd 16800) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3874) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_220[7:0]) +
	( 16'sd 21154) * $signed(input_fmap_221[7:0]) +
	( 15'sd 11491) * $signed(input_fmap_222[7:0]) +
	( 16'sd 20560) * $signed(input_fmap_223[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15136) * $signed(input_fmap_225[7:0]) +
	( 16'sd 25348) * $signed(input_fmap_226[7:0]) +
	( 16'sd 31792) * $signed(input_fmap_227[7:0]) +
	( 16'sd 28247) * $signed(input_fmap_228[7:0]) +
	( 13'sd 2314) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29775) * $signed(input_fmap_230[7:0]) +
	( 16'sd 21393) * $signed(input_fmap_231[7:0]) +
	( 16'sd 32601) * $signed(input_fmap_232[7:0]) +
	( 16'sd 25561) * $signed(input_fmap_233[7:0]) +
	( 16'sd 21325) * $signed(input_fmap_234[7:0]) +
	( 16'sd 28884) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5412) * $signed(input_fmap_236[7:0]) +
	( 15'sd 9694) * $signed(input_fmap_237[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_238[7:0]) +
	( 13'sd 2404) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18895) * $signed(input_fmap_240[7:0]) +
	( 16'sd 27478) * $signed(input_fmap_241[7:0]) +
	( 16'sd 22483) * $signed(input_fmap_242[7:0]) +
	( 15'sd 9889) * $signed(input_fmap_243[7:0]) +
	( 16'sd 23502) * $signed(input_fmap_244[7:0]) +
	( 14'sd 8156) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11408) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20696) * $signed(input_fmap_247[7:0]) +
	( 15'sd 12727) * $signed(input_fmap_248[7:0]) +
	( 11'sd 986) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17534) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13153) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6838) * $signed(input_fmap_252[7:0]) +
	( 12'sd 1616) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2129) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26298) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_170;
assign conv_mac_170 = 
	( 16'sd 25221) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24061) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19865) * $signed(input_fmap_2[7:0]) +
	( 14'sd 8147) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32531) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29008) * $signed(input_fmap_6[7:0]) +
	( 16'sd 30971) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19785) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10014) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19486) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4726) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22648) * $signed(input_fmap_12[7:0]) +
	( 14'sd 7421) * $signed(input_fmap_13[7:0]) +
	( 13'sd 3743) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29423) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15924) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19351) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20861) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10702) * $signed(input_fmap_20[7:0]) +
	( 7'sd 57) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31649) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11609) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12431) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19499) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28521) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27059) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3650) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25240) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21701) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12752) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27078) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1433) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19772) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32017) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19801) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6342) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19603) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24020) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27197) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25379) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29552) * $signed(input_fmap_42[7:0]) +
	( 16'sd 27724) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22269) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7569) * $signed(input_fmap_45[7:0]) +
	( 16'sd 29601) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26469) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16112) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4658) * $signed(input_fmap_50[7:0]) +
	( 14'sd 4287) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19340) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8313) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19025) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17500) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11384) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4410) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18331) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11603) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19538) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28294) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2525) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12209) * $signed(input_fmap_63[7:0]) +
	( 16'sd 30826) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27380) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10512) * $signed(input_fmap_66[7:0]) +
	( 15'sd 16375) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2873) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3899) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23953) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26806) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28218) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24298) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20880) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17376) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12605) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3095) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5849) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23117) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30655) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19849) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10182) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26567) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25017) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25979) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11611) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23839) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22969) * $signed(input_fmap_95[7:0]) +
	( 14'sd 8002) * $signed(input_fmap_96[7:0]) +
	( 16'sd 16881) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29431) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30239) * $signed(input_fmap_99[7:0]) +
	( 15'sd 8494) * $signed(input_fmap_100[7:0]) +
	( 10'sd 305) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24972) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20356) * $signed(input_fmap_103[7:0]) +
	( 16'sd 32620) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30500) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4197) * $signed(input_fmap_106[7:0]) +
	( 16'sd 22542) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19419) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16591) * $signed(input_fmap_109[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12848) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2889) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14563) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27898) * $signed(input_fmap_114[7:0]) +
	( 11'sd 1017) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1995) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28034) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17409) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20786) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9526) * $signed(input_fmap_120[7:0]) +
	( 16'sd 29110) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27837) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5485) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12141) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23634) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28692) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11836) * $signed(input_fmap_127[7:0]) +
	( 15'sd 14809) * $signed(input_fmap_128[7:0]) +
	( 16'sd 18226) * $signed(input_fmap_129[7:0]) +
	( 16'sd 20456) * $signed(input_fmap_130[7:0]) +
	( 16'sd 26177) * $signed(input_fmap_131[7:0]) +
	( 16'sd 26753) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22398) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7194) * $signed(input_fmap_136[7:0]) +
	( 16'sd 29109) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10985) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3168) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28005) * $signed(input_fmap_140[7:0]) +
	( 15'sd 11198) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25454) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26521) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5620) * $signed(input_fmap_144[7:0]) +
	( 15'sd 9796) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15442) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11460) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6647) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12297) * $signed(input_fmap_149[7:0]) +
	( 16'sd 22126) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4725) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2403) * $signed(input_fmap_152[7:0]) +
	( 15'sd 13693) * $signed(input_fmap_153[7:0]) +
	( 16'sd 20317) * $signed(input_fmap_154[7:0]) +
	( 16'sd 32129) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13696) * $signed(input_fmap_156[7:0]) +
	( 16'sd 16821) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1569) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26545) * $signed(input_fmap_159[7:0]) +
	( 16'sd 32092) * $signed(input_fmap_160[7:0]) +
	( 13'sd 3987) * $signed(input_fmap_161[7:0]) +
	( 16'sd 28616) * $signed(input_fmap_162[7:0]) +
	( 14'sd 4459) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11572) * $signed(input_fmap_164[7:0]) +
	( 11'sd 935) * $signed(input_fmap_165[7:0]) +
	( 14'sd 6519) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7223) * $signed(input_fmap_167[7:0]) +
	( 16'sd 30963) * $signed(input_fmap_168[7:0]) +
	( 16'sd 31188) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3998) * $signed(input_fmap_171[7:0]) +
	( 16'sd 30885) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27084) * $signed(input_fmap_173[7:0]) +
	( 16'sd 22561) * $signed(input_fmap_174[7:0]) +
	( 11'sd 782) * $signed(input_fmap_175[7:0]) +
	( 11'sd 701) * $signed(input_fmap_176[7:0]) +
	( 16'sd 28539) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22306) * $signed(input_fmap_178[7:0]) +
	( 14'sd 4623) * $signed(input_fmap_179[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15630) * $signed(input_fmap_181[7:0]) +
	( 12'sd 1448) * $signed(input_fmap_182[7:0]) +
	( 16'sd 20916) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13604) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11632) * $signed(input_fmap_185[7:0]) +
	( 14'sd 7613) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27577) * $signed(input_fmap_187[7:0]) +
	( 14'sd 5130) * $signed(input_fmap_188[7:0]) +
	( 16'sd 28018) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5544) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19903) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28089) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20914) * $signed(input_fmap_193[7:0]) +
	( 16'sd 27360) * $signed(input_fmap_194[7:0]) +
	( 15'sd 9278) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22930) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11432) * $signed(input_fmap_197[7:0]) +
	( 9'sd 136) * $signed(input_fmap_198[7:0]) +
	( 16'sd 18542) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8360) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27971) * $signed(input_fmap_201[7:0]) +
	( 14'sd 4874) * $signed(input_fmap_202[7:0]) +
	( 15'sd 11756) * $signed(input_fmap_203[7:0]) +
	( 16'sd 30179) * $signed(input_fmap_204[7:0]) +
	( 16'sd 25645) * $signed(input_fmap_205[7:0]) +
	( 13'sd 4054) * $signed(input_fmap_206[7:0]) +
	( 15'sd 11876) * $signed(input_fmap_207[7:0]) +
	( 16'sd 21357) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23598) * $signed(input_fmap_209[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30752) * $signed(input_fmap_211[7:0]) +
	( 14'sd 4190) * $signed(input_fmap_212[7:0]) +
	( 10'sd 316) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17395) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9284) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23883) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30260) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8466) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15974) * $signed(input_fmap_219[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1101) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10780) * $signed(input_fmap_222[7:0]) +
	( 15'sd 13973) * $signed(input_fmap_223[7:0]) +
	( 16'sd 18746) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14327) * $signed(input_fmap_225[7:0]) +
	( 16'sd 28350) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22357) * $signed(input_fmap_227[7:0]) +
	( 13'sd 3842) * $signed(input_fmap_228[7:0]) +
	( 16'sd 32023) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_230[7:0]) +
	( 15'sd 16131) * $signed(input_fmap_231[7:0]) +
	( 16'sd 28859) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21650) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5514) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29493) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28223) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29738) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19974) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13971) * $signed(input_fmap_239[7:0]) +
	( 9'sd 184) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25259) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5082) * $signed(input_fmap_242[7:0]) +
	( 16'sd 26773) * $signed(input_fmap_243[7:0]) +
	( 13'sd 3932) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6218) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22246) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11676) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1941) * $signed(input_fmap_248[7:0]) +
	( 16'sd 18295) * $signed(input_fmap_249[7:0]) +
	( 15'sd 13725) * $signed(input_fmap_250[7:0]) +
	( 12'sd 1199) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27029) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24061) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19343) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20021) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_171;
assign conv_mac_171 = 
	( 9'sd 209) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26072) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17549) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17937) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9918) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12496) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27881) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18056) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32729) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29316) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14381) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11310) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5264) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6509) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9817) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16175) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22385) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3046) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23601) * $signed(input_fmap_18[7:0]) +
	( 14'sd 8000) * $signed(input_fmap_19[7:0]) +
	( 15'sd 14277) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13515) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2746) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21795) * $signed(input_fmap_23[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20034) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25777) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1959) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27014) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5729) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21465) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25916) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22512) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23867) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26361) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2256) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21264) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14343) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22433) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21602) * $signed(input_fmap_41[7:0]) +
	( 15'sd 10914) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25807) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20733) * $signed(input_fmap_44[7:0]) +
	( 15'sd 12903) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18163) * $signed(input_fmap_46[7:0]) +
	( 16'sd 23618) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16424) * $signed(input_fmap_49[7:0]) +
	( 9'sd 162) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9213) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25999) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24860) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23169) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31531) * $signed(input_fmap_55[7:0]) +
	( 15'sd 14132) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12473) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16596) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11301) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19982) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3858) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5362) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27361) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4101) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32112) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21570) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26159) * $signed(input_fmap_68[7:0]) +
	( 16'sd 23431) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13180) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8351) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13234) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32732) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16447) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29098) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25575) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13666) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22088) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30832) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9274) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28911) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18527) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22951) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20170) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32562) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9094) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5693) * $signed(input_fmap_90[7:0]) +
	( 8'sd 111) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18913) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2637) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12463) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23361) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2963) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24817) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6718) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28989) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6735) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30962) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12744) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29697) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28257) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32233) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18744) * $signed(input_fmap_109[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_110[7:0]) +
	( 10'sd 382) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10308) * $signed(input_fmap_112[7:0]) +
	( 7'sd 41) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17351) * $signed(input_fmap_114[7:0]) +
	( 15'sd 10689) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8927) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30207) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9246) * $signed(input_fmap_119[7:0]) +
	( 14'sd 5745) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20095) * $signed(input_fmap_121[7:0]) +
	( 16'sd 30001) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13897) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15566) * $signed(input_fmap_124[7:0]) +
	( 14'sd 7815) * $signed(input_fmap_125[7:0]) +
	( 14'sd 8132) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29138) * $signed(input_fmap_127[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_128[7:0]) +
	( 15'sd 8454) * $signed(input_fmap_129[7:0]) +
	( 13'sd 3428) * $signed(input_fmap_130[7:0]) +
	( 15'sd 12045) * $signed(input_fmap_131[7:0]) +
	( 8'sd 117) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32309) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19677) * $signed(input_fmap_135[7:0]) +
	( 16'sd 22319) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4216) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9797) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21599) * $signed(input_fmap_139[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21003) * $signed(input_fmap_142[7:0]) +
	( 15'sd 15861) * $signed(input_fmap_143[7:0]) +
	( 15'sd 15151) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25508) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18428) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9702) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23939) * $signed(input_fmap_148[7:0]) +
	( 15'sd 8244) * $signed(input_fmap_149[7:0]) +
	( 14'sd 6490) * $signed(input_fmap_150[7:0]) +
	( 15'sd 13115) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7991) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14268) * $signed(input_fmap_153[7:0]) +
	( 10'sd 408) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22423) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7147) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11522) * $signed(input_fmap_157[7:0]) +
	( 13'sd 2635) * $signed(input_fmap_158[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_160[7:0]) +
	( 16'sd 26674) * $signed(input_fmap_161[7:0]) +
	( 16'sd 25135) * $signed(input_fmap_162[7:0]) +
	( 16'sd 29897) * $signed(input_fmap_163[7:0]) +
	( 16'sd 31488) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4968) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8572) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17422) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17323) * $signed(input_fmap_169[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11124) * $signed(input_fmap_171[7:0]) +
	( 16'sd 21343) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19208) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19266) * $signed(input_fmap_174[7:0]) +
	( 16'sd 26313) * $signed(input_fmap_175[7:0]) +
	( 16'sd 22988) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29022) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10878) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22062) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15714) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23758) * $signed(input_fmap_181[7:0]) +
	( 14'sd 7469) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17843) * $signed(input_fmap_183[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_184[7:0]) +
	( 16'sd 30045) * $signed(input_fmap_185[7:0]) +
	( 16'sd 27772) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9299) * $signed(input_fmap_187[7:0]) +
	( 15'sd 15300) * $signed(input_fmap_188[7:0]) +
	( 14'sd 4096) * $signed(input_fmap_189[7:0]) +
	( 16'sd 21862) * $signed(input_fmap_190[7:0]) +
	( 15'sd 8996) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27778) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26397) * $signed(input_fmap_193[7:0]) +
	( 16'sd 24675) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1810) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22556) * $signed(input_fmap_197[7:0]) +
	( 16'sd 21520) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5457) * $signed(input_fmap_199[7:0]) +
	( 16'sd 27694) * $signed(input_fmap_200[7:0]) +
	( 16'sd 28702) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19663) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21654) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6045) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5565) * $signed(input_fmap_205[7:0]) +
	( 15'sd 11463) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13575) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22447) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24036) * $signed(input_fmap_209[7:0]) +
	( 16'sd 24259) * $signed(input_fmap_210[7:0]) +
	( 16'sd 31744) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_212[7:0]) +
	( 16'sd 17182) * $signed(input_fmap_213[7:0]) +
	( 15'sd 12674) * $signed(input_fmap_214[7:0]) +
	( 16'sd 31241) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20701) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24755) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31092) * $signed(input_fmap_218[7:0]) +
	( 16'sd 29416) * $signed(input_fmap_219[7:0]) +
	( 15'sd 15371) * $signed(input_fmap_220[7:0]) +
	( 16'sd 22515) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10272) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17794) * $signed(input_fmap_223[7:0]) +
	( 16'sd 20898) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14359) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22272) * $signed(input_fmap_226[7:0]) +
	( 14'sd 7504) * $signed(input_fmap_227[7:0]) +
	( 15'sd 13378) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29952) * $signed(input_fmap_229[7:0]) +
	( 13'sd 2534) * $signed(input_fmap_230[7:0]) +
	( 14'sd 5658) * $signed(input_fmap_231[7:0]) +
	( 16'sd 26714) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1851) * $signed(input_fmap_233[7:0]) +
	( 16'sd 25255) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19739) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30170) * $signed(input_fmap_236[7:0]) +
	( 16'sd 17938) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5156) * $signed(input_fmap_238[7:0]) +
	( 11'sd 699) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10652) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30400) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15833) * $signed(input_fmap_242[7:0]) +
	( 16'sd 26149) * $signed(input_fmap_243[7:0]) +
	( 16'sd 17160) * $signed(input_fmap_244[7:0]) +
	( 11'sd 751) * $signed(input_fmap_245[7:0]) +
	( 13'sd 2628) * $signed(input_fmap_246[7:0]) +
	( 11'sd 561) * $signed(input_fmap_247[7:0]) +
	( 14'sd 6691) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15864) * $signed(input_fmap_249[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_250[7:0]) +
	( 16'sd 23816) * $signed(input_fmap_251[7:0]) +
	( 16'sd 29275) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17361) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31919) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20260) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_172;
assign conv_mac_172 = 
	( 10'sd 317) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10971) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17360) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4456) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19108) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15434) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26915) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31844) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23783) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15946) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15666) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31100) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18525) * $signed(input_fmap_13[7:0]) +
	( 9'sd 218) * $signed(input_fmap_14[7:0]) +
	( 16'sd 16530) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11855) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2652) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3282) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28760) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27703) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27248) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16720) * $signed(input_fmap_22[7:0]) +
	( 16'sd 27448) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2080) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3592) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18064) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21136) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25991) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8843) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15249) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28319) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5380) * $signed(input_fmap_32[7:0]) +
	( 15'sd 14605) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25070) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7113) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21103) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17311) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5894) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20910) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21067) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31456) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24436) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18386) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1508) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19307) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13843) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28255) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14862) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7897) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7346) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31012) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15936) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15379) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5206) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29394) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20215) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14886) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16732) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4420) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7414) * $signed(input_fmap_63[7:0]) +
	( 15'sd 14600) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2737) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8321) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22570) * $signed(input_fmap_67[7:0]) +
	( 16'sd 26239) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18205) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1486) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24148) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14922) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25852) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7122) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6109) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2590) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1219) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8910) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24764) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32489) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3967) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26991) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31670) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29226) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11709) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1650) * $signed(input_fmap_87[7:0]) +
	( 15'sd 15024) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14713) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11610) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9370) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13603) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22200) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7091) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18263) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19414) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25896) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20947) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10040) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10323) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25117) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29903) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31658) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8770) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21575) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15784) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28342) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29445) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29905) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21671) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23540) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4471) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21169) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7185) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18921) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20867) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32011) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9735) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28285) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18319) * $signed(input_fmap_123[7:0]) +
	( 16'sd 25608) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_125[7:0]) +
	( 15'sd 8766) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23156) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_128[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27198) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31861) * $signed(input_fmap_131[7:0]) +
	( 16'sd 28688) * $signed(input_fmap_132[7:0]) +
	( 16'sd 27131) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24735) * $signed(input_fmap_134[7:0]) +
	( 14'sd 7980) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25321) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4673) * $signed(input_fmap_137[7:0]) +
	( 16'sd 21755) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20711) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29458) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10936) * $signed(input_fmap_141[7:0]) +
	( 15'sd 12533) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20493) * $signed(input_fmap_143[7:0]) +
	( 16'sd 26483) * $signed(input_fmap_144[7:0]) +
	( 14'sd 6623) * $signed(input_fmap_145[7:0]) +
	( 15'sd 11905) * $signed(input_fmap_146[7:0]) +
	( 16'sd 32374) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20199) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12280) * $signed(input_fmap_149[7:0]) +
	( 15'sd 14001) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19969) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_152[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25809) * $signed(input_fmap_154[7:0]) +
	( 16'sd 16633) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15267) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25532) * $signed(input_fmap_157[7:0]) +
	( 13'sd 3505) * $signed(input_fmap_158[7:0]) +
	( 14'sd 7453) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24578) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_161[7:0]) +
	( 15'sd 8574) * $signed(input_fmap_162[7:0]) +
	( 16'sd 17085) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19786) * $signed(input_fmap_164[7:0]) +
	( 15'sd 13868) * $signed(input_fmap_165[7:0]) +
	( 16'sd 27634) * $signed(input_fmap_166[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_167[7:0]) +
	( 16'sd 21916) * $signed(input_fmap_168[7:0]) +
	( 16'sd 24890) * $signed(input_fmap_169[7:0]) +
	( 13'sd 3438) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16580) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22247) * $signed(input_fmap_172[7:0]) +
	( 13'sd 2697) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6034) * $signed(input_fmap_174[7:0]) +
	( 16'sd 16774) * $signed(input_fmap_175[7:0]) +
	( 14'sd 8009) * $signed(input_fmap_176[7:0]) +
	( 15'sd 10281) * $signed(input_fmap_177[7:0]) +
	( 16'sd 20878) * $signed(input_fmap_178[7:0]) +
	( 15'sd 14179) * $signed(input_fmap_179[7:0]) +
	( 16'sd 25632) * $signed(input_fmap_180[7:0]) +
	( 16'sd 26105) * $signed(input_fmap_181[7:0]) +
	( 16'sd 24383) * $signed(input_fmap_182[7:0]) +
	( 10'sd 462) * $signed(input_fmap_183[7:0]) +
	( 13'sd 2430) * $signed(input_fmap_184[7:0]) +
	( 16'sd 32660) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17095) * $signed(input_fmap_186[7:0]) +
	( 16'sd 29813) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_189[7:0]) +
	( 16'sd 16939) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23797) * $signed(input_fmap_191[7:0]) +
	( 15'sd 11803) * $signed(input_fmap_192[7:0]) +
	( 16'sd 21389) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21441) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_196[7:0]) +
	( 15'sd 8515) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24416) * $signed(input_fmap_198[7:0]) +
	( 15'sd 8880) * $signed(input_fmap_199[7:0]) +
	( 15'sd 9657) * $signed(input_fmap_200[7:0]) +
	( 14'sd 4637) * $signed(input_fmap_201[7:0]) +
	( 11'sd 844) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6948) * $signed(input_fmap_203[7:0]) +
	( 15'sd 9924) * $signed(input_fmap_204[7:0]) +
	( 14'sd 4990) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31902) * $signed(input_fmap_206[7:0]) +
	( 16'sd 26432) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30567) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7817) * $signed(input_fmap_209[7:0]) +
	( 16'sd 29711) * $signed(input_fmap_210[7:0]) +
	( 15'sd 11136) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24267) * $signed(input_fmap_212[7:0]) +
	( 14'sd 7810) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31611) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1216) * $signed(input_fmap_215[7:0]) +
	( 15'sd 12279) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17574) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13236) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21060) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21977) * $signed(input_fmap_220[7:0]) +
	( 13'sd 3244) * $signed(input_fmap_221[7:0]) +
	( 15'sd 9140) * $signed(input_fmap_222[7:0]) +
	( 15'sd 10063) * $signed(input_fmap_223[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_224[7:0]) +
	( 16'sd 24180) * $signed(input_fmap_225[7:0]) +
	( 16'sd 28299) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13217) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25205) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3645) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7834) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18093) * $signed(input_fmap_231[7:0]) +
	( 14'sd 5354) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23946) * $signed(input_fmap_233[7:0]) +
	( 16'sd 16563) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7675) * $signed(input_fmap_235[7:0]) +
	( 16'sd 20122) * $signed(input_fmap_236[7:0]) +
	( 15'sd 16169) * $signed(input_fmap_237[7:0]) +
	( 14'sd 4133) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12726) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9326) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18460) * $signed(input_fmap_241[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10782) * $signed(input_fmap_243[7:0]) +
	( 16'sd 21255) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5453) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19836) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26398) * $signed(input_fmap_248[7:0]) +
	( 14'sd 5865) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12994) * $signed(input_fmap_250[7:0]) +
	( 10'sd 438) * $signed(input_fmap_251[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_252[7:0]) +
	( 12'sd 1766) * $signed(input_fmap_253[7:0]) +
	( 15'sd 8624) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_173;
assign conv_mac_173 = 
	( 16'sd 29305) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6484) * $signed(input_fmap_1[7:0]) +
	( 16'sd 24931) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29966) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7575) * $signed(input_fmap_4[7:0]) +
	( 10'sd 473) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4967) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12155) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27142) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23590) * $signed(input_fmap_9[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12952) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23664) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11095) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9213) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3186) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18505) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6393) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16738) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9607) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23075) * $signed(input_fmap_22[7:0]) +
	( 16'sd 22390) * $signed(input_fmap_23[7:0]) +
	( 11'sd 869) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30736) * $signed(input_fmap_25[7:0]) +
	( 16'sd 32325) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14493) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31036) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28289) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5363) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28815) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7681) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21178) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18061) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25089) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20800) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32368) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7776) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_39[7:0]) +
	( 15'sd 14722) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1430) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20311) * $signed(input_fmap_42[7:0]) +
	( 14'sd 6276) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30979) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24780) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21967) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7957) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14187) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12630) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28525) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7633) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2367) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17599) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9409) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6188) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30721) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5090) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28364) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11547) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29413) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_62[7:0]) +
	( 15'sd 11134) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32511) * $signed(input_fmap_64[7:0]) +
	( 10'sd 306) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22679) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12056) * $signed(input_fmap_67[7:0]) +
	( 16'sd 32298) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14090) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28725) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4219) * $signed(input_fmap_71[7:0]) +
	( 10'sd 355) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18656) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_74[7:0]) +
	( 16'sd 16924) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12379) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9951) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_78[7:0]) +
	( 16'sd 23277) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17450) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18297) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9029) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21999) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19430) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2298) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19368) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26321) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8210) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25778) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18036) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3690) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26578) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20813) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20875) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29769) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28239) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17568) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6756) * $signed(input_fmap_100[7:0]) +
	( 9'sd 151) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13670) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13298) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9083) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27260) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12939) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24359) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24178) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7288) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27334) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3775) * $signed(input_fmap_111[7:0]) +
	( 15'sd 9413) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11469) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28898) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5529) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20546) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29018) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12155) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14534) * $signed(input_fmap_119[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17890) * $signed(input_fmap_121[7:0]) +
	( 14'sd 6782) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16565) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5372) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2561) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17874) * $signed(input_fmap_128[7:0]) +
	( 15'sd 15028) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_130[7:0]) +
	( 16'sd 25563) * $signed(input_fmap_131[7:0]) +
	( 14'sd 4252) * $signed(input_fmap_132[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_134[7:0]) +
	( 14'sd 8020) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12223) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6267) * $signed(input_fmap_137[7:0]) +
	( 13'sd 2937) * $signed(input_fmap_138[7:0]) +
	( 16'sd 32036) * $signed(input_fmap_139[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_140[7:0]) +
	( 11'sd 770) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14440) * $signed(input_fmap_142[7:0]) +
	( 15'sd 9148) * $signed(input_fmap_143[7:0]) +
	( 15'sd 12494) * $signed(input_fmap_144[7:0]) +
	( 11'sd 822) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14926) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18422) * $signed(input_fmap_147[7:0]) +
	( 16'sd 19204) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12270) * $signed(input_fmap_149[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_150[7:0]) +
	( 16'sd 29797) * $signed(input_fmap_151[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1784) * $signed(input_fmap_153[7:0]) +
	( 16'sd 21684) * $signed(input_fmap_154[7:0]) +
	( 12'sd 1429) * $signed(input_fmap_155[7:0]) +
	( 16'sd 22075) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14275) * $signed(input_fmap_157[7:0]) +
	( 15'sd 14850) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4764) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17820) * $signed(input_fmap_160[7:0]) +
	( 14'sd 8188) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2953) * $signed(input_fmap_162[7:0]) +
	( 14'sd 7881) * $signed(input_fmap_163[7:0]) +
	( 16'sd 32026) * $signed(input_fmap_164[7:0]) +
	( 15'sd 15122) * $signed(input_fmap_165[7:0]) +
	( 15'sd 11800) * $signed(input_fmap_166[7:0]) +
	( 13'sd 3758) * $signed(input_fmap_167[7:0]) +
	( 15'sd 15016) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10780) * $signed(input_fmap_169[7:0]) +
	( 16'sd 25274) * $signed(input_fmap_170[7:0]) +
	( 16'sd 25822) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12174) * $signed(input_fmap_172[7:0]) +
	( 14'sd 4166) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21192) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3677) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15140) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15486) * $signed(input_fmap_178[7:0]) +
	( 15'sd 12729) * $signed(input_fmap_179[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_180[7:0]) +
	( 14'sd 4435) * $signed(input_fmap_181[7:0]) +
	( 12'sd 1180) * $signed(input_fmap_182[7:0]) +
	( 16'sd 25175) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14787) * $signed(input_fmap_184[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_186[7:0]) +
	( 14'sd 6960) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31654) * $signed(input_fmap_188[7:0]) +
	( 16'sd 21525) * $signed(input_fmap_189[7:0]) +
	( 16'sd 32640) * $signed(input_fmap_190[7:0]) +
	( 16'sd 22103) * $signed(input_fmap_191[7:0]) +
	( 15'sd 8295) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23650) * $signed(input_fmap_194[7:0]) +
	( 11'sd 1016) * $signed(input_fmap_195[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25456) * $signed(input_fmap_197[7:0]) +
	( 16'sd 30361) * $signed(input_fmap_198[7:0]) +
	( 15'sd 9224) * $signed(input_fmap_199[7:0]) +
	( 16'sd 28432) * $signed(input_fmap_200[7:0]) +
	( 16'sd 25683) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2811) * $signed(input_fmap_202[7:0]) +
	( 15'sd 14835) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4685) * $signed(input_fmap_204[7:0]) +
	( 16'sd 26933) * $signed(input_fmap_205[7:0]) +
	( 15'sd 16174) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5143) * $signed(input_fmap_207[7:0]) +
	( 16'sd 29829) * $signed(input_fmap_208[7:0]) +
	( 16'sd 30329) * $signed(input_fmap_209[7:0]) +
	( 16'sd 21318) * $signed(input_fmap_210[7:0]) +
	( 15'sd 11120) * $signed(input_fmap_211[7:0]) +
	( 16'sd 22797) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30879) * $signed(input_fmap_214[7:0]) +
	( 10'sd 410) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28570) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10832) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31845) * $signed(input_fmap_218[7:0]) +
	( 16'sd 24258) * $signed(input_fmap_219[7:0]) +
	( 16'sd 17528) * $signed(input_fmap_220[7:0]) +
	( 16'sd 30897) * $signed(input_fmap_221[7:0]) +
	( 15'sd 16311) * $signed(input_fmap_222[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_223[7:0]) +
	( 15'sd 11463) * $signed(input_fmap_224[7:0]) +
	( 16'sd 21164) * $signed(input_fmap_225[7:0]) +
	( 15'sd 9154) * $signed(input_fmap_226[7:0]) +
	( 9'sd 170) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18746) * $signed(input_fmap_228[7:0]) +
	( 10'sd 455) * $signed(input_fmap_229[7:0]) +
	( 10'sd 285) * $signed(input_fmap_230[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_231[7:0]) +
	( 15'sd 13858) * $signed(input_fmap_232[7:0]) +
	( 15'sd 13997) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14079) * $signed(input_fmap_234[7:0]) +
	( 16'sd 23338) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25824) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14139) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_238[7:0]) +
	( 16'sd 28809) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9032) * $signed(input_fmap_240[7:0]) +
	( 15'sd 14506) * $signed(input_fmap_241[7:0]) +
	( 16'sd 25281) * $signed(input_fmap_242[7:0]) +
	( 15'sd 14643) * $signed(input_fmap_243[7:0]) +
	( 14'sd 7352) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12536) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22956) * $signed(input_fmap_246[7:0]) +
	( 16'sd 28781) * $signed(input_fmap_247[7:0]) +
	( 14'sd 7965) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9788) * $signed(input_fmap_249[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6302) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_252[7:0]) +
	( 16'sd 21096) * $signed(input_fmap_253[7:0]) +
	( 14'sd 4677) * $signed(input_fmap_254[7:0]) +
	( 15'sd 13740) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_174;
assign conv_mac_174 = 
	( 15'sd 10612) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29550) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7551) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25536) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26396) * $signed(input_fmap_5[7:0]) +
	( 16'sd 32577) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9019) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22491) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5480) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6661) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10268) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2627) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24331) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27348) * $signed(input_fmap_14[7:0]) +
	( 16'sd 32172) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5658) * $signed(input_fmap_16[7:0]) +
	( 11'sd 944) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3286) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11613) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4876) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3684) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26085) * $signed(input_fmap_23[7:0]) +
	( 15'sd 13891) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1242) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3024) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21720) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20443) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21845) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21824) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1053) * $signed(input_fmap_31[7:0]) +
	( 11'sd 770) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8284) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6313) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12404) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23826) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6480) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27207) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5065) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13271) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18317) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25238) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1299) * $signed(input_fmap_44[7:0]) +
	( 16'sd 16619) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12147) * $signed(input_fmap_47[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_48[7:0]) +
	( 15'sd 10377) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13624) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19914) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24271) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23127) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11769) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19616) * $signed(input_fmap_56[7:0]) +
	( 15'sd 11982) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26679) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6687) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4454) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11787) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16519) * $signed(input_fmap_63[7:0]) +
	( 14'sd 8166) * $signed(input_fmap_64[7:0]) +
	( 11'sd 553) * $signed(input_fmap_65[7:0]) +
	( 14'sd 5192) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24330) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23563) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19194) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2478) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8690) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31879) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12567) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20580) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32242) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7250) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8226) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26523) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22122) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8644) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23125) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15824) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21736) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12136) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9800) * $signed(input_fmap_88[7:0]) +
	( 16'sd 16436) * $signed(input_fmap_89[7:0]) +
	( 15'sd 14767) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26103) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31709) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25647) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12105) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8190) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18504) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15484) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10289) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11622) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8520) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30747) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15019) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32637) * $signed(input_fmap_105[7:0]) +
	( 15'sd 14775) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28004) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18399) * $signed(input_fmap_109[7:0]) +
	( 16'sd 32606) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_111[7:0]) +
	( 16'sd 28540) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11588) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23182) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25962) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31693) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21380) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32269) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3613) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18220) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30170) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22746) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21503) * $signed(input_fmap_127[7:0]) +
	( 16'sd 16508) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31874) * $signed(input_fmap_129[7:0]) +
	( 13'sd 2132) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14223) * $signed(input_fmap_131[7:0]) +
	( 16'sd 28410) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16799) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2416) * $signed(input_fmap_134[7:0]) +
	( 16'sd 25852) * $signed(input_fmap_135[7:0]) +
	( 15'sd 10096) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12545) * $signed(input_fmap_137[7:0]) +
	( 16'sd 28899) * $signed(input_fmap_138[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_139[7:0]) +
	( 16'sd 20132) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10704) * $signed(input_fmap_141[7:0]) +
	( 16'sd 24387) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5898) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13341) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17513) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19026) * $signed(input_fmap_146[7:0]) +
	( 11'sd 556) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21763) * $signed(input_fmap_148[7:0]) +
	( 16'sd 29524) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5184) * $signed(input_fmap_150[7:0]) +
	( 16'sd 16551) * $signed(input_fmap_151[7:0]) +
	( 15'sd 15326) * $signed(input_fmap_152[7:0]) +
	( 14'sd 7791) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11103) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13577) * $signed(input_fmap_155[7:0]) +
	( 16'sd 19134) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31555) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18112) * $signed(input_fmap_158[7:0]) +
	( 12'sd 1996) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21194) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4256) * $signed(input_fmap_161[7:0]) +
	( 15'sd 11218) * $signed(input_fmap_162[7:0]) +
	( 16'sd 21911) * $signed(input_fmap_163[7:0]) +
	( 16'sd 20098) * $signed(input_fmap_164[7:0]) +
	( 16'sd 20090) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8357) * $signed(input_fmap_166[7:0]) +
	( 16'sd 21858) * $signed(input_fmap_167[7:0]) +
	( 16'sd 24565) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21412) * $signed(input_fmap_169[7:0]) +
	( 16'sd 22735) * $signed(input_fmap_170[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14274) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12597) * $signed(input_fmap_173[7:0]) +
	( 15'sd 8487) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15777) * $signed(input_fmap_175[7:0]) +
	( 16'sd 26119) * $signed(input_fmap_176[7:0]) +
	( 15'sd 9718) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9109) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20290) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32704) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18324) * $signed(input_fmap_181[7:0]) +
	( 15'sd 16108) * $signed(input_fmap_182[7:0]) +
	( 16'sd 19213) * $signed(input_fmap_183[7:0]) +
	( 16'sd 29816) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15863) * $signed(input_fmap_185[7:0]) +
	( 16'sd 16525) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1931) * $signed(input_fmap_187[7:0]) +
	( 15'sd 15476) * $signed(input_fmap_188[7:0]) +
	( 16'sd 20899) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31155) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5793) * $signed(input_fmap_191[7:0]) +
	( 16'sd 21011) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10371) * $signed(input_fmap_193[7:0]) +
	( 16'sd 22060) * $signed(input_fmap_194[7:0]) +
	( 16'sd 18397) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12905) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15969) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22570) * $signed(input_fmap_198[7:0]) +
	( 16'sd 27138) * $signed(input_fmap_199[7:0]) +
	( 16'sd 19276) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6942) * $signed(input_fmap_201[7:0]) +
	( 15'sd 12516) * $signed(input_fmap_202[7:0]) +
	( 13'sd 3745) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17329) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12507) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28763) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12777) * $signed(input_fmap_208[7:0]) +
	( 16'sd 30323) * $signed(input_fmap_209[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_210[7:0]) +
	( 16'sd 27953) * $signed(input_fmap_211[7:0]) +
	( 15'sd 15256) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_213[7:0]) +
	( 15'sd 12893) * $signed(input_fmap_214[7:0]) +
	( 16'sd 27406) * $signed(input_fmap_215[7:0]) +
	( 15'sd 9860) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30906) * $signed(input_fmap_217[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_218[7:0]) +
	( 16'sd 29350) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30476) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13350) * $signed(input_fmap_221[7:0]) +
	( 16'sd 30448) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17630) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13161) * $signed(input_fmap_224[7:0]) +
	( 16'sd 19214) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18673) * $signed(input_fmap_226[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25397) * $signed(input_fmap_228[7:0]) +
	( 14'sd 7092) * $signed(input_fmap_229[7:0]) +
	( 12'sd 1153) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31913) * $signed(input_fmap_231[7:0]) +
	( 14'sd 4203) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18456) * $signed(input_fmap_234[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23059) * $signed(input_fmap_236[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12254) * $signed(input_fmap_238[7:0]) +
	( 15'sd 16231) * $signed(input_fmap_239[7:0]) +
	( 16'sd 17530) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21256) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15913) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22146) * $signed(input_fmap_243[7:0]) +
	( 11'sd 666) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5915) * $signed(input_fmap_245[7:0]) +
	( 15'sd 12537) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12634) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4970) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25306) * $signed(input_fmap_249[7:0]) +
	( 16'sd 20263) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_251[7:0]) +
	( 15'sd 11887) * $signed(input_fmap_252[7:0]) +
	( 12'sd 1234) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13212) * $signed(input_fmap_254[7:0]) +
	( 16'sd 18138) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_175;
assign conv_mac_175 = 
	( 12'sd 1994) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2833) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19466) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2216) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11955) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1285) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16954) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32127) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32312) * $signed(input_fmap_8[7:0]) +
	( 15'sd 8527) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6839) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27970) * $signed(input_fmap_11[7:0]) +
	( 16'sd 29530) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17843) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10924) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11357) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9538) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9702) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16715) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9211) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9682) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13149) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12020) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27819) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11401) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3197) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32206) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24421) * $signed(input_fmap_28[7:0]) +
	( 16'sd 27943) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26047) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32137) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17359) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15739) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29615) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32251) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12920) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29054) * $signed(input_fmap_37[7:0]) +
	( 11'sd 923) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6972) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9595) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30237) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3224) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28723) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24668) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31586) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22837) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8987) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16465) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10340) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1822) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6770) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4126) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27306) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16514) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3147) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25328) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18784) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12643) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4460) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11717) * $signed(input_fmap_61[7:0]) +
	( 16'sd 22121) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2205) * $signed(input_fmap_65[7:0]) +
	( 16'sd 31979) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26497) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5156) * $signed(input_fmap_68[7:0]) +
	( 16'sd 17207) * $signed(input_fmap_69[7:0]) +
	( 10'sd 446) * $signed(input_fmap_70[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12551) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7932) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11774) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22333) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3928) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11252) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7674) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30070) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1075) * $signed(input_fmap_80[7:0]) +
	( 11'sd 761) * $signed(input_fmap_81[7:0]) +
	( 15'sd 12431) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31740) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8704) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24008) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23000) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14761) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27107) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29617) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23780) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3369) * $signed(input_fmap_92[7:0]) +
	( 15'sd 9373) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12237) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22410) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22114) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18254) * $signed(input_fmap_97[7:0]) +
	( 14'sd 8086) * $signed(input_fmap_98[7:0]) +
	( 8'sd 118) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17692) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24214) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25472) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9721) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29595) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24695) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18849) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28438) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31387) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18220) * $signed(input_fmap_110[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3176) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18733) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8344) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21502) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11110) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5775) * $signed(input_fmap_117[7:0]) +
	( 11'sd 842) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6479) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11594) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31299) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26453) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15715) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29426) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24825) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30340) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30036) * $signed(input_fmap_127[7:0]) +
	( 16'sd 28026) * $signed(input_fmap_128[7:0]) +
	( 16'sd 18239) * $signed(input_fmap_129[7:0]) +
	( 6'sd 27) * $signed(input_fmap_130[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25583) * $signed(input_fmap_132[7:0]) +
	( 14'sd 4468) * $signed(input_fmap_133[7:0]) +
	( 15'sd 14421) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21634) * $signed(input_fmap_135[7:0]) +
	( 16'sd 20098) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11728) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22179) * $signed(input_fmap_138[7:0]) +
	( 15'sd 9765) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17110) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10353) * $signed(input_fmap_141[7:0]) +
	( 14'sd 7626) * $signed(input_fmap_142[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_143[7:0]) +
	( 16'sd 30496) * $signed(input_fmap_144[7:0]) +
	( 15'sd 9623) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9283) * $signed(input_fmap_146[7:0]) +
	( 14'sd 6597) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20127) * $signed(input_fmap_148[7:0]) +
	( 14'sd 5977) * $signed(input_fmap_149[7:0]) +
	( 15'sd 13616) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17899) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7574) * $signed(input_fmap_152[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_153[7:0]) +
	( 16'sd 18616) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23516) * $signed(input_fmap_155[7:0]) +
	( 16'sd 23022) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29029) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11573) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20917) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31104) * $signed(input_fmap_160[7:0]) +
	( 15'sd 9896) * $signed(input_fmap_161[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2267) * $signed(input_fmap_163[7:0]) +
	( 16'sd 20291) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30813) * $signed(input_fmap_165[7:0]) +
	( 15'sd 10558) * $signed(input_fmap_166[7:0]) +
	( 13'sd 2273) * $signed(input_fmap_167[7:0]) +
	( 15'sd 16001) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17042) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23272) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19417) * $signed(input_fmap_171[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19910) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32596) * $signed(input_fmap_174[7:0]) +
	( 16'sd 24147) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7701) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_177[7:0]) +
	( 15'sd 12906) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3251) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6682) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10933) * $signed(input_fmap_182[7:0]) +
	( 16'sd 24490) * $signed(input_fmap_183[7:0]) +
	( 16'sd 19950) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26094) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2808) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18906) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29232) * $signed(input_fmap_188[7:0]) +
	( 15'sd 8873) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28004) * $signed(input_fmap_190[7:0]) +
	( 14'sd 7178) * $signed(input_fmap_191[7:0]) +
	( 15'sd 8841) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12516) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18417) * $signed(input_fmap_194[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_195[7:0]) +
	( 16'sd 31060) * $signed(input_fmap_196[7:0]) +
	( 16'sd 23446) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19421) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20989) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27294) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14974) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2865) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15512) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6095) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20820) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30327) * $signed(input_fmap_207[7:0]) +
	( 16'sd 27286) * $signed(input_fmap_208[7:0]) +
	( 15'sd 9338) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1580) * $signed(input_fmap_210[7:0]) +
	( 13'sd 2130) * $signed(input_fmap_211[7:0]) +
	( 14'sd 5738) * $signed(input_fmap_212[7:0]) +
	( 16'sd 16716) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31816) * $signed(input_fmap_214[7:0]) +
	( 16'sd 30957) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_216[7:0]) +
	( 16'sd 21543) * $signed(input_fmap_217[7:0]) +
	( 14'sd 4256) * $signed(input_fmap_218[7:0]) +
	( 16'sd 31066) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28939) * $signed(input_fmap_220[7:0]) +
	( 13'sd 4032) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28877) * $signed(input_fmap_222[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_223[7:0]) +
	( 13'sd 2847) * $signed(input_fmap_224[7:0]) +
	( 16'sd 28980) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31541) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9086) * $signed(input_fmap_227[7:0]) +
	( 15'sd 9369) * $signed(input_fmap_228[7:0]) +
	( 15'sd 16009) * $signed(input_fmap_229[7:0]) +
	( 15'sd 9306) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3867) * $signed(input_fmap_231[7:0]) +
	( 16'sd 22893) * $signed(input_fmap_232[7:0]) +
	( 16'sd 30729) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18689) * $signed(input_fmap_234[7:0]) +
	( 16'sd 25719) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23652) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11254) * $signed(input_fmap_237[7:0]) +
	( 16'sd 25147) * $signed(input_fmap_238[7:0]) +
	( 14'sd 4366) * $signed(input_fmap_239[7:0]) +
	( 13'sd 2164) * $signed(input_fmap_240[7:0]) +
	( 16'sd 19496) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17680) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25095) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6306) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1766) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8455) * $signed(input_fmap_247[7:0]) +
	( 16'sd 17822) * $signed(input_fmap_248[7:0]) +
	( 16'sd 20386) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17468) * $signed(input_fmap_250[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_252[7:0]) +
	( 13'sd 4006) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13233) * $signed(input_fmap_254[7:0]) +
	( 13'sd 3806) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_176;
assign conv_mac_176 = 
	( 16'sd 27387) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27601) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25323) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26716) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15014) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2480) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17503) * $signed(input_fmap_6[7:0]) +
	( 14'sd 4555) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31796) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5939) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31273) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18803) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12089) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9364) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3502) * $signed(input_fmap_16[7:0]) +
	( 16'sd 29154) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4784) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1035) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28711) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6300) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11578) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21020) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8195) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28368) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32672) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20972) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3330) * $signed(input_fmap_29[7:0]) +
	( 13'sd 4067) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15330) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10304) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10375) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11684) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22309) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29793) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10571) * $signed(input_fmap_37[7:0]) +
	( 16'sd 28689) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3132) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17713) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18208) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2411) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31767) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10733) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17983) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1309) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10641) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25855) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2360) * $signed(input_fmap_49[7:0]) +
	( 16'sd 24005) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6368) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7871) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10815) * $signed(input_fmap_53[7:0]) +
	( 14'sd 5520) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21925) * $signed(input_fmap_55[7:0]) +
	( 15'sd 11835) * $signed(input_fmap_56[7:0]) +
	( 10'sd 445) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20408) * $signed(input_fmap_58[7:0]) +
	( 15'sd 10667) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17047) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6543) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25134) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23539) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23307) * $signed(input_fmap_65[7:0]) +
	( 15'sd 12019) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10296) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21062) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4773) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1729) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23647) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3025) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11489) * $signed(input_fmap_74[7:0]) +
	( 10'sd 418) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26525) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3814) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24044) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_81[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10174) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20867) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31262) * $signed(input_fmap_85[7:0]) +
	( 8'sd 107) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7539) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16856) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29744) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29600) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18422) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27186) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4398) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2787) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1473) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25230) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7976) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13391) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15396) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17461) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20056) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13563) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10513) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32074) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21652) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23669) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1486) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17172) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12673) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8332) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17637) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19586) * $signed(input_fmap_114[7:0]) +
	( 13'sd 3602) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_116[7:0]) +
	( 16'sd 21756) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15616) * $signed(input_fmap_118[7:0]) +
	( 15'sd 14709) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21914) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13401) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28718) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28602) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28009) * $signed(input_fmap_124[7:0]) +
	( 16'sd 21107) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10888) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28889) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27133) * $signed(input_fmap_130[7:0]) +
	( 15'sd 10473) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14483) * $signed(input_fmap_132[7:0]) +
	( 16'sd 26480) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_134[7:0]) +
	( 13'sd 2886) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31506) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11936) * $signed(input_fmap_137[7:0]) +
	( 16'sd 23789) * $signed(input_fmap_138[7:0]) +
	( 14'sd 6365) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3156) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12007) * $signed(input_fmap_141[7:0]) +
	( 16'sd 26058) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22815) * $signed(input_fmap_145[7:0]) +
	( 16'sd 20464) * $signed(input_fmap_146[7:0]) +
	( 14'sd 5501) * $signed(input_fmap_147[7:0]) +
	( 16'sd 31519) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7795) * $signed(input_fmap_149[7:0]) +
	( 15'sd 16130) * $signed(input_fmap_150[7:0]) +
	( 15'sd 10745) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31085) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10328) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4892) * $signed(input_fmap_154[7:0]) +
	( 12'sd 1533) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10493) * $signed(input_fmap_156[7:0]) +
	( 15'sd 10248) * $signed(input_fmap_157[7:0]) +
	( 15'sd 15841) * $signed(input_fmap_158[7:0]) +
	( 16'sd 18255) * $signed(input_fmap_159[7:0]) +
	( 16'sd 16883) * $signed(input_fmap_160[7:0]) +
	( 15'sd 9992) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27103) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20817) * $signed(input_fmap_163[7:0]) +
	( 15'sd 12207) * $signed(input_fmap_164[7:0]) +
	( 16'sd 24794) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22556) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24048) * $signed(input_fmap_167[7:0]) +
	( 15'sd 16346) * $signed(input_fmap_168[7:0]) +
	( 13'sd 2326) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2184) * $signed(input_fmap_170[7:0]) +
	( 12'sd 1716) * $signed(input_fmap_171[7:0]) +
	( 15'sd 10468) * $signed(input_fmap_172[7:0]) +
	( 16'sd 31493) * $signed(input_fmap_173[7:0]) +
	( 16'sd 30460) * $signed(input_fmap_174[7:0]) +
	( 16'sd 16917) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_176[7:0]) +
	( 16'sd 31384) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9014) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15345) * $signed(input_fmap_179[7:0]) +
	( 14'sd 5335) * $signed(input_fmap_180[7:0]) +
	( 13'sd 2249) * $signed(input_fmap_181[7:0]) +
	( 16'sd 31958) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30577) * $signed(input_fmap_183[7:0]) +
	( 14'sd 5614) * $signed(input_fmap_184[7:0]) +
	( 15'sd 14190) * $signed(input_fmap_185[7:0]) +
	( 15'sd 15004) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25502) * $signed(input_fmap_187[7:0]) +
	( 16'sd 28111) * $signed(input_fmap_188[7:0]) +
	( 15'sd 13606) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4908) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24513) * $signed(input_fmap_191[7:0]) +
	( 15'sd 11730) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30079) * $signed(input_fmap_193[7:0]) +
	( 16'sd 31708) * $signed(input_fmap_194[7:0]) +
	( 15'sd 11287) * $signed(input_fmap_195[7:0]) +
	( 16'sd 29615) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24839) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19815) * $signed(input_fmap_198[7:0]) +
	( 16'sd 25934) * $signed(input_fmap_199[7:0]) +
	( 16'sd 30703) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16825) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31339) * $signed(input_fmap_202[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32297) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5681) * $signed(input_fmap_205[7:0]) +
	( 14'sd 5388) * $signed(input_fmap_206[7:0]) +
	( 16'sd 26952) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_208[7:0]) +
	( 16'sd 27734) * $signed(input_fmap_209[7:0]) +
	( 14'sd 7378) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5723) * $signed(input_fmap_211[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_212[7:0]) +
	( 15'sd 13251) * $signed(input_fmap_213[7:0]) +
	( 16'sd 27708) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10411) * $signed(input_fmap_215[7:0]) +
	( 16'sd 26185) * $signed(input_fmap_216[7:0]) +
	( 16'sd 18655) * $signed(input_fmap_217[7:0]) +
	( 16'sd 16769) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14085) * $signed(input_fmap_219[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_220[7:0]) +
	( 15'sd 14917) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5368) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9631) * $signed(input_fmap_223[7:0]) +
	( 16'sd 16704) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20912) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30388) * $signed(input_fmap_226[7:0]) +
	( 15'sd 15144) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1545) * $signed(input_fmap_228[7:0]) +
	( 14'sd 4284) * $signed(input_fmap_229[7:0]) +
	( 16'sd 26595) * $signed(input_fmap_230[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12848) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_233[7:0]) +
	( 16'sd 25941) * $signed(input_fmap_234[7:0]) +
	( 16'sd 25912) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_236[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_237[7:0]) +
	( 16'sd 21450) * $signed(input_fmap_238[7:0]) +
	( 16'sd 28602) * $signed(input_fmap_239[7:0]) +
	( 15'sd 11789) * $signed(input_fmap_240[7:0]) +
	( 14'sd 4705) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27372) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13712) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20634) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22148) * $signed(input_fmap_245[7:0]) +
	( 14'sd 5805) * $signed(input_fmap_246[7:0]) +
	( 16'sd 23662) * $signed(input_fmap_247[7:0]) +
	( 16'sd 27757) * $signed(input_fmap_248[7:0]) +
	( 16'sd 27539) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_250[7:0]) +
	( 16'sd 24270) * $signed(input_fmap_251[7:0]) +
	( 16'sd 24993) * $signed(input_fmap_252[7:0]) +
	( 15'sd 15674) * $signed(input_fmap_253[7:0]) +
	( 16'sd 27398) * $signed(input_fmap_254[7:0]) +
	( 16'sd 17459) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_177;
assign conv_mac_177 = 
	( 15'sd 13470) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31608) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8612) * $signed(input_fmap_2[7:0]) +
	( 12'sd 1131) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29594) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30223) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13276) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26247) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25987) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2865) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19403) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28029) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10427) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24539) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29739) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21321) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10967) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13076) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8613) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6926) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24809) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19098) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9411) * $signed(input_fmap_23[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25354) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13580) * $signed(input_fmap_26[7:0]) +
	( 14'sd 5803) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25504) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24266) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31094) * $signed(input_fmap_30[7:0]) +
	( 11'sd 996) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3927) * $signed(input_fmap_32[7:0]) +
	( 15'sd 9703) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21775) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2602) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12272) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18862) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19656) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24389) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7275) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2718) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32644) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20413) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21593) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21650) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5329) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21398) * $signed(input_fmap_47[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15280) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13318) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28667) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29684) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13026) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19651) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10043) * $signed(input_fmap_55[7:0]) +
	( 15'sd 9241) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14932) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17644) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10569) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29637) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13443) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13151) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18275) * $signed(input_fmap_64[7:0]) +
	( 16'sd 21613) * $signed(input_fmap_65[7:0]) +
	( 14'sd 7985) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24664) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1384) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8644) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12764) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25224) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7498) * $signed(input_fmap_74[7:0]) +
	( 15'sd 11411) * $signed(input_fmap_75[7:0]) +
	( 15'sd 16250) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28654) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31676) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30353) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20362) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8708) * $signed(input_fmap_82[7:0]) +
	( 9'sd 143) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21155) * $signed(input_fmap_84[7:0]) +
	( 16'sd 28375) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8359) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25507) * $signed(input_fmap_87[7:0]) +
	( 13'sd 3015) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19617) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28591) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27513) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17280) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17963) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14787) * $signed(input_fmap_94[7:0]) +
	( 11'sd 987) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17927) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17774) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30088) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8759) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4316) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4812) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9178) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28313) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19693) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17553) * $signed(input_fmap_105[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29941) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1333) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8790) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18482) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1147) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18193) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15662) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6757) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2399) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10603) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25123) * $signed(input_fmap_117[7:0]) +
	( 14'sd 8165) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16799) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7536) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20366) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20804) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3194) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32044) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29012) * $signed(input_fmap_127[7:0]) +
	( 14'sd 6664) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19567) * $signed(input_fmap_129[7:0]) +
	( 16'sd 27015) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14038) * $signed(input_fmap_131[7:0]) +
	( 14'sd 7247) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11378) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5883) * $signed(input_fmap_134[7:0]) +
	( 7'sd 63) * $signed(input_fmap_135[7:0]) +
	( 15'sd 10267) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26604) * $signed(input_fmap_137[7:0]) +
	( 16'sd 17761) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14993) * $signed(input_fmap_139[7:0]) +
	( 13'sd 2455) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18933) * $signed(input_fmap_141[7:0]) +
	( 16'sd 20109) * $signed(input_fmap_142[7:0]) +
	( 16'sd 32544) * $signed(input_fmap_143[7:0]) +
	( 16'sd 21119) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8989) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9426) * $signed(input_fmap_146[7:0]) +
	( 13'sd 2156) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22521) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27038) * $signed(input_fmap_149[7:0]) +
	( 9'sd 221) * $signed(input_fmap_150[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_151[7:0]) +
	( 16'sd 25299) * $signed(input_fmap_152[7:0]) +
	( 14'sd 5314) * $signed(input_fmap_153[7:0]) +
	( 13'sd 3971) * $signed(input_fmap_154[7:0]) +
	( 16'sd 32239) * $signed(input_fmap_155[7:0]) +
	( 15'sd 9161) * $signed(input_fmap_156[7:0]) +
	( 16'sd 25939) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_158[7:0]) +
	( 15'sd 8856) * $signed(input_fmap_159[7:0]) +
	( 15'sd 10954) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19787) * $signed(input_fmap_161[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15779) * $signed(input_fmap_163[7:0]) +
	( 16'sd 26427) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14738) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13894) * $signed(input_fmap_166[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_167[7:0]) +
	( 16'sd 27817) * $signed(input_fmap_168[7:0]) +
	( 15'sd 13928) * $signed(input_fmap_169[7:0]) +
	( 16'sd 27136) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31617) * $signed(input_fmap_171[7:0]) +
	( 14'sd 5429) * $signed(input_fmap_172[7:0]) +
	( 16'sd 20021) * $signed(input_fmap_173[7:0]) +
	( 10'sd 382) * $signed(input_fmap_174[7:0]) +
	( 16'sd 31029) * $signed(input_fmap_175[7:0]) +
	( 15'sd 9233) * $signed(input_fmap_176[7:0]) +
	( 14'sd 4887) * $signed(input_fmap_177[7:0]) +
	( 14'sd 7978) * $signed(input_fmap_178[7:0]) +
	( 16'sd 24823) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26472) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23165) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12837) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5361) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14615) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26552) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3682) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4657) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23409) * $signed(input_fmap_188[7:0]) +
	( 14'sd 4157) * $signed(input_fmap_189[7:0]) +
	( 15'sd 8652) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_191[7:0]) +
	( 16'sd 26469) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26176) * $signed(input_fmap_193[7:0]) +
	( 15'sd 11495) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_195[7:0]) +
	( 15'sd 8364) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25538) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_198[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_199[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21949) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21719) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6579) * $signed(input_fmap_203[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_204[7:0]) +
	( 15'sd 9543) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2795) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18138) * $signed(input_fmap_207[7:0]) +
	( 16'sd 31971) * $signed(input_fmap_208[7:0]) +
	( 16'sd 28638) * $signed(input_fmap_209[7:0]) +
	( 14'sd 6486) * $signed(input_fmap_210[7:0]) +
	( 15'sd 14405) * $signed(input_fmap_211[7:0]) +
	( 15'sd 10889) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1983) * $signed(input_fmap_213[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25531) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1126) * $signed(input_fmap_216[7:0]) +
	( 15'sd 13422) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31447) * $signed(input_fmap_218[7:0]) +
	( 15'sd 9467) * $signed(input_fmap_219[7:0]) +
	( 14'sd 5182) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28608) * $signed(input_fmap_221[7:0]) +
	( 14'sd 4812) * $signed(input_fmap_222[7:0]) +
	( 14'sd 4201) * $signed(input_fmap_223[7:0]) +
	( 16'sd 26659) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26382) * $signed(input_fmap_225[7:0]) +
	( 14'sd 5488) * $signed(input_fmap_226[7:0]) +
	( 16'sd 25550) * $signed(input_fmap_227[7:0]) +
	( 16'sd 17737) * $signed(input_fmap_228[7:0]) +
	( 13'sd 2584) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30832) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17469) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18967) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24211) * $signed(input_fmap_233[7:0]) +
	( 16'sd 25015) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26398) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28245) * $signed(input_fmap_236[7:0]) +
	( 16'sd 16608) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13860) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9310) * $signed(input_fmap_239[7:0]) +
	( 15'sd 12883) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20809) * $signed(input_fmap_241[7:0]) +
	( 15'sd 14411) * $signed(input_fmap_242[7:0]) +
	( 16'sd 21024) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28010) * $signed(input_fmap_244[7:0]) +
	( 16'sd 16885) * $signed(input_fmap_245[7:0]) +
	( 14'sd 5487) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11676) * $signed(input_fmap_247[7:0]) +
	( 16'sd 31044) * $signed(input_fmap_248[7:0]) +
	( 16'sd 26624) * $signed(input_fmap_249[7:0]) +
	( 16'sd 31288) * $signed(input_fmap_250[7:0]) +
	( 13'sd 3733) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28975) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2634) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19096) * $signed(input_fmap_254[7:0]) +
	( 16'sd 22800) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_178;
assign conv_mac_178 = 
	( 16'sd 24695) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4979) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15025) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_4[7:0]) +
	( 16'sd 28358) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13105) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10361) * $signed(input_fmap_7[7:0]) +
	( 15'sd 10759) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31495) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15091) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31897) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7424) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5228) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5164) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5553) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4578) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16515) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26794) * $signed(input_fmap_21[7:0]) +
	( 9'sd 170) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9033) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12197) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21883) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27273) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6577) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24102) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15794) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16523) * $signed(input_fmap_32[7:0]) +
	( 16'sd 16652) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18035) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31270) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30449) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8805) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29489) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30286) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22377) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28250) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14470) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2410) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22491) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28631) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30634) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12069) * $signed(input_fmap_49[7:0]) +
	( 14'sd 8106) * $signed(input_fmap_50[7:0]) +
	( 13'sd 3717) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17508) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17596) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3144) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7963) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18119) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22620) * $signed(input_fmap_57[7:0]) +
	( 16'sd 22322) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32309) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12036) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6510) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18011) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30324) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9954) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12740) * $signed(input_fmap_67[7:0]) +
	( 16'sd 22701) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7317) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2405) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25133) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14133) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8934) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18158) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6182) * $signed(input_fmap_75[7:0]) +
	( 16'sd 26955) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19280) * $signed(input_fmap_77[7:0]) +
	( 16'sd 25969) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28778) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8032) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19917) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24566) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20830) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8533) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17928) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18941) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5628) * $signed(input_fmap_87[7:0]) +
	( 16'sd 21101) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27593) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16704) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11668) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15738) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27742) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26584) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7398) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2056) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25907) * $signed(input_fmap_98[7:0]) +
	( 15'sd 10831) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2554) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8433) * $signed(input_fmap_101[7:0]) +
	( 15'sd 8421) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25110) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26877) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7041) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5900) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17349) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1728) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7641) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18388) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26196) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14129) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1850) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21893) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23190) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20248) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6037) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24281) * $signed(input_fmap_119[7:0]) +
	( 16'sd 27041) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22359) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29380) * $signed(input_fmap_122[7:0]) +
	( 16'sd 32449) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32227) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29070) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12882) * $signed(input_fmap_126[7:0]) +
	( 15'sd 8862) * $signed(input_fmap_127[7:0]) +
	( 14'sd 6196) * $signed(input_fmap_128[7:0]) +
	( 13'sd 2575) * $signed(input_fmap_129[7:0]) +
	( 16'sd 23969) * $signed(input_fmap_130[7:0]) +
	( 14'sd 7628) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10199) * $signed(input_fmap_132[7:0]) +
	( 16'sd 30809) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2516) * $signed(input_fmap_134[7:0]) +
	( 16'sd 26036) * $signed(input_fmap_135[7:0]) +
	( 16'sd 20540) * $signed(input_fmap_136[7:0]) +
	( 16'sd 28186) * $signed(input_fmap_137[7:0]) +
	( 14'sd 4649) * $signed(input_fmap_138[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_139[7:0]) +
	( 16'sd 31565) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20649) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14545) * $signed(input_fmap_142[7:0]) +
	( 13'sd 3777) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18555) * $signed(input_fmap_144[7:0]) +
	( 15'sd 11917) * $signed(input_fmap_145[7:0]) +
	( 8'sd 109) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9508) * $signed(input_fmap_147[7:0]) +
	( 16'sd 19703) * $signed(input_fmap_148[7:0]) +
	( 14'sd 6463) * $signed(input_fmap_149[7:0]) +
	( 16'sd 32063) * $signed(input_fmap_150[7:0]) +
	( 16'sd 20571) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21870) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31778) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27807) * $signed(input_fmap_155[7:0]) +
	( 15'sd 12021) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15512) * $signed(input_fmap_157[7:0]) +
	( 16'sd 26625) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32457) * $signed(input_fmap_159[7:0]) +
	( 13'sd 3528) * $signed(input_fmap_160[7:0]) +
	( 13'sd 2383) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21282) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2477) * $signed(input_fmap_163[7:0]) +
	( 15'sd 16195) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4189) * $signed(input_fmap_165[7:0]) +
	( 16'sd 29117) * $signed(input_fmap_166[7:0]) +
	( 14'sd 4202) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20012) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14491) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16504) * $signed(input_fmap_171[7:0]) +
	( 15'sd 16253) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18895) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14702) * $signed(input_fmap_174[7:0]) +
	( 16'sd 27431) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21164) * $signed(input_fmap_176[7:0]) +
	( 16'sd 25640) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3368) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28908) * $signed(input_fmap_180[7:0]) +
	( 14'sd 5599) * $signed(input_fmap_181[7:0]) +
	( 7'sd 47) * $signed(input_fmap_182[7:0]) +
	( 14'sd 7779) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24454) * $signed(input_fmap_184[7:0]) +
	( 15'sd 9684) * $signed(input_fmap_185[7:0]) +
	( 15'sd 15011) * $signed(input_fmap_186[7:0]) +
	( 16'sd 32382) * $signed(input_fmap_187[7:0]) +
	( 15'sd 16099) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25439) * $signed(input_fmap_189[7:0]) +
	( 15'sd 14752) * $signed(input_fmap_190[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_191[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20043) * $signed(input_fmap_193[7:0]) +
	( 16'sd 24525) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22067) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_196[7:0]) +
	( 15'sd 12303) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27895) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23932) * $signed(input_fmap_199[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12122) * $signed(input_fmap_201[7:0]) +
	( 16'sd 20487) * $signed(input_fmap_202[7:0]) +
	( 15'sd 14875) * $signed(input_fmap_203[7:0]) +
	( 15'sd 10697) * $signed(input_fmap_204[7:0]) +
	( 15'sd 8485) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3911) * $signed(input_fmap_206[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18851) * $signed(input_fmap_208[7:0]) +
	( 16'sd 16995) * $signed(input_fmap_209[7:0]) +
	( 16'sd 24462) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20891) * $signed(input_fmap_211[7:0]) +
	( 16'sd 31885) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9397) * $signed(input_fmap_213[7:0]) +
	( 16'sd 19198) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9664) * $signed(input_fmap_215[7:0]) +
	( 13'sd 3393) * $signed(input_fmap_216[7:0]) +
	( 16'sd 21454) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21595) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3944) * $signed(input_fmap_219[7:0]) +
	( 15'sd 15627) * $signed(input_fmap_220[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10683) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_223[7:0]) +
	( 16'sd 24054) * $signed(input_fmap_224[7:0]) +
	( 16'sd 25777) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7906) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_227[7:0]) +
	( 15'sd 13413) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8336) * $signed(input_fmap_229[7:0]) +
	( 9'sd 247) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14258) * $signed(input_fmap_231[7:0]) +
	( 16'sd 16713) * $signed(input_fmap_232[7:0]) +
	( 15'sd 8761) * $signed(input_fmap_233[7:0]) +
	( 14'sd 7876) * $signed(input_fmap_234[7:0]) +
	( 16'sd 20089) * $signed(input_fmap_235[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_237[7:0]) +
	( 16'sd 21559) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21627) * $signed(input_fmap_239[7:0]) +
	( 16'sd 30270) * $signed(input_fmap_240[7:0]) +
	( 14'sd 6988) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11667) * $signed(input_fmap_242[7:0]) +
	( 16'sd 18498) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19021) * $signed(input_fmap_244[7:0]) +
	( 15'sd 11508) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31272) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_247[7:0]) +
	( 13'sd 3128) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24712) * $signed(input_fmap_249[7:0]) +
	( 14'sd 6530) * $signed(input_fmap_250[7:0]) +
	( 16'sd 25382) * $signed(input_fmap_251[7:0]) +
	( 12'sd 1954) * $signed(input_fmap_252[7:0]) +
	( 16'sd 16877) * $signed(input_fmap_253[7:0]) +
	( 16'sd 28487) * $signed(input_fmap_254[7:0]) +
	( 16'sd 31760) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_179;
assign conv_mac_179 = 
	( 16'sd 27498) * $signed(input_fmap_0[7:0]) +
	( 16'sd 16837) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14931) * $signed(input_fmap_2[7:0]) +
	( 11'sd 513) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15631) * $signed(input_fmap_4[7:0]) +
	( 14'sd 6186) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29660) * $signed(input_fmap_6[7:0]) +
	( 15'sd 10316) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15139) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18425) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12872) * $signed(input_fmap_10[7:0]) +
	( 11'sd 783) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28070) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12074) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28475) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9445) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20693) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6976) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23530) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20744) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31120) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32259) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29792) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19277) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8560) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14058) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7141) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3068) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27068) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31168) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2961) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28121) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5749) * $signed(input_fmap_32[7:0]) +
	( 16'sd 31117) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23561) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22558) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19593) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25653) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11972) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24644) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19116) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21535) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_43[7:0]) +
	( 16'sd 16937) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26391) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11903) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24509) * $signed(input_fmap_48[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13715) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9636) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20383) * $signed(input_fmap_53[7:0]) +
	( 13'sd 3310) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3282) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23517) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30059) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23900) * $signed(input_fmap_59[7:0]) +
	( 15'sd 12742) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9864) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4677) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16975) * $signed(input_fmap_63[7:0]) +
	( 14'sd 4891) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30768) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30538) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16428) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13009) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3471) * $signed(input_fmap_69[7:0]) +
	( 10'sd 325) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3682) * $signed(input_fmap_71[7:0]) +
	( 16'sd 32551) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4977) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6316) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6724) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11267) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13566) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7710) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9897) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9092) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8359) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17370) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13656) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5520) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26512) * $signed(input_fmap_86[7:0]) +
	( 11'sd 695) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11743) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21629) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13073) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_91[7:0]) +
	( 14'sd 8048) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14001) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15551) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5702) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30961) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22352) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17473) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19889) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25694) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17287) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27532) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7410) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29194) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27219) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28230) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21998) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12287) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23344) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7641) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30536) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16192) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31354) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15682) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9270) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11096) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3609) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24881) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29515) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6613) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5399) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3949) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13882) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17898) * $signed(input_fmap_128[7:0]) +
	( 16'sd 20501) * $signed(input_fmap_129[7:0]) +
	( 13'sd 4051) * $signed(input_fmap_130[7:0]) +
	( 14'sd 7155) * $signed(input_fmap_131[7:0]) +
	( 14'sd 6624) * $signed(input_fmap_132[7:0]) +
	( 15'sd 9604) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25558) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20527) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13539) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9007) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29651) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18413) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_140[7:0]) +
	( 16'sd 28934) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14685) * $signed(input_fmap_142[7:0]) +
	( 15'sd 16120) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22284) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27412) * $signed(input_fmap_145[7:0]) +
	( 13'sd 2863) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8491) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17505) * $signed(input_fmap_148[7:0]) +
	( 9'sd 189) * $signed(input_fmap_149[7:0]) +
	( 11'sd 539) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18887) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21899) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2970) * $signed(input_fmap_153[7:0]) +
	( 15'sd 9287) * $signed(input_fmap_154[7:0]) +
	( 9'sd 244) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15586) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13873) * $signed(input_fmap_157[7:0]) +
	( 13'sd 2161) * $signed(input_fmap_158[7:0]) +
	( 12'sd 1588) * $signed(input_fmap_159[7:0]) +
	( 16'sd 25312) * $signed(input_fmap_160[7:0]) +
	( 15'sd 10467) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27278) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15897) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24751) * $signed(input_fmap_164[7:0]) +
	( 14'sd 6228) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13347) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_167[7:0]) +
	( 15'sd 10372) * $signed(input_fmap_168[7:0]) +
	( 14'sd 4376) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5790) * $signed(input_fmap_170[7:0]) +
	( 14'sd 6891) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1439) * $signed(input_fmap_172[7:0]) +
	( 16'sd 31588) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19196) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5332) * $signed(input_fmap_175[7:0]) +
	( 16'sd 23500) * $signed(input_fmap_176[7:0]) +
	( 16'sd 26383) * $signed(input_fmap_177[7:0]) +
	( 16'sd 16974) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5530) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32379) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30491) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16719) * $signed(input_fmap_182[7:0]) +
	( 16'sd 19102) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13931) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24776) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6426) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1436) * $signed(input_fmap_187[7:0]) +
	( 16'sd 19259) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26939) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5860) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20028) * $signed(input_fmap_191[7:0]) +
	( 16'sd 25696) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9757) * $signed(input_fmap_193[7:0]) +
	( 15'sd 9274) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1534) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6041) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31388) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27908) * $signed(input_fmap_198[7:0]) +
	( 15'sd 15980) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8214) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12703) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8386) * $signed(input_fmap_202[7:0]) +
	( 16'sd 29879) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32101) * $signed(input_fmap_204[7:0]) +
	( 16'sd 19165) * $signed(input_fmap_205[7:0]) +
	( 16'sd 23105) * $signed(input_fmap_206[7:0]) +
	( 15'sd 15172) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30740) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23750) * $signed(input_fmap_209[7:0]) +
	( 16'sd 16811) * $signed(input_fmap_210[7:0]) +
	( 16'sd 31521) * $signed(input_fmap_211[7:0]) +
	( 16'sd 21042) * $signed(input_fmap_212[7:0]) +
	( 16'sd 26821) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31123) * $signed(input_fmap_214[7:0]) +
	( 16'sd 28558) * $signed(input_fmap_215[7:0]) +
	( 14'sd 6810) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25325) * $signed(input_fmap_217[7:0]) +
	( 12'sd 1157) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3132) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14048) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19161) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_223[7:0]) +
	( 16'sd 22548) * $signed(input_fmap_224[7:0]) +
	( 16'sd 30325) * $signed(input_fmap_225[7:0]) +
	( 12'sd 1820) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20729) * $signed(input_fmap_227[7:0]) +
	( 14'sd 6165) * $signed(input_fmap_228[7:0]) +
	( 16'sd 32324) * $signed(input_fmap_229[7:0]) +
	( 15'sd 12305) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7104) * $signed(input_fmap_231[7:0]) +
	( 16'sd 21231) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10578) * $signed(input_fmap_233[7:0]) +
	( 16'sd 17281) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21383) * $signed(input_fmap_235[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_236[7:0]) +
	( 16'sd 17103) * $signed(input_fmap_237[7:0]) +
	( 14'sd 4594) * $signed(input_fmap_238[7:0]) +
	( 16'sd 18710) * $signed(input_fmap_239[7:0]) +
	( 15'sd 12035) * $signed(input_fmap_240[7:0]) +
	( 15'sd 10602) * $signed(input_fmap_241[7:0]) +
	( 14'sd 4757) * $signed(input_fmap_242[7:0]) +
	( 14'sd 5178) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30693) * $signed(input_fmap_244[7:0]) +
	( 15'sd 8804) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17216) * $signed(input_fmap_246[7:0]) +
	( 12'sd 1277) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10660) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3121) * $signed(input_fmap_249[7:0]) +
	( 14'sd 4799) * $signed(input_fmap_250[7:0]) +
	( 16'sd 17496) * $signed(input_fmap_251[7:0]) +
	( 16'sd 16388) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13571) * $signed(input_fmap_253[7:0]) +
	( 15'sd 11373) * $signed(input_fmap_254[7:0]) +
	( 16'sd 31155) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_180;
assign conv_mac_180 = 
	( 15'sd 13948) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29649) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16241) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6511) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8442) * $signed(input_fmap_4[7:0]) +
	( 11'sd 751) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30772) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24513) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18327) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29607) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26389) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28713) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1026) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17879) * $signed(input_fmap_13[7:0]) +
	( 16'sd 23115) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20246) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4177) * $signed(input_fmap_16[7:0]) +
	( 15'sd 9458) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30073) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5731) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5946) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26083) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13483) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16938) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1782) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21300) * $signed(input_fmap_25[7:0]) +
	( 11'sd 791) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6024) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27730) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28112) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1094) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7729) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18120) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28914) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28293) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14410) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21440) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20493) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32067) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22204) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30988) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5507) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18315) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11944) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16301) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31848) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1833) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23616) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16610) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27096) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30142) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2610) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21719) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28613) * $signed(input_fmap_55[7:0]) +
	( 14'sd 6613) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7754) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26837) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2173) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25149) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4272) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12425) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27896) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32512) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27061) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10377) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9902) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30005) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28009) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29393) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_71[7:0]) +
	( 16'sd 27808) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20855) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12283) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24864) * $signed(input_fmap_75[7:0]) +
	( 12'sd 1431) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18004) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30303) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20740) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31095) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18987) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10134) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20959) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3824) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18656) * $signed(input_fmap_87[7:0]) +
	( 10'sd 440) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27683) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8769) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1642) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13413) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_93[7:0]) +
	( 16'sd 27602) * $signed(input_fmap_94[7:0]) +
	( 11'sd 863) * $signed(input_fmap_95[7:0]) +
	( 16'sd 23297) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30413) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15494) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9768) * $signed(input_fmap_99[7:0]) +
	( 11'sd 915) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14308) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21013) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7244) * $signed(input_fmap_103[7:0]) +
	( 16'sd 28429) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29653) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23043) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15501) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2092) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28172) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10657) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12652) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22128) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18749) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20641) * $signed(input_fmap_115[7:0]) +
	( 11'sd 760) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5888) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5605) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5178) * $signed(input_fmap_119[7:0]) +
	( 13'sd 3434) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20464) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26423) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_123[7:0]) +
	( 11'sd 649) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25862) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18974) * $signed(input_fmap_126[7:0]) +
	( 12'sd 2042) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30461) * $signed(input_fmap_128[7:0]) +
	( 16'sd 25446) * $signed(input_fmap_129[7:0]) +
	( 15'sd 16206) * $signed(input_fmap_130[7:0]) +
	( 14'sd 6221) * $signed(input_fmap_131[7:0]) +
	( 15'sd 15876) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29328) * $signed(input_fmap_133[7:0]) +
	( 16'sd 16419) * $signed(input_fmap_134[7:0]) +
	( 14'sd 8183) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21553) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26673) * $signed(input_fmap_137[7:0]) +
	( 14'sd 6208) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21220) * $signed(input_fmap_139[7:0]) +
	( 11'sd 854) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31400) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30984) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1145) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19749) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28898) * $signed(input_fmap_145[7:0]) +
	( 15'sd 11769) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_147[7:0]) +
	( 15'sd 13569) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4702) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21167) * $signed(input_fmap_150[7:0]) +
	( 16'sd 26537) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24574) * $signed(input_fmap_152[7:0]) +
	( 11'sd 807) * $signed(input_fmap_153[7:0]) +
	( 16'sd 17054) * $signed(input_fmap_154[7:0]) +
	( 15'sd 15752) * $signed(input_fmap_155[7:0]) +
	( 16'sd 31530) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29206) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11670) * $signed(input_fmap_158[7:0]) +
	( 16'sd 24676) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11874) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23600) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24161) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22200) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3012) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4676) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31538) * $signed(input_fmap_166[7:0]) +
	( 15'sd 14912) * $signed(input_fmap_167[7:0]) +
	( 16'sd 19737) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20216) * $signed(input_fmap_169[7:0]) +
	( 16'sd 29854) * $signed(input_fmap_170[7:0]) +
	( 16'sd 32224) * $signed(input_fmap_171[7:0]) +
	( 15'sd 15966) * $signed(input_fmap_172[7:0]) +
	( 16'sd 21844) * $signed(input_fmap_173[7:0]) +
	( 11'sd 892) * $signed(input_fmap_174[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15284) * $signed(input_fmap_176[7:0]) +
	( 16'sd 20837) * $signed(input_fmap_177[7:0]) +
	( 13'sd 3416) * $signed(input_fmap_178[7:0]) +
	( 16'sd 30630) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27203) * $signed(input_fmap_180[7:0]) +
	( 16'sd 22284) * $signed(input_fmap_181[7:0]) +
	( 16'sd 31830) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17589) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9503) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27917) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18673) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4282) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1346) * $signed(input_fmap_188[7:0]) +
	( 14'sd 4395) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4527) * $signed(input_fmap_190[7:0]) +
	( 16'sd 16449) * $signed(input_fmap_191[7:0]) +
	( 15'sd 10462) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6612) * $signed(input_fmap_193[7:0]) +
	( 14'sd 7243) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13310) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24924) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26510) * $signed(input_fmap_197[7:0]) +
	( 16'sd 25665) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1477) * $signed(input_fmap_199[7:0]) +
	( 15'sd 15270) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1986) * $signed(input_fmap_201[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_202[7:0]) +
	( 16'sd 16773) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32459) * $signed(input_fmap_204[7:0]) +
	( 15'sd 10549) * $signed(input_fmap_205[7:0]) +
	( 15'sd 11417) * $signed(input_fmap_206[7:0]) +
	( 16'sd 22107) * $signed(input_fmap_207[7:0]) +
	( 16'sd 24495) * $signed(input_fmap_208[7:0]) +
	( 12'sd 1652) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23642) * $signed(input_fmap_210[7:0]) +
	( 16'sd 22782) * $signed(input_fmap_211[7:0]) +
	( 16'sd 27413) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11596) * $signed(input_fmap_213[7:0]) +
	( 16'sd 27027) * $signed(input_fmap_214[7:0]) +
	( 16'sd 21515) * $signed(input_fmap_215[7:0]) +
	( 16'sd 25563) * $signed(input_fmap_216[7:0]) +
	( 16'sd 26659) * $signed(input_fmap_217[7:0]) +
	( 14'sd 7696) * $signed(input_fmap_218[7:0]) +
	( 16'sd 29964) * $signed(input_fmap_219[7:0]) +
	( 15'sd 10026) * $signed(input_fmap_220[7:0]) +
	( 14'sd 4321) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5528) * $signed(input_fmap_222[7:0]) +
	( 16'sd 32374) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6127) * $signed(input_fmap_224[7:0]) +
	( 14'sd 6432) * $signed(input_fmap_225[7:0]) +
	( 13'sd 2828) * $signed(input_fmap_226[7:0]) +
	( 16'sd 16387) * $signed(input_fmap_227[7:0]) +
	( 16'sd 21082) * $signed(input_fmap_228[7:0]) +
	( 16'sd 27248) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15573) * $signed(input_fmap_230[7:0]) +
	( 16'sd 32234) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7104) * $signed(input_fmap_232[7:0]) +
	( 16'sd 25834) * $signed(input_fmap_233[7:0]) +
	( 16'sd 24715) * $signed(input_fmap_234[7:0]) +
	( 13'sd 4059) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28781) * $signed(input_fmap_236[7:0]) +
	( 15'sd 9612) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22391) * $signed(input_fmap_239[7:0]) +
	( 16'sd 30183) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25292) * $signed(input_fmap_241[7:0]) +
	( 15'sd 10552) * $signed(input_fmap_242[7:0]) +
	( 16'sd 20069) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6884) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28368) * $signed(input_fmap_245[7:0]) +
	( 16'sd 26557) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18057) * $signed(input_fmap_247[7:0]) +
	( 15'sd 14591) * $signed(input_fmap_248[7:0]) +
	( 11'sd 929) * $signed(input_fmap_249[7:0]) +
	( 16'sd 20512) * $signed(input_fmap_250[7:0]) +
	( 16'sd 29666) * $signed(input_fmap_251[7:0]) +
	( 16'sd 29117) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27524) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13322) * $signed(input_fmap_254[7:0]) +
	( 16'sd 16805) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_181;
assign conv_mac_181 = 
	( 16'sd 31221) * $signed(input_fmap_0[7:0]) +
	( 16'sd 17773) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7111) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23230) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28943) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30026) * $signed(input_fmap_5[7:0]) +
	( 16'sd 18639) * $signed(input_fmap_6[7:0]) +
	( 16'sd 32097) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24426) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22242) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14491) * $signed(input_fmap_10[7:0]) +
	( 15'sd 15014) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24054) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30886) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12103) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27654) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20981) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30778) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11933) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25726) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12005) * $signed(input_fmap_21[7:0]) +
	( 12'sd 1027) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4959) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25635) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30071) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22566) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22726) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25340) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18939) * $signed(input_fmap_29[7:0]) +
	( 14'sd 6151) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31407) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9114) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28465) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29681) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29212) * $signed(input_fmap_35[7:0]) +
	( 13'sd 3191) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19550) * $signed(input_fmap_37[7:0]) +
	( 16'sd 23531) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8378) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1633) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22681) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3085) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12574) * $signed(input_fmap_43[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30069) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8530) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31454) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25341) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24971) * $signed(input_fmap_49[7:0]) +
	( 16'sd 16641) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26464) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8577) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18852) * $signed(input_fmap_53[7:0]) +
	( 15'sd 16049) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26906) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30474) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7388) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18292) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19395) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20937) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21241) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23608) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29463) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1039) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31636) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26355) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11157) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27198) * $signed(input_fmap_68[7:0]) +
	( 11'sd 607) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11595) * $signed(input_fmap_70[7:0]) +
	( 16'sd 26666) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2064) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30614) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12954) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10351) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13620) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5792) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11882) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7044) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_80[7:0]) +
	( 14'sd 7192) * $signed(input_fmap_81[7:0]) +
	( 16'sd 19300) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10551) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8720) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16728) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31587) * $signed(input_fmap_86[7:0]) +
	( 15'sd 16026) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2854) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27076) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9313) * $signed(input_fmap_90[7:0]) +
	( 16'sd 29467) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_92[7:0]) +
	( 14'sd 5072) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26876) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23842) * $signed(input_fmap_95[7:0]) +
	( 10'sd 486) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9193) * $signed(input_fmap_97[7:0]) +
	( 16'sd 27282) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30984) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27131) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13799) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29427) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27368) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20365) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24999) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16761) * $signed(input_fmap_106[7:0]) +
	( 16'sd 21632) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22763) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1382) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23115) * $signed(input_fmap_110[7:0]) +
	( 16'sd 28405) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6257) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13813) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25625) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5223) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27146) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14401) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17737) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10726) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30445) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17468) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30612) * $signed(input_fmap_123[7:0]) +
	( 14'sd 7636) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31949) * $signed(input_fmap_125[7:0]) +
	( 16'sd 16725) * $signed(input_fmap_126[7:0]) +
	( 13'sd 4012) * $signed(input_fmap_127[7:0]) +
	( 15'sd 14802) * $signed(input_fmap_128[7:0]) +
	( 13'sd 2238) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31416) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13874) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25884) * $signed(input_fmap_132[7:0]) +
	( 16'sd 25429) * $signed(input_fmap_133[7:0]) +
	( 15'sd 12351) * $signed(input_fmap_134[7:0]) +
	( 15'sd 16206) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21959) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25862) * $signed(input_fmap_137[7:0]) +
	( 14'sd 5029) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11053) * $signed(input_fmap_139[7:0]) +
	( 14'sd 7847) * $signed(input_fmap_140[7:0]) +
	( 15'sd 15565) * $signed(input_fmap_141[7:0]) +
	( 16'sd 23893) * $signed(input_fmap_142[7:0]) +
	( 16'sd 18226) * $signed(input_fmap_143[7:0]) +
	( 14'sd 7333) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21446) * $signed(input_fmap_145[7:0]) +
	( 16'sd 25637) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19193) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4909) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7802) * $signed(input_fmap_149[7:0]) +
	( 16'sd 19878) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4738) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23631) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2140) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10308) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12570) * $signed(input_fmap_155[7:0]) +
	( 16'sd 32072) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29676) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28385) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5018) * $signed(input_fmap_159[7:0]) +
	( 11'sd 821) * $signed(input_fmap_160[7:0]) +
	( 15'sd 15093) * $signed(input_fmap_161[7:0]) +
	( 16'sd 20358) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26037) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25687) * $signed(input_fmap_164[7:0]) +
	( 16'sd 18797) * $signed(input_fmap_165[7:0]) +
	( 16'sd 27342) * $signed(input_fmap_166[7:0]) +
	( 16'sd 29436) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20120) * $signed(input_fmap_168[7:0]) +
	( 14'sd 5160) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20417) * $signed(input_fmap_170[7:0]) +
	( 12'sd 1244) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22050) * $signed(input_fmap_172[7:0]) +
	( 10'sd 492) * $signed(input_fmap_173[7:0]) +
	( 16'sd 25959) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25006) * $signed(input_fmap_175[7:0]) +
	( 14'sd 4518) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22624) * $signed(input_fmap_177[7:0]) +
	( 15'sd 16367) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6459) * $signed(input_fmap_179[7:0]) +
	( 16'sd 27105) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28423) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29772) * $signed(input_fmap_182[7:0]) +
	( 16'sd 31801) * $signed(input_fmap_183[7:0]) +
	( 16'sd 28516) * $signed(input_fmap_184[7:0]) +
	( 13'sd 2549) * $signed(input_fmap_185[7:0]) +
	( 15'sd 8394) * $signed(input_fmap_186[7:0]) +
	( 15'sd 8649) * $signed(input_fmap_187[7:0]) +
	( 15'sd 8276) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5265) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5844) * $signed(input_fmap_190[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_191[7:0]) +
	( 15'sd 11871) * $signed(input_fmap_192[7:0]) +
	( 13'sd 2660) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26352) * $signed(input_fmap_194[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_195[7:0]) +
	( 16'sd 18456) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19923) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24538) * $signed(input_fmap_198[7:0]) +
	( 16'sd 18843) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20684) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11050) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2820) * $signed(input_fmap_202[7:0]) +
	( 15'sd 14269) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6481) * $signed(input_fmap_204[7:0]) +
	( 15'sd 14700) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31803) * $signed(input_fmap_206[7:0]) +
	( 16'sd 27632) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18326) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23334) * $signed(input_fmap_209[7:0]) +
	( 14'sd 6163) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12329) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29402) * $signed(input_fmap_212[7:0]) +
	( 15'sd 15941) * $signed(input_fmap_213[7:0]) +
	( 14'sd 5563) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5740) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19191) * $signed(input_fmap_216[7:0]) +
	( 13'sd 3749) * $signed(input_fmap_217[7:0]) +
	( 15'sd 14083) * $signed(input_fmap_218[7:0]) +
	( 16'sd 17374) * $signed(input_fmap_219[7:0]) +
	( 13'sd 3784) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8954) * $signed(input_fmap_223[7:0]) +
	( 15'sd 11691) * $signed(input_fmap_224[7:0]) +
	( 16'sd 23723) * $signed(input_fmap_225[7:0]) +
	( 16'sd 17787) * $signed(input_fmap_226[7:0]) +
	( 16'sd 28278) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31375) * $signed(input_fmap_228[7:0]) +
	( 15'sd 11186) * $signed(input_fmap_229[7:0]) +
	( 15'sd 8558) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1498) * $signed(input_fmap_231[7:0]) +
	( 15'sd 11349) * $signed(input_fmap_232[7:0]) +
	( 15'sd 16014) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3139) * $signed(input_fmap_234[7:0]) +
	( 14'sd 5004) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31195) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_237[7:0]) +
	( 14'sd 8010) * $signed(input_fmap_238[7:0]) +
	( 15'sd 10740) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23583) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15358) * $signed(input_fmap_241[7:0]) +
	( 15'sd 14108) * $signed(input_fmap_242[7:0]) +
	( 12'sd 2024) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30315) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28047) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28990) * $signed(input_fmap_246[7:0]) +
	( 16'sd 22434) * $signed(input_fmap_247[7:0]) +
	( 16'sd 16818) * $signed(input_fmap_248[7:0]) +
	( 15'sd 11520) * $signed(input_fmap_249[7:0]) +
	( 16'sd 16932) * $signed(input_fmap_250[7:0]) +
	( 13'sd 3968) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27586) * $signed(input_fmap_252[7:0]) +
	( 16'sd 26904) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1661) * $signed(input_fmap_254[7:0]) +
	( 15'sd 15558) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_182;
assign conv_mac_182 = 
	( 15'sd 9984) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22956) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26797) * $signed(input_fmap_2[7:0]) +
	( 16'sd 20227) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11625) * $signed(input_fmap_4[7:0]) +
	( 16'sd 16858) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6993) * $signed(input_fmap_6[7:0]) +
	( 15'sd 12492) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1209) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2958) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32688) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10146) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32104) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3579) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13398) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30778) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3124) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23157) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12570) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31589) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12731) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10652) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5942) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25027) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28178) * $signed(input_fmap_24[7:0]) +
	( 16'sd 30959) * $signed(input_fmap_25[7:0]) +
	( 16'sd 31634) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26887) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4859) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5283) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21348) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31472) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_33[7:0]) +
	( 16'sd 22284) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8316) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29391) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32189) * $signed(input_fmap_37[7:0]) +
	( 16'sd 17926) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3301) * $signed(input_fmap_39[7:0]) +
	( 12'sd 1149) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1223) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20253) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5698) * $signed(input_fmap_44[7:0]) +
	( 11'sd 745) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26611) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21076) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28165) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18628) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29288) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15927) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21121) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18434) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27126) * $signed(input_fmap_54[7:0]) +
	( 15'sd 14382) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2169) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3462) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17015) * $signed(input_fmap_59[7:0]) +
	( 13'sd 3569) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31684) * $signed(input_fmap_61[7:0]) +
	( 14'sd 5586) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_63[7:0]) +
	( 16'sd 16493) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31288) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25965) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2643) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4454) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28518) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23166) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2457) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11577) * $signed(input_fmap_73[7:0]) +
	( 11'sd 729) * $signed(input_fmap_74[7:0]) +
	( 15'sd 16205) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19985) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9103) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5147) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13995) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25680) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27536) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22476) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10926) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18129) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7549) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26888) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19637) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27512) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11365) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14024) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10435) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3735) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18650) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11625) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13209) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19557) * $signed(input_fmap_99[7:0]) +
	( 10'sd 470) * $signed(input_fmap_100[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29284) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13743) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30295) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30375) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8238) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9712) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8767) * $signed(input_fmap_110[7:0]) +
	( 11'sd 990) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_112[7:0]) +
	( 16'sd 28274) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18257) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2245) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_117[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3069) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12887) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16398) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18977) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9299) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22146) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20191) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10267) * $signed(input_fmap_127[7:0]) +
	( 16'sd 25342) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28997) * $signed(input_fmap_129[7:0]) +
	( 14'sd 4180) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20219) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11190) * $signed(input_fmap_132[7:0]) +
	( 16'sd 20924) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32642) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32651) * $signed(input_fmap_135[7:0]) +
	( 14'sd 6811) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9387) * $signed(input_fmap_137[7:0]) +
	( 16'sd 16902) * $signed(input_fmap_138[7:0]) +
	( 15'sd 13732) * $signed(input_fmap_139[7:0]) +
	( 16'sd 27672) * $signed(input_fmap_140[7:0]) +
	( 16'sd 26523) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31025) * $signed(input_fmap_142[7:0]) +
	( 16'sd 19831) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2369) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17617) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24745) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27248) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11819) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2904) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31461) * $signed(input_fmap_150[7:0]) +
	( 15'sd 8992) * $signed(input_fmap_151[7:0]) +
	( 15'sd 9391) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31263) * $signed(input_fmap_153[7:0]) +
	( 14'sd 5041) * $signed(input_fmap_154[7:0]) +
	( 15'sd 8284) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18339) * $signed(input_fmap_156[7:0]) +
	( 16'sd 16866) * $signed(input_fmap_157[7:0]) +
	( 14'sd 6381) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27129) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24236) * $signed(input_fmap_160[7:0]) +
	( 10'sd 461) * $signed(input_fmap_161[7:0]) +
	( 12'sd 1273) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2155) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13652) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28722) * $signed(input_fmap_165[7:0]) +
	( 16'sd 17644) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26695) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9517) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11616) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7157) * $signed(input_fmap_170[7:0]) +
	( 15'sd 16239) * $signed(input_fmap_171[7:0]) +
	( 8'sd 91) * $signed(input_fmap_172[7:0]) +
	( 15'sd 9045) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19227) * $signed(input_fmap_174[7:0]) +
	( 15'sd 16068) * $signed(input_fmap_175[7:0]) +
	( 15'sd 14506) * $signed(input_fmap_176[7:0]) +
	( 15'sd 14136) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32526) * $signed(input_fmap_178[7:0]) +
	( 13'sd 4024) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26058) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3975) * $signed(input_fmap_181[7:0]) +
	( 16'sd 24036) * $signed(input_fmap_182[7:0]) +
	( 13'sd 3267) * $signed(input_fmap_183[7:0]) +
	( 15'sd 15744) * $signed(input_fmap_184[7:0]) +
	( 16'sd 31198) * $signed(input_fmap_185[7:0]) +
	( 8'sd 96) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2205) * $signed(input_fmap_187[7:0]) +
	( 14'sd 7905) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11008) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13856) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29704) * $signed(input_fmap_191[7:0]) +
	( 13'sd 3033) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_193[7:0]) +
	( 13'sd 2802) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29845) * $signed(input_fmap_195[7:0]) +
	( 13'sd 2096) * $signed(input_fmap_196[7:0]) +
	( 16'sd 16561) * $signed(input_fmap_197[7:0]) +
	( 16'sd 21386) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29212) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13880) * $signed(input_fmap_200[7:0]) +
	( 16'sd 20781) * $signed(input_fmap_201[7:0]) +
	( 16'sd 20783) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30757) * $signed(input_fmap_203[7:0]) +
	( 16'sd 28556) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29131) * $signed(input_fmap_205[7:0]) +
	( 12'sd 1793) * $signed(input_fmap_206[7:0]) +
	( 14'sd 6554) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_208[7:0]) +
	( 12'sd 1109) * $signed(input_fmap_209[7:0]) +
	( 15'sd 16055) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6320) * $signed(input_fmap_211[7:0]) +
	( 15'sd 13594) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5167) * $signed(input_fmap_213[7:0]) +
	( 16'sd 20405) * $signed(input_fmap_214[7:0]) +
	( 16'sd 32714) * $signed(input_fmap_215[7:0]) +
	( 15'sd 8386) * $signed(input_fmap_216[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21563) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15497) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22912) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13432) * $signed(input_fmap_221[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_222[7:0]) +
	( 14'sd 7655) * $signed(input_fmap_223[7:0]) +
	( 16'sd 18057) * $signed(input_fmap_224[7:0]) +
	( 15'sd 9924) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32224) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9491) * $signed(input_fmap_227[7:0]) +
	( 15'sd 12061) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_229[7:0]) +
	( 10'sd 509) * $signed(input_fmap_230[7:0]) +
	( 11'sd 854) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14055) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15864) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14316) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7576) * $signed(input_fmap_235[7:0]) +
	( 14'sd 7990) * $signed(input_fmap_236[7:0]) +
	( 15'sd 8385) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14885) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26056) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15561) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28574) * $signed(input_fmap_242[7:0]) +
	( 16'sd 23664) * $signed(input_fmap_243[7:0]) +
	( 16'sd 20809) * $signed(input_fmap_244[7:0]) +
	( 16'sd 18257) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28321) * $signed(input_fmap_246[7:0]) +
	( 14'sd 6918) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32020) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12624) * $signed(input_fmap_249[7:0]) +
	( 16'sd 24963) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21572) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12014) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3911) * $signed(input_fmap_253[7:0]) +
	( 16'sd 25841) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5491) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_183;
assign conv_mac_183 = 
	( 16'sd 26671) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20260) * $signed(input_fmap_1[7:0]) +
	( 15'sd 16188) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24823) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13227) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18329) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27505) * $signed(input_fmap_6[7:0]) +
	( 10'sd 510) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28825) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10869) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5534) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26282) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10227) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10384) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11367) * $signed(input_fmap_14[7:0]) +
	( 16'sd 27574) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2724) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25050) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26874) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15811) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5954) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10474) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23531) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5849) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27340) * $signed(input_fmap_25[7:0]) +
	( 11'sd 939) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31125) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4336) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1388) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3905) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29492) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28597) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30057) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18629) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4614) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15731) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24445) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9203) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21190) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32310) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3528) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17126) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8098) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15790) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11581) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20204) * $signed(input_fmap_47[7:0]) +
	( 14'sd 4656) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9456) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28882) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26684) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2115) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4470) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13986) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15402) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29489) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15916) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10023) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2828) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25374) * $signed(input_fmap_60[7:0]) +
	( 16'sd 26081) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15382) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18296) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12185) * $signed(input_fmap_65[7:0]) +
	( 13'sd 2645) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19917) * $signed(input_fmap_67[7:0]) +
	( 11'sd 581) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29298) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5128) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2953) * $signed(input_fmap_71[7:0]) +
	( 15'sd 14037) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29797) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7003) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29178) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17304) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10852) * $signed(input_fmap_78[7:0]) +
	( 16'sd 26957) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14545) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26221) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8414) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15209) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25300) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17520) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8736) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11539) * $signed(input_fmap_87[7:0]) +
	( 10'sd 472) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17824) * $signed(input_fmap_89[7:0]) +
	( 16'sd 27941) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28911) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27373) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12191) * $signed(input_fmap_94[7:0]) +
	( 13'sd 2431) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9655) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31704) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24096) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12436) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23528) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_102[7:0]) +
	( 14'sd 7688) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16938) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11695) * $signed(input_fmap_105[7:0]) +
	( 11'sd 612) * $signed(input_fmap_106[7:0]) +
	( 11'sd 672) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_109[7:0]) +
	( 15'sd 8474) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20987) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25900) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15125) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11078) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13281) * $signed(input_fmap_115[7:0]) +
	( 6'sd 20) * $signed(input_fmap_116[7:0]) +
	( 15'sd 12001) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4868) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26890) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18714) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24758) * $signed(input_fmap_121[7:0]) +
	( 15'sd 14879) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20122) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20018) * $signed(input_fmap_124[7:0]) +
	( 16'sd 17086) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27632) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19621) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8362) * $signed(input_fmap_128[7:0]) +
	( 16'sd 26086) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22515) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31632) * $signed(input_fmap_131[7:0]) +
	( 16'sd 22961) * $signed(input_fmap_132[7:0]) +
	( 15'sd 14772) * $signed(input_fmap_133[7:0]) +
	( 14'sd 7586) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19799) * $signed(input_fmap_135[7:0]) +
	( 13'sd 3042) * $signed(input_fmap_136[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_137[7:0]) +
	( 16'sd 25874) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28104) * $signed(input_fmap_139[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22344) * $signed(input_fmap_141[7:0]) +
	( 10'sd 479) * $signed(input_fmap_142[7:0]) +
	( 13'sd 2333) * $signed(input_fmap_143[7:0]) +
	( 16'sd 23740) * $signed(input_fmap_144[7:0]) +
	( 16'sd 19368) * $signed(input_fmap_145[7:0]) +
	( 15'sd 10538) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18571) * $signed(input_fmap_147[7:0]) +
	( 16'sd 19843) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27337) * $signed(input_fmap_149[7:0]) +
	( 16'sd 24780) * $signed(input_fmap_150[7:0]) +
	( 16'sd 25470) * $signed(input_fmap_151[7:0]) +
	( 13'sd 3541) * $signed(input_fmap_152[7:0]) +
	( 15'sd 15395) * $signed(input_fmap_153[7:0]) +
	( 15'sd 14557) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12494) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18063) * $signed(input_fmap_156[7:0]) +
	( 9'sd 195) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20312) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27754) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6720) * $signed(input_fmap_160[7:0]) +
	( 16'sd 27615) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_162[7:0]) +
	( 14'sd 5997) * $signed(input_fmap_163[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_165[7:0]) +
	( 15'sd 16316) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26087) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20968) * $signed(input_fmap_169[7:0]) +
	( 15'sd 13624) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18113) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1467) * $signed(input_fmap_172[7:0]) +
	( 15'sd 14765) * $signed(input_fmap_173[7:0]) +
	( 12'sd 1046) * $signed(input_fmap_174[7:0]) +
	( 15'sd 11264) * $signed(input_fmap_175[7:0]) +
	( 16'sd 24941) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19185) * $signed(input_fmap_177[7:0]) +
	( 15'sd 9833) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22444) * $signed(input_fmap_179[7:0]) +
	( 16'sd 25562) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11076) * $signed(input_fmap_181[7:0]) +
	( 16'sd 22995) * $signed(input_fmap_182[7:0]) +
	( 16'sd 18549) * $signed(input_fmap_183[7:0]) +
	( 15'sd 10454) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6701) * $signed(input_fmap_185[7:0]) +
	( 16'sd 22694) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9235) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2521) * $signed(input_fmap_188[7:0]) +
	( 16'sd 18671) * $signed(input_fmap_189[7:0]) +
	( 15'sd 9579) * $signed(input_fmap_190[7:0]) +
	( 16'sd 21162) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28395) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5326) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23200) * $signed(input_fmap_194[7:0]) +
	( 15'sd 12168) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22105) * $signed(input_fmap_197[7:0]) +
	( 16'sd 28700) * $signed(input_fmap_198[7:0]) +
	( 16'sd 31963) * $signed(input_fmap_199[7:0]) +
	( 16'sd 24735) * $signed(input_fmap_200[7:0]) +
	( 16'sd 30966) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19013) * $signed(input_fmap_202[7:0]) +
	( 15'sd 9562) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6424) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15345) * $signed(input_fmap_205[7:0]) +
	( 16'sd 18470) * $signed(input_fmap_206[7:0]) +
	( 16'sd 27847) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8865) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26635) * $signed(input_fmap_209[7:0]) +
	( 15'sd 12653) * $signed(input_fmap_210[7:0]) +
	( 16'sd 18970) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26008) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12416) * $signed(input_fmap_213[7:0]) +
	( 16'sd 27411) * $signed(input_fmap_214[7:0]) +
	( 16'sd 28652) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23984) * $signed(input_fmap_216[7:0]) +
	( 13'sd 2531) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26427) * $signed(input_fmap_218[7:0]) +
	( 16'sd 30690) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21693) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5106) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14489) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8364) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12224) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2538) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22109) * $signed(input_fmap_226[7:0]) +
	( 16'sd 28741) * $signed(input_fmap_227[7:0]) +
	( 16'sd 30939) * $signed(input_fmap_228[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27462) * $signed(input_fmap_230[7:0]) +
	( 16'sd 21477) * $signed(input_fmap_231[7:0]) +
	( 16'sd 25327) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_233[7:0]) +
	( 16'sd 25457) * $signed(input_fmap_234[7:0]) +
	( 14'sd 8075) * $signed(input_fmap_235[7:0]) +
	( 16'sd 32307) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11256) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12552) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23320) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25570) * $signed(input_fmap_240[7:0]) +
	( 13'sd 2438) * $signed(input_fmap_241[7:0]) +
	( 15'sd 14523) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28925) * $signed(input_fmap_243[7:0]) +
	( 13'sd 3064) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2226) * $signed(input_fmap_245[7:0]) +
	( 14'sd 4705) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17467) * $signed(input_fmap_247[7:0]) +
	( 15'sd 15817) * $signed(input_fmap_248[7:0]) +
	( 14'sd 8115) * $signed(input_fmap_249[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_250[7:0]) +
	( 9'sd 164) * $signed(input_fmap_251[7:0]) +
	( 15'sd 16135) * $signed(input_fmap_252[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_253[7:0]) +
	( 16'sd 30148) * $signed(input_fmap_254[7:0]) +
	( 16'sd 18735) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_184;
assign conv_mac_184 = 
	( 11'sd 975) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8258) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8822) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17015) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14425) * $signed(input_fmap_6[7:0]) +
	( 15'sd 16365) * $signed(input_fmap_7[7:0]) +
	( 16'sd 31325) * $signed(input_fmap_8[7:0]) +
	( 15'sd 14820) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24034) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19336) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7194) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28633) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13794) * $signed(input_fmap_14[7:0]) +
	( 16'sd 26561) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10537) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30515) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4962) * $signed(input_fmap_18[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_20[7:0]) +
	( 16'sd 28169) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11148) * $signed(input_fmap_22[7:0]) +
	( 15'sd 13879) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10337) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4308) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30675) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1052) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13630) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17931) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13059) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2986) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21959) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5842) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25867) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27800) * $signed(input_fmap_36[7:0]) +
	( 15'sd 16353) * $signed(input_fmap_37[7:0]) +
	( 16'sd 21466) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30048) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22801) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14745) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2658) * $signed(input_fmap_43[7:0]) +
	( 14'sd 8081) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20652) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8518) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2978) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22216) * $signed(input_fmap_48[7:0]) +
	( 16'sd 22917) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6955) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12880) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19566) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28823) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26129) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26892) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15257) * $signed(input_fmap_57[7:0]) +
	( 14'sd 5051) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18212) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20967) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17712) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20653) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_63[7:0]) +
	( 9'sd 245) * $signed(input_fmap_64[7:0]) +
	( 16'sd 27896) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19999) * $signed(input_fmap_66[7:0]) +
	( 16'sd 18843) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30786) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32158) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2573) * $signed(input_fmap_70[7:0]) +
	( 15'sd 15058) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20098) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_73[7:0]) +
	( 10'sd 419) * $signed(input_fmap_74[7:0]) +
	( 16'sd 28766) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16961) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2846) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17620) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13656) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19098) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8514) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21413) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27951) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19674) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18908) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29419) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32096) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7184) * $signed(input_fmap_89[7:0]) +
	( 16'sd 30767) * $signed(input_fmap_90[7:0]) +
	( 9'sd 226) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31399) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11943) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15198) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3550) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6400) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18857) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27176) * $signed(input_fmap_99[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22507) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3698) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14783) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25087) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12897) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28639) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26153) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28167) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24720) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30988) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30337) * $signed(input_fmap_111[7:0]) +
	( 11'sd 714) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29650) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4329) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30128) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32407) * $signed(input_fmap_116[7:0]) +
	( 12'sd 1764) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12848) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17779) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32535) * $signed(input_fmap_120[7:0]) +
	( 15'sd 13942) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26274) * $signed(input_fmap_122[7:0]) +
	( 16'sd 29644) * $signed(input_fmap_123[7:0]) +
	( 14'sd 4468) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28902) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19944) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20606) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23516) * $signed(input_fmap_128[7:0]) +
	( 16'sd 32561) * $signed(input_fmap_129[7:0]) +
	( 13'sd 3519) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31357) * $signed(input_fmap_131[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_132[7:0]) +
	( 15'sd 13623) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5811) * $signed(input_fmap_134[7:0]) +
	( 14'sd 4798) * $signed(input_fmap_135[7:0]) +
	( 14'sd 4096) * $signed(input_fmap_136[7:0]) +
	( 15'sd 10435) * $signed(input_fmap_137[7:0]) +
	( 16'sd 23672) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31901) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17617) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5459) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27262) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1294) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13891) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26820) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14145) * $signed(input_fmap_147[7:0]) +
	( 16'sd 16969) * $signed(input_fmap_148[7:0]) +
	( 15'sd 10770) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18220) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_151[7:0]) +
	( 16'sd 25106) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14613) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7030) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12347) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17980) * $signed(input_fmap_156[7:0]) +
	( 9'sd 245) * $signed(input_fmap_157[7:0]) +
	( 15'sd 10825) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21260) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26698) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4206) * $signed(input_fmap_161[7:0]) +
	( 10'sd 504) * $signed(input_fmap_162[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3168) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2505) * $signed(input_fmap_165[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13040) * $signed(input_fmap_167[7:0]) +
	( 16'sd 30745) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6861) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7435) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9831) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19529) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6805) * $signed(input_fmap_174[7:0]) +
	( 16'sd 31618) * $signed(input_fmap_175[7:0]) +
	( 16'sd 22661) * $signed(input_fmap_176[7:0]) +
	( 16'sd 21861) * $signed(input_fmap_177[7:0]) +
	( 11'sd 610) * $signed(input_fmap_178[7:0]) +
	( 15'sd 15666) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3943) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15469) * $signed(input_fmap_181[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_182[7:0]) +
	( 16'sd 20406) * $signed(input_fmap_183[7:0]) +
	( 16'sd 21260) * $signed(input_fmap_184[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_185[7:0]) +
	( 16'sd 30600) * $signed(input_fmap_186[7:0]) +
	( 15'sd 12573) * $signed(input_fmap_187[7:0]) +
	( 16'sd 22594) * $signed(input_fmap_188[7:0]) +
	( 16'sd 32644) * $signed(input_fmap_189[7:0]) +
	( 14'sd 6131) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24803) * $signed(input_fmap_192[7:0]) +
	( 13'sd 3583) * $signed(input_fmap_193[7:0]) +
	( 16'sd 17420) * $signed(input_fmap_194[7:0]) +
	( 16'sd 19048) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5228) * $signed(input_fmap_196[7:0]) +
	( 14'sd 4301) * $signed(input_fmap_197[7:0]) +
	( 14'sd 7631) * $signed(input_fmap_198[7:0]) +
	( 15'sd 8268) * $signed(input_fmap_199[7:0]) +
	( 15'sd 11160) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9997) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5541) * $signed(input_fmap_203[7:0]) +
	( 16'sd 18001) * $signed(input_fmap_204[7:0]) +
	( 16'sd 19424) * $signed(input_fmap_205[7:0]) +
	( 15'sd 13175) * $signed(input_fmap_206[7:0]) +
	( 16'sd 16686) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30990) * $signed(input_fmap_208[7:0]) +
	( 15'sd 12297) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18139) * $signed(input_fmap_210[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12997) * $signed(input_fmap_212[7:0]) +
	( 16'sd 21462) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23907) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6269) * $signed(input_fmap_215[7:0]) +
	( 16'sd 30665) * $signed(input_fmap_216[7:0]) +
	( 16'sd 23532) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10543) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19208) * $signed(input_fmap_219[7:0]) +
	( 14'sd 7215) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25404) * $signed(input_fmap_221[7:0]) +
	( 16'sd 30062) * $signed(input_fmap_222[7:0]) +
	( 16'sd 21444) * $signed(input_fmap_223[7:0]) +
	( 16'sd 28023) * $signed(input_fmap_224[7:0]) +
	( 15'sd 9409) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7721) * $signed(input_fmap_226[7:0]) +
	( 16'sd 19398) * $signed(input_fmap_227[7:0]) +
	( 15'sd 15806) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17040) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15375) * $signed(input_fmap_230[7:0]) +
	( 16'sd 27132) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18589) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10947) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3332) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11809) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10331) * $signed(input_fmap_237[7:0]) +
	( 10'sd 502) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21852) * $signed(input_fmap_239[7:0]) +
	( 16'sd 27800) * $signed(input_fmap_240[7:0]) +
	( 16'sd 24100) * $signed(input_fmap_241[7:0]) +
	( 11'sd 735) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31422) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1269) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6189) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9849) * $signed(input_fmap_246[7:0]) +
	( 16'sd 16813) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21845) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24963) * $signed(input_fmap_249[7:0]) +
	( 10'sd 424) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22810) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26859) * $signed(input_fmap_252[7:0]) +
	( 13'sd 2110) * $signed(input_fmap_253[7:0]) +
	( 16'sd 18701) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23266) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_185;
assign conv_mac_185 = 
	( 16'sd 21920) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30282) * $signed(input_fmap_1[7:0]) +
	( 15'sd 10440) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25588) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7620) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21959) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27552) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25398) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12617) * $signed(input_fmap_9[7:0]) +
	( 11'sd 544) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22489) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1838) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20282) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16264) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2978) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28237) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18219) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24853) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13746) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14959) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7122) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17957) * $signed(input_fmap_25[7:0]) +
	( 9'sd 180) * $signed(input_fmap_26[7:0]) +
	( 15'sd 15260) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3918) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16189) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1108) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13585) * $signed(input_fmap_32[7:0]) +
	( 5'sd 9) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14819) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21733) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6506) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7381) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31334) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19459) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31717) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16390) * $signed(input_fmap_41[7:0]) +
	( 13'sd 4030) * $signed(input_fmap_42[7:0]) +
	( 15'sd 9505) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5856) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27564) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4138) * $signed(input_fmap_46[7:0]) +
	( 10'sd 486) * $signed(input_fmap_47[7:0]) +
	( 15'sd 11430) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31329) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15796) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6435) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16215) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1930) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7106) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30267) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19026) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31148) * $signed(input_fmap_58[7:0]) +
	( 10'sd 367) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5571) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12055) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14048) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3808) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31486) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14058) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19061) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11468) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12455) * $signed(input_fmap_70[7:0]) +
	( 15'sd 12909) * $signed(input_fmap_71[7:0]) +
	( 13'sd 4091) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3600) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30312) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24918) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26992) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11741) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5431) * $signed(input_fmap_79[7:0]) +
	( 16'sd 25210) * $signed(input_fmap_80[7:0]) +
	( 14'sd 4147) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29077) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8228) * $signed(input_fmap_83[7:0]) +
	( 16'sd 25932) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30574) * $signed(input_fmap_85[7:0]) +
	( 16'sd 30899) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10136) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20371) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10182) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25195) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4520) * $signed(input_fmap_91[7:0]) +
	( 16'sd 29305) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20511) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25143) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12851) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27447) * $signed(input_fmap_96[7:0]) +
	( 16'sd 26890) * $signed(input_fmap_97[7:0]) +
	( 10'sd 355) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17340) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27651) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30549) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11582) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5333) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15833) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7450) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16389) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9222) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28306) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18683) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26872) * $signed(input_fmap_111[7:0]) +
	( 14'sd 7541) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19629) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4843) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20154) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27129) * $signed(input_fmap_116[7:0]) +
	( 15'sd 11165) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22726) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31990) * $signed(input_fmap_119[7:0]) +
	( 16'sd 19146) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25172) * $signed(input_fmap_121[7:0]) +
	( 16'sd 20937) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24564) * $signed(input_fmap_123[7:0]) +
	( 16'sd 26483) * $signed(input_fmap_124[7:0]) +
	( 10'sd 281) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28833) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20716) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8413) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10640) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30348) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_131[7:0]) +
	( 16'sd 32475) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12716) * $signed(input_fmap_136[7:0]) +
	( 16'sd 17015) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22883) * $signed(input_fmap_138[7:0]) +
	( 14'sd 4366) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30534) * $signed(input_fmap_140[7:0]) +
	( 16'sd 17661) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11455) * $signed(input_fmap_142[7:0]) +
	( 16'sd 30892) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3231) * $signed(input_fmap_144[7:0]) +
	( 16'sd 32008) * $signed(input_fmap_145[7:0]) +
	( 14'sd 4165) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8404) * $signed(input_fmap_147[7:0]) +
	( 12'sd 1469) * $signed(input_fmap_148[7:0]) +
	( 14'sd 5760) * $signed(input_fmap_149[7:0]) +
	( 15'sd 13170) * $signed(input_fmap_150[7:0]) +
	( 13'sd 2190) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16679) * $signed(input_fmap_152[7:0]) +
	( 15'sd 15412) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6572) * $signed(input_fmap_154[7:0]) +
	( 13'sd 3481) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7578) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14829) * $signed(input_fmap_157[7:0]) +
	( 16'sd 19778) * $signed(input_fmap_158[7:0]) +
	( 16'sd 24527) * $signed(input_fmap_159[7:0]) +
	( 15'sd 8950) * $signed(input_fmap_160[7:0]) +
	( 15'sd 10347) * $signed(input_fmap_161[7:0]) +
	( 14'sd 6281) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24448) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8798) * $signed(input_fmap_164[7:0]) +
	( 13'sd 3113) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13875) * $signed(input_fmap_166[7:0]) +
	( 15'sd 14811) * $signed(input_fmap_167[7:0]) +
	( 16'sd 22223) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25625) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24925) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30624) * $signed(input_fmap_171[7:0]) +
	( 15'sd 13767) * $signed(input_fmap_172[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_173[7:0]) +
	( 16'sd 24389) * $signed(input_fmap_174[7:0]) +
	( 15'sd 12297) * $signed(input_fmap_175[7:0]) +
	( 16'sd 27159) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29634) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2101) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25687) * $signed(input_fmap_179[7:0]) +
	( 16'sd 30672) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_181[7:0]) +
	( 16'sd 24937) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2479) * $signed(input_fmap_183[7:0]) +
	( 14'sd 6276) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11304) * $signed(input_fmap_185[7:0]) +
	( 15'sd 14242) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28713) * $signed(input_fmap_187[7:0]) +
	( 15'sd 14437) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7383) * $signed(input_fmap_189[7:0]) +
	( 16'sd 23976) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31967) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19222) * $signed(input_fmap_192[7:0]) +
	( 16'sd 31433) * $signed(input_fmap_193[7:0]) +
	( 16'sd 19295) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25643) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19998) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10663) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5200) * $signed(input_fmap_198[7:0]) +
	( 14'sd 4175) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13246) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18929) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24689) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14954) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1952) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12942) * $signed(input_fmap_206[7:0]) +
	( 11'sd 566) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4832) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13776) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9176) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26433) * $signed(input_fmap_211[7:0]) +
	( 14'sd 6740) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11648) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28140) * $signed(input_fmap_214[7:0]) +
	( 16'sd 30482) * $signed(input_fmap_215[7:0]) +
	( 14'sd 7492) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26731) * $signed(input_fmap_218[7:0]) +
	( 16'sd 23370) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25570) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6490) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28343) * $signed(input_fmap_222[7:0]) +
	( 16'sd 27635) * $signed(input_fmap_223[7:0]) +
	( 15'sd 11979) * $signed(input_fmap_224[7:0]) +
	( 14'sd 6606) * $signed(input_fmap_225[7:0]) +
	( 7'sd 45) * $signed(input_fmap_226[7:0]) +
	( 16'sd 25715) * $signed(input_fmap_227[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_228[7:0]) +
	( 15'sd 12426) * $signed(input_fmap_229[7:0]) +
	( 16'sd 17919) * $signed(input_fmap_230[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_231[7:0]) +
	( 16'sd 22303) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3439) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13034) * $signed(input_fmap_234[7:0]) +
	( 16'sd 20288) * $signed(input_fmap_235[7:0]) +
	( 16'sd 18739) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28087) * $signed(input_fmap_237[7:0]) +
	( 16'sd 26833) * $signed(input_fmap_238[7:0]) +
	( 16'sd 27523) * $signed(input_fmap_239[7:0]) +
	( 15'sd 8531) * $signed(input_fmap_240[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_241[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_242[7:0]) +
	( 16'sd 17687) * $signed(input_fmap_243[7:0]) +
	( 15'sd 14995) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19710) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17014) * $signed(input_fmap_246[7:0]) +
	( 11'sd 889) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21325) * $signed(input_fmap_248[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26948) * $signed(input_fmap_250[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17951) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24897) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26816) * $signed(input_fmap_254[7:0]) +
	( 12'sd 1442) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_186;
assign conv_mac_186 = 
	( 15'sd 12367) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2178) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15217) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30613) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15130) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11901) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8326) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32733) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2328) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10119) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1794) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4523) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2587) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32239) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27051) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6923) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8192) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4478) * $signed(input_fmap_20[7:0]) +
	( 14'sd 7021) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27047) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10795) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2233) * $signed(input_fmap_24[7:0]) +
	( 15'sd 11687) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15300) * $signed(input_fmap_26[7:0]) +
	( 5'sd 13) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31185) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16615) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18307) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25644) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5526) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4782) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12787) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24184) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14305) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31726) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21999) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2824) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29207) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16686) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30047) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7045) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10346) * $signed(input_fmap_47[7:0]) +
	( 15'sd 10067) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23086) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2216) * $signed(input_fmap_50[7:0]) +
	( 16'sd 21920) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25731) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7485) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7807) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3376) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4244) * $signed(input_fmap_56[7:0]) +
	( 16'sd 32190) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28946) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25074) * $signed(input_fmap_59[7:0]) +
	( 15'sd 10088) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6779) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10879) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28923) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2373) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13120) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11058) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23966) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13955) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11446) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29461) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30250) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2840) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10108) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23412) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15744) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16223) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23396) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14388) * $signed(input_fmap_79[7:0]) +
	( 16'sd 22751) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18740) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28527) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11665) * $signed(input_fmap_83[7:0]) +
	( 15'sd 10452) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7578) * $signed(input_fmap_85[7:0]) +
	( 11'sd 955) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3795) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13670) * $signed(input_fmap_89[7:0]) +
	( 10'sd 465) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13266) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12804) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25515) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30855) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11523) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11279) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6258) * $signed(input_fmap_97[7:0]) +
	( 16'sd 31783) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31995) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5587) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28078) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22739) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8983) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7875) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9089) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9117) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28934) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9563) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11540) * $signed(input_fmap_109[7:0]) +
	( 15'sd 14775) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5696) * $signed(input_fmap_111[7:0]) +
	( 15'sd 14303) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31701) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17382) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15135) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6585) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28662) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2251) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3332) * $signed(input_fmap_119[7:0]) +
	( 16'sd 16465) * $signed(input_fmap_120[7:0]) +
	( 14'sd 8030) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21491) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24750) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10156) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20260) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26946) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_127[7:0]) +
	( 14'sd 5247) * $signed(input_fmap_128[7:0]) +
	( 16'sd 29910) * $signed(input_fmap_129[7:0]) +
	( 16'sd 23349) * $signed(input_fmap_130[7:0]) +
	( 16'sd 29630) * $signed(input_fmap_131[7:0]) +
	( 7'sd 51) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10402) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2161) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23008) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1774) * $signed(input_fmap_136[7:0]) +
	( 12'sd 1748) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7260) * $signed(input_fmap_138[7:0]) +
	( 15'sd 12702) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24968) * $signed(input_fmap_140[7:0]) +
	( 16'sd 17514) * $signed(input_fmap_141[7:0]) +
	( 15'sd 15477) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23141) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_144[7:0]) +
	( 16'sd 32755) * $signed(input_fmap_145[7:0]) +
	( 14'sd 4665) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13321) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4472) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27445) * $signed(input_fmap_149[7:0]) +
	( 14'sd 8111) * $signed(input_fmap_150[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16527) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17250) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30630) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22458) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15261) * $signed(input_fmap_157[7:0]) +
	( 16'sd 30582) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20242) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6174) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20566) * $signed(input_fmap_161[7:0]) +
	( 13'sd 4047) * $signed(input_fmap_162[7:0]) +
	( 16'sd 25356) * $signed(input_fmap_163[7:0]) +
	( 16'sd 29202) * $signed(input_fmap_164[7:0]) +
	( 16'sd 20058) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18495) * $signed(input_fmap_166[7:0]) +
	( 16'sd 22399) * $signed(input_fmap_167[7:0]) +
	( 15'sd 8214) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20425) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24705) * $signed(input_fmap_170[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_171[7:0]) +
	( 16'sd 30132) * $signed(input_fmap_172[7:0]) +
	( 16'sd 30204) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32061) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7282) * $signed(input_fmap_175[7:0]) +
	( 15'sd 14904) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15314) * $signed(input_fmap_177[7:0]) +
	( 13'sd 3885) * $signed(input_fmap_178[7:0]) +
	( 16'sd 30430) * $signed(input_fmap_179[7:0]) +
	( 15'sd 13748) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_181[7:0]) +
	( 8'sd 115) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30334) * $signed(input_fmap_183[7:0]) +
	( 11'sd 1015) * $signed(input_fmap_184[7:0]) +
	( 15'sd 9379) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_186[7:0]) +
	( 16'sd 24214) * $signed(input_fmap_187[7:0]) +
	( 14'sd 7249) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5488) * $signed(input_fmap_189[7:0]) +
	( 16'sd 23532) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5813) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19287) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28285) * $signed(input_fmap_193[7:0]) +
	( 16'sd 21869) * $signed(input_fmap_194[7:0]) +
	( 16'sd 18387) * $signed(input_fmap_195[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5851) * $signed(input_fmap_197[7:0]) +
	( 16'sd 17745) * $signed(input_fmap_198[7:0]) +
	( 15'sd 15227) * $signed(input_fmap_199[7:0]) +
	( 11'sd 596) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1535) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14501) * $signed(input_fmap_202[7:0]) +
	( 15'sd 11553) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15691) * $signed(input_fmap_204[7:0]) +
	( 16'sd 21421) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2723) * $signed(input_fmap_206[7:0]) +
	( 15'sd 14901) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14494) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11501) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10523) * $signed(input_fmap_211[7:0]) +
	( 14'sd 4390) * $signed(input_fmap_212[7:0]) +
	( 15'sd 14886) * $signed(input_fmap_213[7:0]) +
	( 16'sd 26291) * $signed(input_fmap_214[7:0]) +
	( 15'sd 12411) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17791) * $signed(input_fmap_216[7:0]) +
	( 14'sd 6462) * $signed(input_fmap_217[7:0]) +
	( 16'sd 18391) * $signed(input_fmap_218[7:0]) +
	( 16'sd 28090) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13594) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1517) * $signed(input_fmap_221[7:0]) +
	( 15'sd 10119) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25023) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1962) * $signed(input_fmap_224[7:0]) +
	( 15'sd 11272) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18125) * $signed(input_fmap_226[7:0]) +
	( 14'sd 4434) * $signed(input_fmap_227[7:0]) +
	( 16'sd 21059) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20994) * $signed(input_fmap_229[7:0]) +
	( 12'sd 1575) * $signed(input_fmap_230[7:0]) +
	( 14'sd 4572) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12892) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28887) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18297) * $signed(input_fmap_234[7:0]) +
	( 16'sd 20910) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_236[7:0]) +
	( 16'sd 32555) * $signed(input_fmap_237[7:0]) +
	( 16'sd 31839) * $signed(input_fmap_238[7:0]) +
	( 16'sd 30077) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25961) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25284) * $signed(input_fmap_241[7:0]) +
	( 11'sd 794) * $signed(input_fmap_242[7:0]) +
	( 16'sd 20534) * $signed(input_fmap_243[7:0]) +
	( 15'sd 15120) * $signed(input_fmap_244[7:0]) +
	( 16'sd 26098) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20361) * $signed(input_fmap_246[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_247[7:0]) +
	( 16'sd 28194) * $signed(input_fmap_248[7:0]) +
	( 15'sd 10589) * $signed(input_fmap_249[7:0]) +
	( 16'sd 23473) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22909) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13027) * $signed(input_fmap_252[7:0]) +
	( 16'sd 20682) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31481) * $signed(input_fmap_254[7:0]) +
	( 13'sd 4016) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_187;
assign conv_mac_187 = 
	( 16'sd 18730) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3062) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8847) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7812) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26137) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22912) * $signed(input_fmap_5[7:0]) +
	( 16'sd 16629) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23806) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12443) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11883) * $signed(input_fmap_9[7:0]) +
	( 16'sd 24104) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6463) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20988) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2870) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30172) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26981) * $signed(input_fmap_17[7:0]) +
	( 15'sd 11778) * $signed(input_fmap_18[7:0]) +
	( 14'sd 8089) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1714) * $signed(input_fmap_20[7:0]) +
	( 16'sd 32609) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29251) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5861) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7378) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3023) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17866) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28741) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31178) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27320) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18018) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27965) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15038) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26762) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12418) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24521) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25596) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26910) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28460) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1054) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29948) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23852) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22180) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6261) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18270) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28259) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14654) * $signed(input_fmap_50[7:0]) +
	( 15'sd 9919) * $signed(input_fmap_51[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14841) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2876) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3465) * $signed(input_fmap_55[7:0]) +
	( 16'sd 27691) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2310) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19495) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1933) * $signed(input_fmap_59[7:0]) +
	( 9'sd 135) * $signed(input_fmap_60[7:0]) +
	( 16'sd 18889) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10441) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22757) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_65[7:0]) +
	( 16'sd 24847) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18747) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5381) * $signed(input_fmap_69[7:0]) +
	( 15'sd 8327) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23063) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11513) * $signed(input_fmap_72[7:0]) +
	( 11'sd 571) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29856) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6403) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9849) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19559) * $signed(input_fmap_77[7:0]) +
	( 11'sd 754) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28297) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2643) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27153) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32757) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12867) * $signed(input_fmap_84[7:0]) +
	( 15'sd 13229) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21232) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30524) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31621) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_89[7:0]) +
	( 10'sd 315) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6514) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21952) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13301) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12719) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23568) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14077) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3921) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10184) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8207) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27425) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30366) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12817) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17474) * $signed(input_fmap_104[7:0]) +
	( 11'sd 987) * $signed(input_fmap_105[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26544) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19933) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7619) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23838) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18966) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19642) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8322) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22266) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12894) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27454) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25736) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2445) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3227) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15274) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3565) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17866) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20838) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22226) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13870) * $signed(input_fmap_125[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21549) * $signed(input_fmap_127[7:0]) +
	( 16'sd 22484) * $signed(input_fmap_128[7:0]) +
	( 15'sd 8306) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1342) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24891) * $signed(input_fmap_131[7:0]) +
	( 16'sd 19957) * $signed(input_fmap_132[7:0]) +
	( 14'sd 5512) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_134[7:0]) +
	( 16'sd 22601) * $signed(input_fmap_135[7:0]) +
	( 15'sd 11249) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_137[7:0]) +
	( 15'sd 14472) * $signed(input_fmap_138[7:0]) +
	( 12'sd 1758) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29974) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5228) * $signed(input_fmap_141[7:0]) +
	( 13'sd 3969) * $signed(input_fmap_142[7:0]) +
	( 16'sd 21197) * $signed(input_fmap_143[7:0]) +
	( 16'sd 17812) * $signed(input_fmap_144[7:0]) +
	( 14'sd 8167) * $signed(input_fmap_145[7:0]) +
	( 15'sd 13126) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27899) * $signed(input_fmap_147[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_148[7:0]) +
	( 16'sd 24157) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15844) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4365) * $signed(input_fmap_151[7:0]) +
	( 16'sd 17107) * $signed(input_fmap_152[7:0]) +
	( 16'sd 19276) * $signed(input_fmap_153[7:0]) +
	( 15'sd 14454) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22873) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24057) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5475) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9319) * $signed(input_fmap_158[7:0]) +
	( 16'sd 23289) * $signed(input_fmap_159[7:0]) +
	( 15'sd 13924) * $signed(input_fmap_160[7:0]) +
	( 15'sd 15690) * $signed(input_fmap_161[7:0]) +
	( 16'sd 27288) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24482) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11971) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14985) * $signed(input_fmap_165[7:0]) +
	( 15'sd 14027) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26494) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27301) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7013) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30593) * $signed(input_fmap_171[7:0]) +
	( 16'sd 23962) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5338) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7196) * $signed(input_fmap_175[7:0]) +
	( 16'sd 17214) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29253) * $signed(input_fmap_177[7:0]) +
	( 10'sd 452) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28676) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26945) * $signed(input_fmap_180[7:0]) +
	( 16'sd 23247) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4317) * $signed(input_fmap_182[7:0]) +
	( 16'sd 27395) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11374) * $signed(input_fmap_184[7:0]) +
	( 16'sd 28637) * $signed(input_fmap_185[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22110) * $signed(input_fmap_187[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_188[7:0]) +
	( 15'sd 8354) * $signed(input_fmap_189[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_190[7:0]) +
	( 15'sd 9152) * $signed(input_fmap_191[7:0]) +
	( 16'sd 30802) * $signed(input_fmap_192[7:0]) +
	( 16'sd 24354) * $signed(input_fmap_193[7:0]) +
	( 10'sd 444) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5401) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19362) * $signed(input_fmap_196[7:0]) +
	( 15'sd 9276) * $signed(input_fmap_197[7:0]) +
	( 12'sd 1231) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20358) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13318) * $signed(input_fmap_200[7:0]) +
	( 16'sd 30620) * $signed(input_fmap_201[7:0]) +
	( 14'sd 4461) * $signed(input_fmap_202[7:0]) +
	( 16'sd 28479) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17194) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24477) * $signed(input_fmap_205[7:0]) +
	( 16'sd 30186) * $signed(input_fmap_206[7:0]) +
	( 16'sd 26506) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30119) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23691) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31245) * $signed(input_fmap_210[7:0]) +
	( 15'sd 9393) * $signed(input_fmap_211[7:0]) +
	( 13'sd 2199) * $signed(input_fmap_212[7:0]) +
	( 16'sd 31551) * $signed(input_fmap_213[7:0]) +
	( 14'sd 4554) * $signed(input_fmap_214[7:0]) +
	( 16'sd 25074) * $signed(input_fmap_215[7:0]) +
	( 16'sd 27281) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19908) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3661) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24023) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1883) * $signed(input_fmap_221[7:0]) +
	( 12'sd 1198) * $signed(input_fmap_222[7:0]) +
	( 15'sd 16379) * $signed(input_fmap_223[7:0]) +
	( 16'sd 28509) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3075) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11707) * $signed(input_fmap_226[7:0]) +
	( 15'sd 10526) * $signed(input_fmap_227[7:0]) +
	( 13'sd 2347) * $signed(input_fmap_228[7:0]) +
	( 16'sd 18608) * $signed(input_fmap_229[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_230[7:0]) +
	( 15'sd 9191) * $signed(input_fmap_231[7:0]) +
	( 15'sd 13957) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24361) * $signed(input_fmap_233[7:0]) +
	( 15'sd 10906) * $signed(input_fmap_234[7:0]) +
	( 16'sd 30570) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5372) * $signed(input_fmap_236[7:0]) +
	( 14'sd 4843) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16759) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5664) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21247) * $signed(input_fmap_241[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_242[7:0]) +
	( 16'sd 17432) * $signed(input_fmap_243[7:0]) +
	( 15'sd 9312) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24170) * $signed(input_fmap_245[7:0]) +
	( 16'sd 27842) * $signed(input_fmap_246[7:0]) +
	( 16'sd 28890) * $signed(input_fmap_247[7:0]) +
	( 16'sd 30579) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4881) * $signed(input_fmap_249[7:0]) +
	( 16'sd 27872) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14290) * $signed(input_fmap_251[7:0]) +
	( 16'sd 19461) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27458) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_254[7:0]) +
	( 16'sd 30909) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_188;
assign conv_mac_188 = 
	( 16'sd 31410) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8876) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23269) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30875) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26577) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11720) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24748) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8441) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4298) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17079) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15885) * $signed(input_fmap_10[7:0]) +
	( 16'sd 18270) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31072) * $signed(input_fmap_12[7:0]) +
	( 15'sd 12778) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8346) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14631) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24553) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22700) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29077) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19159) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11074) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23706) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8362) * $signed(input_fmap_23[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25423) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25573) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14971) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3777) * $signed(input_fmap_28[7:0]) +
	( 10'sd 495) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30338) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26818) * $signed(input_fmap_32[7:0]) +
	( 15'sd 11747) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2887) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15790) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15714) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30421) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13452) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21999) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8371) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21071) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19238) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23855) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13086) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17026) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27260) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19627) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20634) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15000) * $signed(input_fmap_52[7:0]) +
	( 11'sd 539) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23331) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19303) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8778) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28155) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2135) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17753) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27013) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25071) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19335) * $signed(input_fmap_63[7:0]) +
	( 14'sd 7438) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2875) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18878) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11864) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17570) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14753) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28796) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3720) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14434) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30950) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17877) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32431) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30394) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24709) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11382) * $signed(input_fmap_79[7:0]) +
	( 15'sd 10328) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2366) * $signed(input_fmap_81[7:0]) +
	( 9'sd 141) * $signed(input_fmap_82[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31089) * $signed(input_fmap_84[7:0]) +
	( 16'sd 29857) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1599) * $signed(input_fmap_86[7:0]) +
	( 15'sd 12546) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30440) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13974) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20992) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4660) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11502) * $signed(input_fmap_92[7:0]) +
	( 16'sd 23008) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31510) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14767) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11237) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10601) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28389) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2695) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30389) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24277) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5191) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31755) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10795) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22630) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_108[7:0]) +
	( 15'sd 10653) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26920) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6046) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23729) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15593) * $signed(input_fmap_114[7:0]) +
	( 15'sd 16239) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20850) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16657) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15134) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18484) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15793) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28126) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5916) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7677) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27807) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28953) * $signed(input_fmap_125[7:0]) +
	( 14'sd 7565) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4558) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9612) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14574) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19052) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20406) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10897) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22525) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11084) * $signed(input_fmap_134[7:0]) +
	( 13'sd 3715) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2824) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15488) * $signed(input_fmap_137[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_138[7:0]) +
	( 15'sd 16351) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17889) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3819) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22218) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12151) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11023) * $signed(input_fmap_144[7:0]) +
	( 12'sd 1064) * $signed(input_fmap_145[7:0]) +
	( 16'sd 28292) * $signed(input_fmap_146[7:0]) +
	( 16'sd 25740) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28212) * $signed(input_fmap_148[7:0]) +
	( 16'sd 20274) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25042) * $signed(input_fmap_150[7:0]) +
	( 16'sd 21080) * $signed(input_fmap_151[7:0]) +
	( 15'sd 9546) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24773) * $signed(input_fmap_153[7:0]) +
	( 15'sd 14822) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23888) * $signed(input_fmap_155[7:0]) +
	( 13'sd 2877) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5087) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25492) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20398) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31916) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23595) * $signed(input_fmap_161[7:0]) +
	( 16'sd 19874) * $signed(input_fmap_162[7:0]) +
	( 15'sd 14618) * $signed(input_fmap_163[7:0]) +
	( 16'sd 31008) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30032) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9904) * $signed(input_fmap_166[7:0]) +
	( 13'sd 3353) * $signed(input_fmap_167[7:0]) +
	( 16'sd 23957) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2611) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30214) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14538) * $signed(input_fmap_172[7:0]) +
	( 16'sd 26023) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7893) * $signed(input_fmap_174[7:0]) +
	( 14'sd 6666) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18236) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24803) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1291) * $signed(input_fmap_178[7:0]) +
	( 14'sd 7553) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32576) * $signed(input_fmap_180[7:0]) +
	( 14'sd 4992) * $signed(input_fmap_181[7:0]) +
	( 16'sd 24300) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29304) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26849) * $signed(input_fmap_184[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_185[7:0]) +
	( 15'sd 10525) * $signed(input_fmap_186[7:0]) +
	( 16'sd 29586) * $signed(input_fmap_187[7:0]) +
	( 16'sd 20936) * $signed(input_fmap_188[7:0]) +
	( 14'sd 4869) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4284) * $signed(input_fmap_190[7:0]) +
	( 16'sd 27321) * $signed(input_fmap_191[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_192[7:0]) +
	( 16'sd 23221) * $signed(input_fmap_193[7:0]) +
	( 14'sd 7182) * $signed(input_fmap_194[7:0]) +
	( 16'sd 31731) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25692) * $signed(input_fmap_196[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_197[7:0]) +
	( 14'sd 6501) * $signed(input_fmap_198[7:0]) +
	( 15'sd 9682) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_200[7:0]) +
	( 11'sd 688) * $signed(input_fmap_201[7:0]) +
	( 16'sd 22642) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19410) * $signed(input_fmap_203[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_204[7:0]) +
	( 15'sd 16311) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31352) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21853) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12593) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3633) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5924) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6636) * $signed(input_fmap_211[7:0]) +
	( 14'sd 5904) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24647) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23808) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23313) * $signed(input_fmap_215[7:0]) +
	( 16'sd 32197) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9316) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30198) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21221) * $signed(input_fmap_219[7:0]) +
	( 15'sd 12208) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13273) * $signed(input_fmap_221[7:0]) +
	( 15'sd 13393) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24153) * $signed(input_fmap_223[7:0]) +
	( 15'sd 15761) * $signed(input_fmap_224[7:0]) +
	( 11'sd 750) * $signed(input_fmap_225[7:0]) +
	( 15'sd 9553) * $signed(input_fmap_226[7:0]) +
	( 15'sd 16181) * $signed(input_fmap_227[7:0]) +
	( 16'sd 23458) * $signed(input_fmap_228[7:0]) +
	( 16'sd 25738) * $signed(input_fmap_229[7:0]) +
	( 14'sd 7519) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_231[7:0]) +
	( 16'sd 16733) * $signed(input_fmap_232[7:0]) +
	( 16'sd 25672) * $signed(input_fmap_233[7:0]) +
	( 15'sd 8215) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29993) * $signed(input_fmap_235[7:0]) +
	( 16'sd 20687) * $signed(input_fmap_236[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17047) * $signed(input_fmap_238[7:0]) +
	( 16'sd 24056) * $signed(input_fmap_239[7:0]) +
	( 16'sd 17471) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15749) * $signed(input_fmap_242[7:0]) +
	( 16'sd 30185) * $signed(input_fmap_243[7:0]) +
	( 15'sd 14974) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10291) * $signed(input_fmap_245[7:0]) +
	( 16'sd 18019) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8659) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18178) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3516) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12011) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28282) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29125) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31153) * $signed(input_fmap_254[7:0]) +
	( 15'sd 13195) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_189;
assign conv_mac_189 = 
	( 15'sd 13163) * $signed(input_fmap_0[7:0]) +
	( 13'sd 2143) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5437) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14499) * $signed(input_fmap_3[7:0]) +
	( 16'sd 18870) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27464) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28256) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29145) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7624) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23803) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20978) * $signed(input_fmap_10[7:0]) +
	( 16'sd 32060) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12799) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13347) * $signed(input_fmap_13[7:0]) +
	( 15'sd 16258) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14358) * $signed(input_fmap_15[7:0]) +
	( 11'sd 784) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1949) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4348) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10990) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27688) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20964) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13037) * $signed(input_fmap_22[7:0]) +
	( 16'sd 31359) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11336) * $signed(input_fmap_24[7:0]) +
	( 16'sd 29759) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11416) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18243) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28310) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28689) * $signed(input_fmap_29[7:0]) +
	( 16'sd 24654) * $signed(input_fmap_30[7:0]) +
	( 15'sd 9709) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15602) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32643) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27702) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19451) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2594) * $signed(input_fmap_36[7:0]) +
	( 8'sd 75) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6335) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12802) * $signed(input_fmap_39[7:0]) +
	( 10'sd 477) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24228) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29790) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16089) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21026) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2630) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9118) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26794) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6338) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7890) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20056) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13127) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19562) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10706) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4713) * $signed(input_fmap_54[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3696) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14170) * $signed(input_fmap_57[7:0]) +
	( 16'sd 25432) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18837) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19444) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11115) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25196) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10175) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19621) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29583) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21196) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7401) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30481) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5859) * $signed(input_fmap_69[7:0]) +
	( 16'sd 28245) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21964) * $signed(input_fmap_71[7:0]) +
	( 16'sd 22856) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26420) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23264) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20385) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9808) * $signed(input_fmap_77[7:0]) +
	( 15'sd 8269) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7730) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23005) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11825) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4440) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21205) * $signed(input_fmap_83[7:0]) +
	( 16'sd 29926) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19319) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8639) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17229) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23436) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13335) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10910) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13892) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9923) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1592) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29947) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2061) * $signed(input_fmap_99[7:0]) +
	( 15'sd 9263) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15423) * $signed(input_fmap_101[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28943) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9761) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14142) * $signed(input_fmap_105[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13613) * $signed(input_fmap_107[7:0]) +
	( 15'sd 15064) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22059) * $signed(input_fmap_109[7:0]) +
	( 15'sd 16296) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19077) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2535) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32062) * $signed(input_fmap_113[7:0]) +
	( 12'sd 1703) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30823) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12290) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29399) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26429) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24068) * $signed(input_fmap_119[7:0]) +
	( 16'sd 24624) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25977) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1833) * $signed(input_fmap_122[7:0]) +
	( 12'sd 1653) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23222) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1150) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13867) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25567) * $signed(input_fmap_127[7:0]) +
	( 16'sd 22670) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5657) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14496) * $signed(input_fmap_130[7:0]) +
	( 16'sd 30443) * $signed(input_fmap_131[7:0]) +
	( 16'sd 21354) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28850) * $signed(input_fmap_133[7:0]) +
	( 14'sd 7486) * $signed(input_fmap_134[7:0]) +
	( 15'sd 13639) * $signed(input_fmap_135[7:0]) +
	( 14'sd 5447) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6709) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7427) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18148) * $signed(input_fmap_139[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_140[7:0]) +
	( 14'sd 4146) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30790) * $signed(input_fmap_142[7:0]) +
	( 16'sd 19063) * $signed(input_fmap_143[7:0]) +
	( 16'sd 30867) * $signed(input_fmap_144[7:0]) +
	( 14'sd 4607) * $signed(input_fmap_145[7:0]) +
	( 16'sd 17922) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9615) * $signed(input_fmap_147[7:0]) +
	( 15'sd 9644) * $signed(input_fmap_148[7:0]) +
	( 14'sd 6946) * $signed(input_fmap_149[7:0]) +
	( 9'sd 248) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4222) * $signed(input_fmap_151[7:0]) +
	( 16'sd 26241) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25051) * $signed(input_fmap_153[7:0]) +
	( 16'sd 32422) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10227) * $signed(input_fmap_155[7:0]) +
	( 16'sd 22568) * $signed(input_fmap_156[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18230) * $signed(input_fmap_158[7:0]) +
	( 15'sd 11508) * $signed(input_fmap_159[7:0]) +
	( 16'sd 20844) * $signed(input_fmap_160[7:0]) +
	( 13'sd 2360) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2124) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27046) * $signed(input_fmap_163[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_164[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_165[7:0]) +
	( 16'sd 32415) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26102) * $signed(input_fmap_167[7:0]) +
	( 16'sd 23539) * $signed(input_fmap_168[7:0]) +
	( 16'sd 23108) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23078) * $signed(input_fmap_170[7:0]) +
	( 13'sd 2415) * $signed(input_fmap_171[7:0]) +
	( 16'sd 26374) * $signed(input_fmap_172[7:0]) +
	( 15'sd 8740) * $signed(input_fmap_173[7:0]) +
	( 15'sd 16045) * $signed(input_fmap_174[7:0]) +
	( 16'sd 16520) * $signed(input_fmap_175[7:0]) +
	( 8'sd 79) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_177[7:0]) +
	( 16'sd 28838) * $signed(input_fmap_178[7:0]) +
	( 16'sd 19307) * $signed(input_fmap_179[7:0]) +
	( 15'sd 11152) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6004) * $signed(input_fmap_181[7:0]) +
	( 16'sd 29714) * $signed(input_fmap_182[7:0]) +
	( 16'sd 18063) * $signed(input_fmap_183[7:0]) +
	( 13'sd 2772) * $signed(input_fmap_184[7:0]) +
	( 16'sd 19552) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9247) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28018) * $signed(input_fmap_187[7:0]) +
	( 15'sd 9372) * $signed(input_fmap_188[7:0]) +
	( 15'sd 15758) * $signed(input_fmap_189[7:0]) +
	( 14'sd 8002) * $signed(input_fmap_190[7:0]) +
	( 15'sd 16295) * $signed(input_fmap_191[7:0]) +
	( 16'sd 23708) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11026) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3560) * $signed(input_fmap_194[7:0]) +
	( 14'sd 7098) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20395) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24780) * $signed(input_fmap_197[7:0]) +
	( 11'sd 583) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16136) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18376) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15766) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21736) * $signed(input_fmap_202[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19445) * $signed(input_fmap_204[7:0]) +
	( 16'sd 27550) * $signed(input_fmap_205[7:0]) +
	( 15'sd 16245) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13285) * $signed(input_fmap_207[7:0]) +
	( 15'sd 10411) * $signed(input_fmap_208[7:0]) +
	( 16'sd 19739) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5150) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23894) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24376) * $signed(input_fmap_212[7:0]) +
	( 16'sd 18732) * $signed(input_fmap_213[7:0]) +
	( 16'sd 16587) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17066) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20467) * $signed(input_fmap_216[7:0]) +
	( 14'sd 7574) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30893) * $signed(input_fmap_218[7:0]) +
	( 16'sd 23433) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4107) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6758) * $signed(input_fmap_221[7:0]) +
	( 13'sd 2626) * $signed(input_fmap_222[7:0]) +
	( 16'sd 18864) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17582) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5254) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30495) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10685) * $signed(input_fmap_228[7:0]) +
	( 15'sd 11010) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14018) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10316) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_232[7:0]) +
	( 15'sd 11585) * $signed(input_fmap_233[7:0]) +
	( 12'sd 1107) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19901) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11884) * $signed(input_fmap_236[7:0]) +
	( 14'sd 6241) * $signed(input_fmap_237[7:0]) +
	( 13'sd 2068) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20355) * $signed(input_fmap_239[7:0]) +
	( 16'sd 27555) * $signed(input_fmap_240[7:0]) +
	( 16'sd 27669) * $signed(input_fmap_241[7:0]) +
	( 16'sd 19186) * $signed(input_fmap_242[7:0]) +
	( 13'sd 3399) * $signed(input_fmap_243[7:0]) +
	( 16'sd 16607) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2540) * $signed(input_fmap_245[7:0]) +
	( 11'sd 548) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9663) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18451) * $signed(input_fmap_248[7:0]) +
	( 12'sd 1158) * $signed(input_fmap_249[7:0]) +
	( 16'sd 18102) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14882) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17962) * $signed(input_fmap_252[7:0]) +
	( 16'sd 30936) * $signed(input_fmap_253[7:0]) +
	( 16'sd 17199) * $signed(input_fmap_254[7:0]) +
	( 16'sd 30318) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_190;
assign conv_mac_190 = 
	( 16'sd 26157) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14368) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11669) * $signed(input_fmap_2[7:0]) +
	( 10'sd 312) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13983) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4459) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25545) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29177) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28850) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21446) * $signed(input_fmap_9[7:0]) +
	( 16'sd 18957) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3856) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6130) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14730) * $signed(input_fmap_14[7:0]) +
	( 16'sd 23818) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12222) * $signed(input_fmap_16[7:0]) +
	( 15'sd 8522) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28088) * $signed(input_fmap_18[7:0]) +
	( 15'sd 16030) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5313) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_21[7:0]) +
	( 15'sd 15995) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15766) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26048) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14340) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27747) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11918) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31721) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31955) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29007) * $signed(input_fmap_32[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19863) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24556) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15147) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28611) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6830) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30030) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5534) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10806) * $signed(input_fmap_41[7:0]) +
	( 13'sd 2991) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13503) * $signed(input_fmap_43[7:0]) +
	( 16'sd 27358) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27948) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14130) * $signed(input_fmap_46[7:0]) +
	( 15'sd 8747) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1104) * $signed(input_fmap_48[7:0]) +
	( 15'sd 14135) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19761) * $signed(input_fmap_50[7:0]) +
	( 15'sd 10037) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28245) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24588) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13621) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9094) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10066) * $signed(input_fmap_56[7:0]) +
	( 8'sd 111) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_58[7:0]) +
	( 13'sd 3692) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32560) * $signed(input_fmap_60[7:0]) +
	( 16'sd 22432) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10769) * $signed(input_fmap_62[7:0]) +
	( 15'sd 8587) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6879) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19008) * $signed(input_fmap_65[7:0]) +
	( 11'sd 592) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30941) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27270) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1846) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20812) * $signed(input_fmap_70[7:0]) +
	( 15'sd 10186) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5763) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18827) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29072) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3049) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11236) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29886) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24768) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3297) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1286) * $signed(input_fmap_80[7:0]) +
	( 15'sd 8627) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20622) * $signed(input_fmap_82[7:0]) +
	( 11'sd 936) * $signed(input_fmap_83[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6470) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14051) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24747) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27785) * $signed(input_fmap_88[7:0]) +
	( 14'sd 4625) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16844) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22403) * $signed(input_fmap_91[7:0]) +
	( 13'sd 2542) * $signed(input_fmap_92[7:0]) +
	( 14'sd 7616) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18146) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30320) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5880) * $signed(input_fmap_96[7:0]) +
	( 15'sd 9708) * $signed(input_fmap_97[7:0]) +
	( 14'sd 5376) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32036) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28323) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26356) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14424) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12480) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24661) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2192) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10139) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4626) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20164) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24118) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13365) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14292) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11552) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12738) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13204) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20308) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_116[7:0]) +
	( 16'sd 30376) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20270) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18331) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18117) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1264) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1493) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11619) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24882) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5925) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11275) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29388) * $signed(input_fmap_127[7:0]) +
	( 16'sd 20309) * $signed(input_fmap_128[7:0]) +
	( 15'sd 15668) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10867) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14811) * $signed(input_fmap_132[7:0]) +
	( 11'sd 918) * $signed(input_fmap_133[7:0]) +
	( 16'sd 27790) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19075) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21233) * $signed(input_fmap_136[7:0]) +
	( 15'sd 14825) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32549) * $signed(input_fmap_138[7:0]) +
	( 11'sd 727) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_140[7:0]) +
	( 16'sd 28064) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11484) * $signed(input_fmap_142[7:0]) +
	( 11'sd 531) * $signed(input_fmap_143[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21753) * $signed(input_fmap_145[7:0]) +
	( 16'sd 22320) * $signed(input_fmap_146[7:0]) +
	( 16'sd 20288) * $signed(input_fmap_147[7:0]) +
	( 14'sd 5540) * $signed(input_fmap_148[7:0]) +
	( 16'sd 19396) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25126) * $signed(input_fmap_150[7:0]) +
	( 16'sd 31622) * $signed(input_fmap_151[7:0]) +
	( 14'sd 5503) * $signed(input_fmap_152[7:0]) +
	( 16'sd 22498) * $signed(input_fmap_153[7:0]) +
	( 15'sd 13118) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30777) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22042) * $signed(input_fmap_157[7:0]) +
	( 16'sd 28586) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6010) * $signed(input_fmap_159[7:0]) +
	( 16'sd 16406) * $signed(input_fmap_160[7:0]) +
	( 15'sd 9579) * $signed(input_fmap_161[7:0]) +
	( 14'sd 8083) * $signed(input_fmap_162[7:0]) +
	( 16'sd 29398) * $signed(input_fmap_163[7:0]) +
	( 16'sd 20123) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28697) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4796) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_167[7:0]) +
	( 16'sd 19542) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26319) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_170[7:0]) +
	( 13'sd 4076) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14716) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23228) * $signed(input_fmap_173[7:0]) +
	( 16'sd 23412) * $signed(input_fmap_174[7:0]) +
	( 16'sd 27618) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15973) * $signed(input_fmap_176[7:0]) +
	( 15'sd 11593) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32304) * $signed(input_fmap_178[7:0]) +
	( 15'sd 14505) * $signed(input_fmap_179[7:0]) +
	( 14'sd 4307) * $signed(input_fmap_180[7:0]) +
	( 13'sd 2305) * $signed(input_fmap_181[7:0]) +
	( 16'sd 28013) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12476) * $signed(input_fmap_183[7:0]) +
	( 16'sd 16598) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17694) * $signed(input_fmap_185[7:0]) +
	( 15'sd 8195) * $signed(input_fmap_186[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_187[7:0]) +
	( 16'sd 25197) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5106) * $signed(input_fmap_189[7:0]) +
	( 13'sd 3765) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14437) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31930) * $signed(input_fmap_192[7:0]) +
	( 12'sd 1067) * $signed(input_fmap_193[7:0]) +
	( 16'sd 24018) * $signed(input_fmap_194[7:0]) +
	( 16'sd 20159) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22358) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21136) * $signed(input_fmap_197[7:0]) +
	( 16'sd 21421) * $signed(input_fmap_198[7:0]) +
	( 15'sd 11963) * $signed(input_fmap_199[7:0]) +
	( 11'sd 524) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3642) * $signed(input_fmap_201[7:0]) +
	( 14'sd 4355) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17113) * $signed(input_fmap_204[7:0]) +
	( 16'sd 21762) * $signed(input_fmap_205[7:0]) +
	( 16'sd 24806) * $signed(input_fmap_206[7:0]) +
	( 15'sd 14661) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18959) * $signed(input_fmap_208[7:0]) +
	( 13'sd 2959) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18771) * $signed(input_fmap_210[7:0]) +
	( 16'sd 29343) * $signed(input_fmap_211[7:0]) +
	( 16'sd 28807) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28596) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28944) * $signed(input_fmap_214[7:0]) +
	( 16'sd 27332) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5878) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32321) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10862) * $signed(input_fmap_218[7:0]) +
	( 16'sd 16692) * $signed(input_fmap_219[7:0]) +
	( 15'sd 11717) * $signed(input_fmap_220[7:0]) +
	( 16'sd 20406) * $signed(input_fmap_221[7:0]) +
	( 11'sd 629) * $signed(input_fmap_222[7:0]) +
	( 15'sd 16077) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6640) * $signed(input_fmap_224[7:0]) +
	( 16'sd 19618) * $signed(input_fmap_225[7:0]) +
	( 16'sd 17239) * $signed(input_fmap_226[7:0]) +
	( 15'sd 8265) * $signed(input_fmap_227[7:0]) +
	( 15'sd 16338) * $signed(input_fmap_228[7:0]) +
	( 14'sd 4357) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30027) * $signed(input_fmap_230[7:0]) +
	( 8'sd 114) * $signed(input_fmap_231[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27748) * $signed(input_fmap_233[7:0]) +
	( 16'sd 30335) * $signed(input_fmap_234[7:0]) +
	( 14'sd 4814) * $signed(input_fmap_235[7:0]) +
	( 16'sd 22352) * $signed(input_fmap_236[7:0]) +
	( 16'sd 18982) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19729) * $signed(input_fmap_238[7:0]) +
	( 16'sd 29581) * $signed(input_fmap_239[7:0]) +
	( 16'sd 21747) * $signed(input_fmap_240[7:0]) +
	( 16'sd 22151) * $signed(input_fmap_241[7:0]) +
	( 16'sd 20546) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28319) * $signed(input_fmap_243[7:0]) +
	( 15'sd 14803) * $signed(input_fmap_244[7:0]) +
	( 16'sd 29393) * $signed(input_fmap_245[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17683) * $signed(input_fmap_247[7:0]) +
	( 16'sd 27810) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28262) * $signed(input_fmap_249[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_250[7:0]) +
	( 15'sd 11793) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13262) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17549) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23866) * $signed(input_fmap_254[7:0]) +
	( 14'sd 4907) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_191;
assign conv_mac_191 = 
	( 16'sd 31185) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32522) * $signed(input_fmap_1[7:0]) +
	( 11'sd 907) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19431) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32327) * $signed(input_fmap_4[7:0]) +
	( 13'sd 4066) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22020) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31560) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3331) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22392) * $signed(input_fmap_9[7:0]) +
	( 11'sd 951) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19080) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28736) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3529) * $signed(input_fmap_13[7:0]) +
	( 15'sd 13123) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2487) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27489) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26430) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14031) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23045) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20337) * $signed(input_fmap_21[7:0]) +
	( 13'sd 3342) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21218) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9239) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5024) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7073) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4296) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5639) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19889) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32093) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4854) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8638) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10187) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21410) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17449) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7665) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14285) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6041) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13250) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5952) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30453) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14603) * $signed(input_fmap_43[7:0]) +
	( 10'sd 505) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18965) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22545) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6938) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3244) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28541) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32120) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22642) * $signed(input_fmap_51[7:0]) +
	( 16'sd 17070) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1521) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6997) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10158) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23113) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4151) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28629) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27177) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25548) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16122) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5463) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3091) * $signed(input_fmap_64[7:0]) +
	( 15'sd 11341) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22462) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23136) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14914) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24296) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11895) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28355) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_73[7:0]) +
	( 16'sd 30965) * $signed(input_fmap_74[7:0]) +
	( 16'sd 21854) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27617) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31242) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30521) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31742) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17021) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18168) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7465) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14416) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6869) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9472) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3720) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27094) * $signed(input_fmap_88[7:0]) +
	( 15'sd 8900) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10838) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12897) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21871) * $signed(input_fmap_93[7:0]) +
	( 16'sd 24385) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26880) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10311) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25818) * $signed(input_fmap_97[7:0]) +
	( 16'sd 18734) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9316) * $signed(input_fmap_99[7:0]) +
	( 12'sd 1183) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27532) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28196) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20430) * $signed(input_fmap_103[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11957) * $signed(input_fmap_105[7:0]) +
	( 15'sd 12521) * $signed(input_fmap_106[7:0]) +
	( 15'sd 15911) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20978) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22586) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20982) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15348) * $signed(input_fmap_112[7:0]) +
	( 11'sd 553) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26990) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31380) * $signed(input_fmap_115[7:0]) +
	( 14'sd 8023) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23708) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20325) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18318) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30034) * $signed(input_fmap_121[7:0]) +
	( 15'sd 8529) * $signed(input_fmap_122[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11517) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32585) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30259) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12776) * $signed(input_fmap_127[7:0]) +
	( 15'sd 10201) * $signed(input_fmap_128[7:0]) +
	( 16'sd 20577) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15407) * $signed(input_fmap_131[7:0]) +
	( 16'sd 23151) * $signed(input_fmap_132[7:0]) +
	( 16'sd 32687) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2211) * $signed(input_fmap_134[7:0]) +
	( 14'sd 7172) * $signed(input_fmap_135[7:0]) +
	( 16'sd 20954) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9853) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9199) * $signed(input_fmap_138[7:0]) +
	( 14'sd 5824) * $signed(input_fmap_139[7:0]) +
	( 14'sd 6989) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24178) * $signed(input_fmap_141[7:0]) +
	( 16'sd 20061) * $signed(input_fmap_142[7:0]) +
	( 11'sd 761) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2229) * $signed(input_fmap_144[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_145[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17896) * $signed(input_fmap_148[7:0]) +
	( 15'sd 10141) * $signed(input_fmap_149[7:0]) +
	( 16'sd 25977) * $signed(input_fmap_150[7:0]) +
	( 14'sd 6926) * $signed(input_fmap_151[7:0]) +
	( 16'sd 18673) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11906) * $signed(input_fmap_153[7:0]) +
	( 16'sd 32588) * $signed(input_fmap_154[7:0]) +
	( 16'sd 24074) * $signed(input_fmap_155[7:0]) +
	( 14'sd 5722) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11010) * $signed(input_fmap_157[7:0]) +
	( 16'sd 18131) * $signed(input_fmap_158[7:0]) +
	( 16'sd 22416) * $signed(input_fmap_159[7:0]) +
	( 15'sd 16369) * $signed(input_fmap_160[7:0]) +
	( 10'sd 430) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10239) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8798) * $signed(input_fmap_163[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_164[7:0]) +
	( 16'sd 32298) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22952) * $signed(input_fmap_166[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5343) * $signed(input_fmap_168[7:0]) +
	( 11'sd 921) * $signed(input_fmap_169[7:0]) +
	( 16'sd 29182) * $signed(input_fmap_170[7:0]) +
	( 13'sd 3169) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31326) * $signed(input_fmap_172[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_173[7:0]) +
	( 16'sd 19312) * $signed(input_fmap_174[7:0]) +
	( 16'sd 18349) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20627) * $signed(input_fmap_176[7:0]) +
	( 15'sd 11209) * $signed(input_fmap_177[7:0]) +
	( 14'sd 7961) * $signed(input_fmap_178[7:0]) +
	( 16'sd 24369) * $signed(input_fmap_179[7:0]) +
	( 16'sd 19125) * $signed(input_fmap_180[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30623) * $signed(input_fmap_182[7:0]) +
	( 15'sd 13073) * $signed(input_fmap_183[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_185[7:0]) +
	( 16'sd 28912) * $signed(input_fmap_186[7:0]) +
	( 13'sd 4035) * $signed(input_fmap_187[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30235) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20296) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23686) * $signed(input_fmap_191[7:0]) +
	( 14'sd 5972) * $signed(input_fmap_192[7:0]) +
	( 16'sd 32168) * $signed(input_fmap_193[7:0]) +
	( 16'sd 24099) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5461) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20275) * $signed(input_fmap_196[7:0]) +
	( 13'sd 2950) * $signed(input_fmap_197[7:0]) +
	( 15'sd 11182) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20909) * $signed(input_fmap_200[7:0]) +
	( 16'sd 21459) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5556) * $signed(input_fmap_202[7:0]) +
	( 15'sd 9126) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_204[7:0]) +
	( 15'sd 9835) * $signed(input_fmap_205[7:0]) +
	( 16'sd 30217) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29204) * $signed(input_fmap_207[7:0]) +
	( 16'sd 16803) * $signed(input_fmap_208[7:0]) +
	( 14'sd 4142) * $signed(input_fmap_209[7:0]) +
	( 16'sd 28772) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30877) * $signed(input_fmap_211[7:0]) +
	( 16'sd 30902) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1597) * $signed(input_fmap_213[7:0]) +
	( 14'sd 6009) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17538) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18548) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17659) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21943) * $signed(input_fmap_218[7:0]) +
	( 16'sd 22481) * $signed(input_fmap_219[7:0]) +
	( 16'sd 29211) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5118) * $signed(input_fmap_221[7:0]) +
	( 15'sd 16006) * $signed(input_fmap_222[7:0]) +
	( 16'sd 27225) * $signed(input_fmap_223[7:0]) +
	( 16'sd 26378) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13226) * $signed(input_fmap_225[7:0]) +
	( 16'sd 28263) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2575) * $signed(input_fmap_227[7:0]) +
	( 16'sd 32048) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6830) * $signed(input_fmap_229[7:0]) +
	( 16'sd 26512) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1590) * $signed(input_fmap_231[7:0]) +
	( 15'sd 15643) * $signed(input_fmap_232[7:0]) +
	( 16'sd 19626) * $signed(input_fmap_233[7:0]) +
	( 13'sd 2151) * $signed(input_fmap_234[7:0]) +
	( 6'sd 17) * $signed(input_fmap_235[7:0]) +
	( 15'sd 13100) * $signed(input_fmap_236[7:0]) +
	( 14'sd 5758) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14435) * $signed(input_fmap_238[7:0]) +
	( 12'sd 1863) * $signed(input_fmap_239[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_240[7:0]) +
	( 15'sd 16154) * $signed(input_fmap_241[7:0]) +
	( 16'sd 30235) * $signed(input_fmap_242[7:0]) +
	( 16'sd 26254) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19926) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3015) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23607) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15467) * $signed(input_fmap_247[7:0]) +
	( 16'sd 20712) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12778) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_251[7:0]) +
	( 16'sd 29373) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_253[7:0]) +
	( 14'sd 5004) * $signed(input_fmap_254[7:0]) +
	( 14'sd 8077) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_192;
assign conv_mac_192 = 
	( 15'sd 8735) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16140) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13347) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10494) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27590) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2589) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9061) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19989) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26630) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10125) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26454) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17110) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17119) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15589) * $signed(input_fmap_15[7:0]) +
	( 13'sd 4009) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16665) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14674) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20162) * $signed(input_fmap_19[7:0]) +
	( 15'sd 10934) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20920) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24458) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19550) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12287) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15243) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17956) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6889) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13175) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24384) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15799) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24051) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15203) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32665) * $signed(input_fmap_33[7:0]) +
	( 16'sd 20114) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12517) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32133) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13092) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8666) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13891) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10853) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27049) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19577) * $signed(input_fmap_42[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7963) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16170) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26252) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25937) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26299) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29141) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18031) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11344) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29842) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21063) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25660) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15036) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24535) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12571) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31391) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11005) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25590) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26769) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9205) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19298) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6545) * $signed(input_fmap_65[7:0]) +
	( 10'sd 358) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5805) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19472) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24695) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24451) * $signed(input_fmap_71[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_72[7:0]) +
	( 16'sd 18921) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9168) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13244) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4931) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18701) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22852) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29916) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28557) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28947) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31929) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7831) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28960) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26235) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31832) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13328) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10596) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6403) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12348) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13378) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25141) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24160) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6878) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32531) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11132) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27532) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31267) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1072) * $signed(input_fmap_101[7:0]) +
	( 9'sd 176) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17095) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25218) * $signed(input_fmap_104[7:0]) +
	( 16'sd 18461) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27265) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10312) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5511) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4411) * $signed(input_fmap_109[7:0]) +
	( 14'sd 6527) * $signed(input_fmap_110[7:0]) +
	( 16'sd 31048) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11839) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26399) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30443) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5889) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14307) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17935) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16783) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17088) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11081) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28360) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23035) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2781) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3437) * $signed(input_fmap_124[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13284) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28573) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2196) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14823) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19595) * $signed(input_fmap_130[7:0]) +
	( 15'sd 11421) * $signed(input_fmap_131[7:0]) +
	( 15'sd 13859) * $signed(input_fmap_132[7:0]) +
	( 15'sd 11587) * $signed(input_fmap_133[7:0]) +
	( 16'sd 30916) * $signed(input_fmap_134[7:0]) +
	( 16'sd 24604) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13987) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26219) * $signed(input_fmap_137[7:0]) +
	( 16'sd 26074) * $signed(input_fmap_138[7:0]) +
	( 15'sd 9643) * $signed(input_fmap_139[7:0]) +
	( 16'sd 31049) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19189) * $signed(input_fmap_141[7:0]) +
	( 16'sd 16676) * $signed(input_fmap_142[7:0]) +
	( 16'sd 29882) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3844) * $signed(input_fmap_144[7:0]) +
	( 14'sd 7240) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7012) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17026) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23205) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25296) * $signed(input_fmap_149[7:0]) +
	( 16'sd 29105) * $signed(input_fmap_150[7:0]) +
	( 16'sd 21057) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20401) * $signed(input_fmap_152[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4615) * $signed(input_fmap_154[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_155[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20836) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25771) * $signed(input_fmap_158[7:0]) +
	( 15'sd 16342) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27017) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22965) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2377) * $signed(input_fmap_162[7:0]) +
	( 16'sd 21672) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11813) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2622) * $signed(input_fmap_165[7:0]) +
	( 15'sd 15994) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26435) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20735) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14407) * $signed(input_fmap_170[7:0]) +
	( 16'sd 20291) * $signed(input_fmap_171[7:0]) +
	( 10'sd 430) * $signed(input_fmap_172[7:0]) +
	( 16'sd 16849) * $signed(input_fmap_173[7:0]) +
	( 16'sd 28526) * $signed(input_fmap_174[7:0]) +
	( 16'sd 30060) * $signed(input_fmap_175[7:0]) +
	( 16'sd 28196) * $signed(input_fmap_176[7:0]) +
	( 16'sd 17510) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22222) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28646) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24670) * $signed(input_fmap_180[7:0]) +
	( 16'sd 22228) * $signed(input_fmap_181[7:0]) +
	( 15'sd 13901) * $signed(input_fmap_182[7:0]) +
	( 16'sd 19265) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26287) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24341) * $signed(input_fmap_185[7:0]) +
	( 11'sd 629) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9964) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17781) * $signed(input_fmap_188[7:0]) +
	( 16'sd 24455) * $signed(input_fmap_189[7:0]) +
	( 14'sd 8048) * $signed(input_fmap_190[7:0]) +
	( 16'sd 18333) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19101) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26778) * $signed(input_fmap_193[7:0]) +
	( 16'sd 19653) * $signed(input_fmap_194[7:0]) +
	( 16'sd 30425) * $signed(input_fmap_195[7:0]) +
	( 16'sd 23251) * $signed(input_fmap_196[7:0]) +
	( 16'sd 16740) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29667) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10285) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26095) * $signed(input_fmap_200[7:0]) +
	( 14'sd 4634) * $signed(input_fmap_201[7:0]) +
	( 13'sd 4090) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_203[7:0]) +
	( 13'sd 3158) * $signed(input_fmap_204[7:0]) +
	( 16'sd 25041) * $signed(input_fmap_205[7:0]) +
	( 16'sd 19435) * $signed(input_fmap_206[7:0]) +
	( 15'sd 15188) * $signed(input_fmap_207[7:0]) +
	( 16'sd 20484) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18982) * $signed(input_fmap_209[7:0]) +
	( 15'sd 13233) * $signed(input_fmap_210[7:0]) +
	( 15'sd 14489) * $signed(input_fmap_211[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_212[7:0]) +
	( 16'sd 19905) * $signed(input_fmap_213[7:0]) +
	( 16'sd 26883) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22426) * $signed(input_fmap_215[7:0]) +
	( 16'sd 26353) * $signed(input_fmap_216[7:0]) +
	( 15'sd 15435) * $signed(input_fmap_217[7:0]) +
	( 16'sd 32072) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15564) * $signed(input_fmap_219[7:0]) +
	( 16'sd 23230) * $signed(input_fmap_220[7:0]) +
	( 14'sd 7986) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3661) * $signed(input_fmap_222[7:0]) +
	( 16'sd 18731) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12316) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1109) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10311) * $signed(input_fmap_226[7:0]) +
	( 16'sd 30681) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18563) * $signed(input_fmap_228[7:0]) +
	( 16'sd 19748) * $signed(input_fmap_229[7:0]) +
	( 13'sd 2598) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17228) * $signed(input_fmap_231[7:0]) +
	( 15'sd 16144) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18477) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4680) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_235[7:0]) +
	( 15'sd 16236) * $signed(input_fmap_236[7:0]) +
	( 13'sd 4046) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22446) * $signed(input_fmap_238[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25983) * $signed(input_fmap_240[7:0]) +
	( 15'sd 16114) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27358) * $signed(input_fmap_242[7:0]) +
	( 15'sd 14409) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24382) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23322) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12951) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21882) * $signed(input_fmap_248[7:0]) +
	( 16'sd 27939) * $signed(input_fmap_249[7:0]) +
	( 16'sd 31873) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21857) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10760) * $signed(input_fmap_252[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_253[7:0]) +
	( 15'sd 8622) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20470) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_193;
assign conv_mac_193 = 
	( 16'sd 17879) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8716) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27122) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12217) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29486) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30770) * $signed(input_fmap_6[7:0]) +
	( 16'sd 27242) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22427) * $signed(input_fmap_8[7:0]) +
	( 7'sd 57) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23360) * $signed(input_fmap_10[7:0]) +
	( 15'sd 16257) * $signed(input_fmap_11[7:0]) +
	( 16'sd 19008) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13089) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19668) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6563) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16152) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7232) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25627) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11422) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23449) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21610) * $signed(input_fmap_21[7:0]) +
	( 7'sd 40) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10399) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11499) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20642) * $signed(input_fmap_25[7:0]) +
	( 15'sd 12340) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20534) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9912) * $signed(input_fmap_28[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10517) * $signed(input_fmap_30[7:0]) +
	( 16'sd 23185) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5884) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2815) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23793) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31533) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30259) * $signed(input_fmap_36[7:0]) +
	( 16'sd 27790) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27715) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19737) * $signed(input_fmap_39[7:0]) +
	( 11'sd 599) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_41[7:0]) +
	( 16'sd 17421) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14432) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19851) * $signed(input_fmap_44[7:0]) +
	( 9'sd 197) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4750) * $signed(input_fmap_46[7:0]) +
	( 16'sd 30312) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7969) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20048) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1832) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19498) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2135) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1427) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_54[7:0]) +
	( 9'sd 253) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23364) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5840) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_58[7:0]) +
	( 15'sd 13425) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18345) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9389) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9802) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19362) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1577) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30785) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11349) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6343) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11787) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12833) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_71[7:0]) +
	( 16'sd 21255) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29137) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31734) * $signed(input_fmap_74[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11592) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22331) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23191) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7496) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29984) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16820) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5917) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2800) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2897) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8280) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7934) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24078) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32255) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32269) * $signed(input_fmap_90[7:0]) +
	( 16'sd 23342) * $signed(input_fmap_91[7:0]) +
	( 15'sd 13225) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25331) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11919) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4842) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13239) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5478) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21386) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11197) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27778) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4695) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2240) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31372) * $signed(input_fmap_103[7:0]) +
	( 16'sd 26535) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12277) * $signed(input_fmap_105[7:0]) +
	( 10'sd 272) * $signed(input_fmap_106[7:0]) +
	( 12'sd 1565) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27852) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16652) * $signed(input_fmap_109[7:0]) +
	( 16'sd 17029) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16061) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7854) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19678) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30027) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30878) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26775) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6906) * $signed(input_fmap_118[7:0]) +
	( 16'sd 29324) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11935) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10690) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31307) * $signed(input_fmap_122[7:0]) +
	( 16'sd 17165) * $signed(input_fmap_123[7:0]) +
	( 13'sd 3252) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24349) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17697) * $signed(input_fmap_127[7:0]) +
	( 16'sd 24486) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17800) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1668) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14514) * $signed(input_fmap_131[7:0]) +
	( 16'sd 20886) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10505) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19577) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28625) * $signed(input_fmap_135[7:0]) +
	( 14'sd 6940) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11760) * $signed(input_fmap_137[7:0]) +
	( 14'sd 6480) * $signed(input_fmap_138[7:0]) +
	( 16'sd 25929) * $signed(input_fmap_139[7:0]) +
	( 16'sd 23292) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3234) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19307) * $signed(input_fmap_142[7:0]) +
	( 16'sd 22196) * $signed(input_fmap_143[7:0]) +
	( 14'sd 8016) * $signed(input_fmap_144[7:0]) +
	( 16'sd 30126) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7346) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19133) * $signed(input_fmap_147[7:0]) +
	( 15'sd 10679) * $signed(input_fmap_148[7:0]) +
	( 10'sd 402) * $signed(input_fmap_149[7:0]) +
	( 12'sd 1285) * $signed(input_fmap_150[7:0]) +
	( 15'sd 13374) * $signed(input_fmap_151[7:0]) +
	( 12'sd 1898) * $signed(input_fmap_152[7:0]) +
	( 7'sd 37) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22889) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28746) * $signed(input_fmap_155[7:0]) +
	( 15'sd 12917) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23827) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8401) * $signed(input_fmap_158[7:0]) +
	( 15'sd 9442) * $signed(input_fmap_159[7:0]) +
	( 15'sd 14629) * $signed(input_fmap_160[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_161[7:0]) +
	( 16'sd 17389) * $signed(input_fmap_162[7:0]) +
	( 15'sd 9365) * $signed(input_fmap_163[7:0]) +
	( 15'sd 11904) * $signed(input_fmap_164[7:0]) +
	( 15'sd 16300) * $signed(input_fmap_165[7:0]) +
	( 15'sd 11781) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31158) * $signed(input_fmap_167[7:0]) +
	( 15'sd 13218) * $signed(input_fmap_168[7:0]) +
	( 15'sd 13584) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5360) * $signed(input_fmap_170[7:0]) +
	( 11'sd 729) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6952) * $signed(input_fmap_172[7:0]) +
	( 15'sd 9197) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7334) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4926) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10487) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7336) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31509) * $signed(input_fmap_178[7:0]) +
	( 14'sd 8023) * $signed(input_fmap_179[7:0]) +
	( 13'sd 4069) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30677) * $signed(input_fmap_181[7:0]) +
	( 14'sd 7316) * $signed(input_fmap_182[7:0]) +
	( 14'sd 8142) * $signed(input_fmap_183[7:0]) +
	( 13'sd 2221) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27938) * $signed(input_fmap_185[7:0]) +
	( 16'sd 31958) * $signed(input_fmap_186[7:0]) +
	( 16'sd 31186) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1425) * $signed(input_fmap_188[7:0]) +
	( 16'sd 21606) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28332) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24255) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12065) * $signed(input_fmap_193[7:0]) +
	( 16'sd 17133) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17448) * $signed(input_fmap_195[7:0]) +
	( 15'sd 13331) * $signed(input_fmap_196[7:0]) +
	( 16'sd 18426) * $signed(input_fmap_197[7:0]) +
	( 16'sd 19220) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29103) * $signed(input_fmap_199[7:0]) +
	( 16'sd 26973) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27377) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21933) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2934) * $signed(input_fmap_205[7:0]) +
	( 16'sd 23897) * $signed(input_fmap_206[7:0]) +
	( 14'sd 4619) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28727) * $signed(input_fmap_208[7:0]) +
	( 16'sd 28209) * $signed(input_fmap_209[7:0]) +
	( 16'sd 28623) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17389) * $signed(input_fmap_211[7:0]) +
	( 16'sd 28205) * $signed(input_fmap_212[7:0]) +
	( 15'sd 13794) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15887) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22420) * $signed(input_fmap_215[7:0]) +
	( 15'sd 15741) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_217[7:0]) +
	( 15'sd 14817) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5026) * $signed(input_fmap_219[7:0]) +
	( 16'sd 32423) * $signed(input_fmap_220[7:0]) +
	( 15'sd 8727) * $signed(input_fmap_221[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17987) * $signed(input_fmap_224[7:0]) +
	( 16'sd 29470) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32529) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27678) * $signed(input_fmap_227[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_228[7:0]) +
	( 11'sd 849) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6198) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10058) * $signed(input_fmap_231[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_233[7:0]) +
	( 15'sd 8927) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22422) * $signed(input_fmap_235[7:0]) +
	( 13'sd 3927) * $signed(input_fmap_236[7:0]) +
	( 15'sd 16203) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14799) * $signed(input_fmap_238[7:0]) +
	( 16'sd 27599) * $signed(input_fmap_239[7:0]) +
	( 14'sd 5974) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18817) * $signed(input_fmap_241[7:0]) +
	( 15'sd 10016) * $signed(input_fmap_242[7:0]) +
	( 13'sd 3109) * $signed(input_fmap_243[7:0]) +
	( 16'sd 17831) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28994) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30101) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21658) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3569) * $signed(input_fmap_249[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_250[7:0]) +
	( 16'sd 28040) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4897) * $signed(input_fmap_252[7:0]) +
	( 12'sd 1568) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10865) * $signed(input_fmap_254[7:0]) +
	( 12'sd 1412) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_194;
assign conv_mac_194 = 
	( 15'sd 13574) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23655) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9993) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6693) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20594) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27256) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31705) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20513) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30444) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2831) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27951) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24093) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21102) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10730) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4721) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31406) * $signed(input_fmap_15[7:0]) +
	( 16'sd 26339) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30139) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28749) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11562) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29198) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10689) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7023) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26334) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26667) * $signed(input_fmap_24[7:0]) +
	( 16'sd 28417) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8252) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31866) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11630) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4796) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5245) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19176) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17703) * $signed(input_fmap_32[7:0]) +
	( 16'sd 32128) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19082) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1239) * $signed(input_fmap_35[7:0]) +
	( 16'sd 24760) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10991) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15186) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20343) * $signed(input_fmap_39[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12389) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30066) * $signed(input_fmap_42[7:0]) +
	( 16'sd 29905) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20101) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11611) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28007) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27210) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26884) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30181) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11533) * $signed(input_fmap_52[7:0]) +
	( 16'sd 21899) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15012) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30922) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26799) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22959) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2472) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21806) * $signed(input_fmap_59[7:0]) +
	( 15'sd 14345) * $signed(input_fmap_60[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14420) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27321) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11870) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29036) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25789) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6074) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19271) * $signed(input_fmap_68[7:0]) +
	( 11'sd 740) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27267) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24810) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17435) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25880) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29014) * $signed(input_fmap_75[7:0]) +
	( 16'sd 32095) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19596) * $signed(input_fmap_77[7:0]) +
	( 15'sd 15087) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12750) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26891) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25308) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7126) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20299) * $signed(input_fmap_83[7:0]) +
	( 16'sd 32721) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10076) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31562) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5060) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2070) * $signed(input_fmap_88[7:0]) +
	( 16'sd 21838) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13722) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8364) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27964) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10208) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12472) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29701) * $signed(input_fmap_95[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10641) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2417) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25648) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13087) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27284) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3102) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13932) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16735) * $signed(input_fmap_104[7:0]) +
	( 15'sd 12487) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28452) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10593) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18722) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13996) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3973) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15761) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21130) * $signed(input_fmap_113[7:0]) +
	( 15'sd 8651) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24706) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6564) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26066) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15129) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3250) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17613) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15470) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10317) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30469) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18065) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26643) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2732) * $signed(input_fmap_126[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_127[7:0]) +
	( 16'sd 19122) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31667) * $signed(input_fmap_129[7:0]) +
	( 11'sd 810) * $signed(input_fmap_130[7:0]) +
	( 16'sd 16673) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25743) * $signed(input_fmap_132[7:0]) +
	( 15'sd 14054) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3261) * $signed(input_fmap_134[7:0]) +
	( 14'sd 4344) * $signed(input_fmap_135[7:0]) +
	( 16'sd 20010) * $signed(input_fmap_136[7:0]) +
	( 16'sd 31082) * $signed(input_fmap_137[7:0]) +
	( 15'sd 15595) * $signed(input_fmap_138[7:0]) +
	( 12'sd 1634) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9341) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13688) * $signed(input_fmap_141[7:0]) +
	( 16'sd 17234) * $signed(input_fmap_142[7:0]) +
	( 16'sd 29719) * $signed(input_fmap_143[7:0]) +
	( 15'sd 12097) * $signed(input_fmap_144[7:0]) +
	( 13'sd 3413) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29787) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30955) * $signed(input_fmap_147[7:0]) +
	( 16'sd 18025) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25008) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_150[7:0]) +
	( 16'sd 26896) * $signed(input_fmap_151[7:0]) +
	( 16'sd 18703) * $signed(input_fmap_152[7:0]) +
	( 16'sd 18696) * $signed(input_fmap_153[7:0]) +
	( 15'sd 13244) * $signed(input_fmap_154[7:0]) +
	( 16'sd 16551) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18232) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18202) * $signed(input_fmap_157[7:0]) +
	( 16'sd 31268) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5930) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22248) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31075) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_162[7:0]) +
	( 14'sd 6751) * $signed(input_fmap_163[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_164[7:0]) +
	( 16'sd 21323) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22216) * $signed(input_fmap_166[7:0]) +
	( 11'sd 598) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29888) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_169[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_170[7:0]) +
	( 14'sd 6397) * $signed(input_fmap_171[7:0]) +
	( 16'sd 25024) * $signed(input_fmap_172[7:0]) +
	( 15'sd 10815) * $signed(input_fmap_173[7:0]) +
	( 16'sd 24154) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1162) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10849) * $signed(input_fmap_176[7:0]) +
	( 16'sd 23063) * $signed(input_fmap_177[7:0]) +
	( 14'sd 8136) * $signed(input_fmap_178[7:0]) +
	( 8'sd 82) * $signed(input_fmap_179[7:0]) +
	( 15'sd 14463) * $signed(input_fmap_180[7:0]) +
	( 14'sd 5305) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30258) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5490) * $signed(input_fmap_183[7:0]) +
	( 16'sd 19885) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6001) * $signed(input_fmap_185[7:0]) +
	( 16'sd 27407) * $signed(input_fmap_186[7:0]) +
	( 16'sd 29817) * $signed(input_fmap_187[7:0]) +
	( 14'sd 7375) * $signed(input_fmap_188[7:0]) +
	( 13'sd 4041) * $signed(input_fmap_189[7:0]) +
	( 14'sd 6403) * $signed(input_fmap_190[7:0]) +
	( 15'sd 9529) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22315) * $signed(input_fmap_192[7:0]) +
	( 16'sd 31739) * $signed(input_fmap_193[7:0]) +
	( 16'sd 28819) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25356) * $signed(input_fmap_196[7:0]) +
	( 14'sd 6217) * $signed(input_fmap_197[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16267) * $signed(input_fmap_199[7:0]) +
	( 11'sd 957) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12410) * $signed(input_fmap_201[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_202[7:0]) +
	( 16'sd 27272) * $signed(input_fmap_203[7:0]) +
	( 12'sd 1489) * $signed(input_fmap_204[7:0]) +
	( 15'sd 14276) * $signed(input_fmap_205[7:0]) +
	( 12'sd 1413) * $signed(input_fmap_206[7:0]) +
	( 15'sd 15688) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6876) * $signed(input_fmap_208[7:0]) +
	( 16'sd 21333) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10317) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1629) * $signed(input_fmap_212[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_214[7:0]) +
	( 16'sd 24946) * $signed(input_fmap_215[7:0]) +
	( 16'sd 25893) * $signed(input_fmap_216[7:0]) +
	( 16'sd 31862) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22026) * $signed(input_fmap_218[7:0]) +
	( 16'sd 22744) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24107) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25270) * $signed(input_fmap_221[7:0]) +
	( 15'sd 8836) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15707) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17342) * $signed(input_fmap_224[7:0]) +
	( 16'sd 32405) * $signed(input_fmap_225[7:0]) +
	( 11'sd 673) * $signed(input_fmap_226[7:0]) +
	( 16'sd 16661) * $signed(input_fmap_227[7:0]) +
	( 14'sd 5792) * $signed(input_fmap_228[7:0]) +
	( 16'sd 28034) * $signed(input_fmap_229[7:0]) +
	( 13'sd 4028) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10959) * $signed(input_fmap_231[7:0]) +
	( 16'sd 30206) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27305) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23779) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26803) * $signed(input_fmap_235[7:0]) +
	( 16'sd 32603) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19156) * $signed(input_fmap_237[7:0]) +
	( 16'sd 16504) * $signed(input_fmap_238[7:0]) +
	( 15'sd 12726) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9699) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21279) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28870) * $signed(input_fmap_242[7:0]) +
	( 16'sd 32204) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19343) * $signed(input_fmap_244[7:0]) +
	( 16'sd 21243) * $signed(input_fmap_245[7:0]) +
	( 16'sd 32161) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9347) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1244) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28644) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25756) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13255) * $signed(input_fmap_251[7:0]) +
	( 16'sd 19405) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25777) * $signed(input_fmap_253[7:0]) +
	( 9'sd 210) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11236) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_195;
assign conv_mac_195 = 
	( 16'sd 31365) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23779) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27467) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28402) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9987) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23738) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4267) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1093) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17425) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10050) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9300) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20382) * $signed(input_fmap_11[7:0]) +
	( 16'sd 26328) * $signed(input_fmap_12[7:0]) +
	( 16'sd 17840) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20480) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10896) * $signed(input_fmap_15[7:0]) +
	( 14'sd 7011) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1497) * $signed(input_fmap_18[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30788) * $signed(input_fmap_20[7:0]) +
	( 11'sd 788) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31024) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24777) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20409) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17185) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29486) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31313) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30272) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7483) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15704) * $signed(input_fmap_30[7:0]) +
	( 15'sd 10252) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_32[7:0]) +
	( 11'sd 824) * $signed(input_fmap_33[7:0]) +
	( 16'sd 17296) * $signed(input_fmap_34[7:0]) +
	( 16'sd 31124) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9010) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18356) * $signed(input_fmap_37[7:0]) +
	( 11'sd 591) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4447) * $signed(input_fmap_39[7:0]) +
	( 14'sd 5304) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15114) * $signed(input_fmap_41[7:0]) +
	( 10'sd 384) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_43[7:0]) +
	( 10'sd 339) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30891) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22984) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17396) * $signed(input_fmap_47[7:0]) +
	( 14'sd 5575) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19083) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26272) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13060) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13829) * $signed(input_fmap_53[7:0]) +
	( 16'sd 32090) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15859) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3545) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1377) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1660) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12175) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18879) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31825) * $signed(input_fmap_64[7:0]) +
	( 16'sd 26959) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29067) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28090) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30073) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1256) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4970) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24966) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11814) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3439) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21284) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13687) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12632) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31537) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29913) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30298) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27652) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6314) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6784) * $signed(input_fmap_82[7:0]) +
	( 16'sd 16448) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5668) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6159) * $signed(input_fmap_85[7:0]) +
	( 15'sd 12307) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20468) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16048) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19627) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15912) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30365) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9989) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11456) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9128) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20986) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14350) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25614) * $signed(input_fmap_98[7:0]) +
	( 12'sd 1959) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27186) * $signed(input_fmap_100[7:0]) +
	( 13'sd 2293) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1259) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9288) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24360) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17246) * $signed(input_fmap_105[7:0]) +
	( 15'sd 10598) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25892) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14720) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4204) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9062) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3279) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10716) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9862) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2962) * $signed(input_fmap_115[7:0]) +
	( 14'sd 5873) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20631) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_118[7:0]) +
	( 14'sd 8018) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7324) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6721) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19284) * $signed(input_fmap_122[7:0]) +
	( 11'sd 713) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10312) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20674) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18856) * $signed(input_fmap_127[7:0]) +
	( 16'sd 28913) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1536) * $signed(input_fmap_129[7:0]) +
	( 15'sd 9285) * $signed(input_fmap_130[7:0]) +
	( 16'sd 29244) * $signed(input_fmap_131[7:0]) +
	( 14'sd 6127) * $signed(input_fmap_132[7:0]) +
	( 16'sd 18731) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18824) * $signed(input_fmap_134[7:0]) +
	( 16'sd 24353) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1513) * $signed(input_fmap_136[7:0]) +
	( 11'sd 721) * $signed(input_fmap_137[7:0]) +
	( 13'sd 2642) * $signed(input_fmap_138[7:0]) +
	( 16'sd 19776) * $signed(input_fmap_139[7:0]) +
	( 13'sd 2368) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19945) * $signed(input_fmap_141[7:0]) +
	( 9'sd 247) * $signed(input_fmap_142[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11634) * $signed(input_fmap_144[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_145[7:0]) +
	( 14'sd 5023) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27392) * $signed(input_fmap_147[7:0]) +
	( 14'sd 7853) * $signed(input_fmap_148[7:0]) +
	( 13'sd 3385) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9288) * $signed(input_fmap_150[7:0]) +
	( 16'sd 27581) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7971) * $signed(input_fmap_152[7:0]) +
	( 16'sd 30402) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25381) * $signed(input_fmap_154[7:0]) +
	( 13'sd 2679) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25499) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20112) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11096) * $signed(input_fmap_158[7:0]) +
	( 15'sd 10100) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6906) * $signed(input_fmap_160[7:0]) +
	( 15'sd 8717) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29921) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15299) * $signed(input_fmap_163[7:0]) +
	( 16'sd 32677) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19304) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22685) * $signed(input_fmap_166[7:0]) +
	( 15'sd 12218) * $signed(input_fmap_167[7:0]) +
	( 16'sd 25521) * $signed(input_fmap_168[7:0]) +
	( 16'sd 32666) * $signed(input_fmap_169[7:0]) +
	( 16'sd 25905) * $signed(input_fmap_170[7:0]) +
	( 16'sd 21149) * $signed(input_fmap_171[7:0]) +
	( 15'sd 11738) * $signed(input_fmap_172[7:0]) +
	( 14'sd 7925) * $signed(input_fmap_173[7:0]) +
	( 15'sd 16218) * $signed(input_fmap_174[7:0]) +
	( 16'sd 19288) * $signed(input_fmap_175[7:0]) +
	( 16'sd 25506) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6872) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32312) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25161) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21994) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30273) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6331) * $signed(input_fmap_182[7:0]) +
	( 15'sd 16259) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11031) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6529) * $signed(input_fmap_186[7:0]) +
	( 16'sd 31665) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_188[7:0]) +
	( 16'sd 23432) * $signed(input_fmap_189[7:0]) +
	( 15'sd 12783) * $signed(input_fmap_190[7:0]) +
	( 16'sd 16728) * $signed(input_fmap_191[7:0]) +
	( 15'sd 9329) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11546) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14586) * $signed(input_fmap_194[7:0]) +
	( 14'sd 7488) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6399) * $signed(input_fmap_196[7:0]) +
	( 12'sd 1042) * $signed(input_fmap_197[7:0]) +
	( 16'sd 21498) * $signed(input_fmap_198[7:0]) +
	( 11'sd 804) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29319) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11372) * $signed(input_fmap_201[7:0]) +
	( 16'sd 16768) * $signed(input_fmap_202[7:0]) +
	( 14'sd 4796) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12981) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30175) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9525) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13931) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12844) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18788) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5118) * $signed(input_fmap_210[7:0]) +
	( 14'sd 4401) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11632) * $signed(input_fmap_212[7:0]) +
	( 16'sd 20611) * $signed(input_fmap_213[7:0]) +
	( 13'sd 3168) * $signed(input_fmap_214[7:0]) +
	( 16'sd 20299) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20639) * $signed(input_fmap_216[7:0]) +
	( 15'sd 8197) * $signed(input_fmap_217[7:0]) +
	( 16'sd 27901) * $signed(input_fmap_218[7:0]) +
	( 12'sd 1175) * $signed(input_fmap_219[7:0]) +
	( 15'sd 10500) * $signed(input_fmap_220[7:0]) +
	( 15'sd 10970) * $signed(input_fmap_221[7:0]) +
	( 16'sd 22411) * $signed(input_fmap_222[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14424) * $signed(input_fmap_224[7:0]) +
	( 15'sd 12788) * $signed(input_fmap_225[7:0]) +
	( 16'sd 20861) * $signed(input_fmap_226[7:0]) +
	( 16'sd 18442) * $signed(input_fmap_227[7:0]) +
	( 11'sd 778) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6994) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6220) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7363) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9402) * $signed(input_fmap_232[7:0]) +
	( 16'sd 30488) * $signed(input_fmap_233[7:0]) +
	( 16'sd 30782) * $signed(input_fmap_234[7:0]) +
	( 15'sd 9282) * $signed(input_fmap_235[7:0]) +
	( 16'sd 21344) * $signed(input_fmap_236[7:0]) +
	( 16'sd 27761) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17752) * $signed(input_fmap_238[7:0]) +
	( 14'sd 6613) * $signed(input_fmap_239[7:0]) +
	( 15'sd 12646) * $signed(input_fmap_240[7:0]) +
	( 14'sd 6749) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23488) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6329) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30743) * $signed(input_fmap_244[7:0]) +
	( 14'sd 5969) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11050) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17807) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18977) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30622) * $signed(input_fmap_249[7:0]) +
	( 16'sd 31945) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19381) * $signed(input_fmap_251[7:0]) +
	( 15'sd 15169) * $signed(input_fmap_252[7:0]) +
	( 15'sd 8984) * $signed(input_fmap_253[7:0]) +
	( 15'sd 12689) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26141) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_196;
assign conv_mac_196 = 
	( 15'sd 10745) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29712) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12749) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2462) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29958) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9365) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12757) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21323) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23977) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7347) * $signed(input_fmap_9[7:0]) +
	( 11'sd 1005) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9902) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25419) * $signed(input_fmap_12[7:0]) +
	( 16'sd 32294) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27478) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1192) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27499) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_17[7:0]) +
	( 16'sd 18583) * $signed(input_fmap_18[7:0]) +
	( 15'sd 15914) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23520) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10020) * $signed(input_fmap_21[7:0]) +
	( 10'sd 356) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11097) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11353) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12615) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26317) * $signed(input_fmap_26[7:0]) +
	( 9'sd 250) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19639) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24473) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1786) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24206) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4441) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1601) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26781) * $signed(input_fmap_34[7:0]) +
	( 10'sd 506) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4268) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28770) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7836) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17509) * $signed(input_fmap_39[7:0]) +
	( 16'sd 30382) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11502) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16256) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2345) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21876) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23868) * $signed(input_fmap_46[7:0]) +
	( 14'sd 7441) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30692) * $signed(input_fmap_48[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15811) * $signed(input_fmap_52[7:0]) +
	( 11'sd 867) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31310) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15798) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17675) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4298) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24126) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19161) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31899) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21442) * $signed(input_fmap_61[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14677) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18247) * $signed(input_fmap_64[7:0]) +
	( 15'sd 13820) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18200) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12653) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1960) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26145) * $signed(input_fmap_69[7:0]) +
	( 15'sd 9789) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16710) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_72[7:0]) +
	( 16'sd 31342) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29381) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13072) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23022) * $signed(input_fmap_76[7:0]) +
	( 11'sd 772) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13089) * $signed(input_fmap_79[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10438) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6052) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10511) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4821) * $signed(input_fmap_84[7:0]) +
	( 16'sd 26380) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18510) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_87[7:0]) +
	( 16'sd 32655) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7717) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17083) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15558) * $signed(input_fmap_91[7:0]) +
	( 15'sd 16229) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15239) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12412) * $signed(input_fmap_94[7:0]) +
	( 16'sd 25440) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12543) * $signed(input_fmap_96[7:0]) +
	( 15'sd 10803) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21367) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9090) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29767) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6645) * $signed(input_fmap_101[7:0]) +
	( 16'sd 25618) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23376) * $signed(input_fmap_104[7:0]) +
	( 13'sd 3130) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3828) * $signed(input_fmap_106[7:0]) +
	( 16'sd 20408) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8283) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11425) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23423) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22396) * $signed(input_fmap_112[7:0]) +
	( 11'sd 603) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14926) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23762) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3865) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15494) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4631) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20330) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6294) * $signed(input_fmap_120[7:0]) +
	( 14'sd 8018) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12044) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6134) * $signed(input_fmap_123[7:0]) +
	( 14'sd 6902) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3405) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6454) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4938) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13877) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6204) * $signed(input_fmap_130[7:0]) +
	( 16'sd 20469) * $signed(input_fmap_131[7:0]) +
	( 16'sd 30739) * $signed(input_fmap_132[7:0]) +
	( 16'sd 23419) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24167) * $signed(input_fmap_134[7:0]) +
	( 15'sd 13522) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25275) * $signed(input_fmap_136[7:0]) +
	( 13'sd 2525) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7039) * $signed(input_fmap_138[7:0]) +
	( 16'sd 26680) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28074) * $signed(input_fmap_140[7:0]) +
	( 16'sd 25217) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19025) * $signed(input_fmap_142[7:0]) +
	( 15'sd 14774) * $signed(input_fmap_143[7:0]) +
	( 15'sd 12999) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23848) * $signed(input_fmap_145[7:0]) +
	( 15'sd 8685) * $signed(input_fmap_146[7:0]) +
	( 14'sd 4963) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_148[7:0]) +
	( 15'sd 13502) * $signed(input_fmap_149[7:0]) +
	( 12'sd 1423) * $signed(input_fmap_150[7:0]) +
	( 15'sd 15837) * $signed(input_fmap_151[7:0]) +
	( 16'sd 17340) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23388) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22598) * $signed(input_fmap_154[7:0]) +
	( 13'sd 4006) * $signed(input_fmap_155[7:0]) +
	( 16'sd 30160) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6224) * $signed(input_fmap_157[7:0]) +
	( 14'sd 6056) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26936) * $signed(input_fmap_159[7:0]) +
	( 16'sd 17383) * $signed(input_fmap_160[7:0]) +
	( 13'sd 3295) * $signed(input_fmap_161[7:0]) +
	( 13'sd 3136) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9480) * $signed(input_fmap_164[7:0]) +
	( 15'sd 8254) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19905) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26151) * $signed(input_fmap_167[7:0]) +
	( 16'sd 16689) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28432) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24404) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3411) * $signed(input_fmap_172[7:0]) +
	( 13'sd 3004) * $signed(input_fmap_173[7:0]) +
	( 16'sd 20468) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17628) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15509) * $signed(input_fmap_176[7:0]) +
	( 16'sd 19075) * $signed(input_fmap_177[7:0]) +
	( 16'sd 28155) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22866) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24457) * $signed(input_fmap_180[7:0]) +
	( 16'sd 27687) * $signed(input_fmap_181[7:0]) +
	( 16'sd 22372) * $signed(input_fmap_182[7:0]) +
	( 12'sd 1125) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13000) * $signed(input_fmap_184[7:0]) +
	( 16'sd 23824) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23062) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5259) * $signed(input_fmap_187[7:0]) +
	( 16'sd 19003) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_189[7:0]) +
	( 16'sd 21664) * $signed(input_fmap_190[7:0]) +
	( 15'sd 9923) * $signed(input_fmap_191[7:0]) +
	( 10'sd 401) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5687) * $signed(input_fmap_193[7:0]) +
	( 14'sd 5754) * $signed(input_fmap_194[7:0]) +
	( 15'sd 15707) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7004) * $signed(input_fmap_196[7:0]) +
	( 16'sd 27300) * $signed(input_fmap_197[7:0]) +
	( 15'sd 13825) * $signed(input_fmap_198[7:0]) +
	( 10'sd 354) * $signed(input_fmap_199[7:0]) +
	( 13'sd 2278) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18375) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7796) * $signed(input_fmap_202[7:0]) +
	( 16'sd 20462) * $signed(input_fmap_203[7:0]) +
	( 15'sd 13092) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11247) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21308) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6734) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18960) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_210[7:0]) +
	( 16'sd 29344) * $signed(input_fmap_211[7:0]) +
	( 16'sd 16709) * $signed(input_fmap_212[7:0]) +
	( 16'sd 26924) * $signed(input_fmap_213[7:0]) +
	( 16'sd 26673) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11646) * $signed(input_fmap_215[7:0]) +
	( 10'sd 440) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25053) * $signed(input_fmap_217[7:0]) +
	( 15'sd 11467) * $signed(input_fmap_218[7:0]) +
	( 13'sd 2340) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22682) * $signed(input_fmap_220[7:0]) +
	( 13'sd 2167) * $signed(input_fmap_221[7:0]) +
	( 16'sd 29741) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9150) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30181) * $signed(input_fmap_224[7:0]) +
	( 16'sd 28872) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6784) * $signed(input_fmap_226[7:0]) +
	( 15'sd 15518) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31734) * $signed(input_fmap_228[7:0]) +
	( 15'sd 13412) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18940) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25156) * $signed(input_fmap_231[7:0]) +
	( 15'sd 13106) * $signed(input_fmap_232[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_233[7:0]) +
	( 16'sd 29190) * $signed(input_fmap_234[7:0]) +
	( 15'sd 11355) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30459) * $signed(input_fmap_236[7:0]) +
	( 12'sd 1871) * $signed(input_fmap_237[7:0]) +
	( 16'sd 25510) * $signed(input_fmap_238[7:0]) +
	( 16'sd 32458) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31847) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3523) * $signed(input_fmap_241[7:0]) +
	( 15'sd 8969) * $signed(input_fmap_242[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_243[7:0]) +
	( 15'sd 16076) * $signed(input_fmap_244[7:0]) +
	( 14'sd 4205) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15149) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30484) * $signed(input_fmap_247[7:0]) +
	( 16'sd 16955) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4951) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_250[7:0]) +
	( 16'sd 32137) * $signed(input_fmap_251[7:0]) +
	( 16'sd 31302) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29732) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26650) * $signed(input_fmap_254[7:0]) +
	( 13'sd 4025) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_197;
assign conv_mac_197 = 
	( 16'sd 28713) * $signed(input_fmap_0[7:0]) +
	( 16'sd 29048) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7149) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14208) * $signed(input_fmap_4[7:0]) +
	( 14'sd 5693) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24216) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32318) * $signed(input_fmap_8[7:0]) +
	( 16'sd 17539) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29160) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9933) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22151) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18368) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28735) * $signed(input_fmap_15[7:0]) +
	( 16'sd 18153) * $signed(input_fmap_16[7:0]) +
	( 13'sd 3535) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27233) * $signed(input_fmap_19[7:0]) +
	( 14'sd 6167) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5429) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14202) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23515) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32389) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22685) * $signed(input_fmap_25[7:0]) +
	( 6'sd 27) * $signed(input_fmap_26[7:0]) +
	( 16'sd 19995) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18956) * $signed(input_fmap_28[7:0]) +
	( 16'sd 30876) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23081) * $signed(input_fmap_30[7:0]) +
	( 16'sd 31433) * $signed(input_fmap_31[7:0]) +
	( 15'sd 16133) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26940) * $signed(input_fmap_33[7:0]) +
	( 12'sd 1957) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13314) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18473) * $signed(input_fmap_36[7:0]) +
	( 15'sd 12972) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13963) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32671) * $signed(input_fmap_40[7:0]) +
	( 13'sd 3311) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30707) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7900) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12133) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28771) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19492) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5932) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28824) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28544) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6212) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26877) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23126) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4257) * $signed(input_fmap_54[7:0]) +
	( 15'sd 16046) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1626) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25292) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28623) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31241) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8722) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27269) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20286) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25910) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19898) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16217) * $signed(input_fmap_65[7:0]) +
	( 16'sd 28307) * $signed(input_fmap_66[7:0]) +
	( 16'sd 30353) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3019) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16529) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7933) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20549) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19443) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21219) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19182) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20526) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7871) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27961) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18200) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29668) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12070) * $signed(input_fmap_81[7:0]) +
	( 11'sd 701) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19678) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11873) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19635) * $signed(input_fmap_85[7:0]) +
	( 16'sd 25120) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3498) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23681) * $signed(input_fmap_88[7:0]) +
	( 15'sd 15942) * $signed(input_fmap_89[7:0]) +
	( 16'sd 25037) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7497) * $signed(input_fmap_91[7:0]) +
	( 15'sd 14524) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8375) * $signed(input_fmap_93[7:0]) +
	( 15'sd 9519) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26873) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6450) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20711) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26406) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19826) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3019) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17738) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11706) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20314) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1291) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6527) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13066) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11504) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12488) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1645) * $signed(input_fmap_111[7:0]) +
	( 16'sd 32158) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21474) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_114[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18341) * $signed(input_fmap_116[7:0]) +
	( 10'sd 495) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12117) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25994) * $signed(input_fmap_120[7:0]) +
	( 15'sd 10941) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24502) * $signed(input_fmap_122[7:0]) +
	( 11'sd 585) * $signed(input_fmap_123[7:0]) +
	( 15'sd 8278) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16722) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21521) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29481) * $signed(input_fmap_127[7:0]) +
	( 16'sd 21364) * $signed(input_fmap_128[7:0]) +
	( 16'sd 25172) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10836) * $signed(input_fmap_130[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11289) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21854) * $signed(input_fmap_133[7:0]) +
	( 16'sd 24416) * $signed(input_fmap_134[7:0]) +
	( 12'sd 1852) * $signed(input_fmap_135[7:0]) +
	( 15'sd 12561) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7330) * $signed(input_fmap_138[7:0]) +
	( 14'sd 7379) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28924) * $signed(input_fmap_140[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11369) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26328) * $signed(input_fmap_143[7:0]) +
	( 16'sd 25598) * $signed(input_fmap_144[7:0]) +
	( 16'sd 18288) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3223) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18152) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11400) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25904) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31805) * $signed(input_fmap_150[7:0]) +
	( 15'sd 15230) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6703) * $signed(input_fmap_152[7:0]) +
	( 13'sd 3889) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22488) * $signed(input_fmap_154[7:0]) +
	( 16'sd 29026) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17318) * $signed(input_fmap_156[7:0]) +
	( 16'sd 19622) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9578) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4933) * $signed(input_fmap_159[7:0]) +
	( 15'sd 10072) * $signed(input_fmap_160[7:0]) +
	( 15'sd 16009) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21536) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24418) * $signed(input_fmap_163[7:0]) +
	( 10'sd 378) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30702) * $signed(input_fmap_165[7:0]) +
	( 16'sd 23699) * $signed(input_fmap_166[7:0]) +
	( 12'sd 2034) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20314) * $signed(input_fmap_169[7:0]) +
	( 16'sd 29868) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31441) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19513) * $signed(input_fmap_172[7:0]) +
	( 13'sd 2703) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14509) * $signed(input_fmap_174[7:0]) +
	( 16'sd 18622) * $signed(input_fmap_175[7:0]) +
	( 16'sd 31755) * $signed(input_fmap_176[7:0]) +
	( 16'sd 16520) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17919) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5450) * $signed(input_fmap_179[7:0]) +
	( 16'sd 18963) * $signed(input_fmap_180[7:0]) +
	( 16'sd 17874) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26839) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5388) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24232) * $signed(input_fmap_185[7:0]) +
	( 16'sd 20266) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22225) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21608) * $signed(input_fmap_188[7:0]) +
	( 15'sd 15181) * $signed(input_fmap_189[7:0]) +
	( 15'sd 16113) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5640) * $signed(input_fmap_191[7:0]) +
	( 15'sd 8927) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30877) * $signed(input_fmap_193[7:0]) +
	( 14'sd 4592) * $signed(input_fmap_194[7:0]) +
	( 16'sd 18973) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17251) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11211) * $signed(input_fmap_197[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_198[7:0]) +
	( 16'sd 22106) * $signed(input_fmap_199[7:0]) +
	( 16'sd 24707) * $signed(input_fmap_200[7:0]) +
	( 14'sd 7816) * $signed(input_fmap_201[7:0]) +
	( 16'sd 20990) * $signed(input_fmap_202[7:0]) +
	( 15'sd 15749) * $signed(input_fmap_203[7:0]) +
	( 11'sd 923) * $signed(input_fmap_204[7:0]) +
	( 16'sd 32286) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27443) * $signed(input_fmap_206[7:0]) +
	( 16'sd 19887) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4607) * $signed(input_fmap_208[7:0]) +
	( 13'sd 2910) * $signed(input_fmap_209[7:0]) +
	( 16'sd 25244) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28503) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17948) * $signed(input_fmap_212[7:0]) +
	( 16'sd 25182) * $signed(input_fmap_213[7:0]) +
	( 16'sd 26350) * $signed(input_fmap_214[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_215[7:0]) +
	( 16'sd 22435) * $signed(input_fmap_216[7:0]) +
	( 14'sd 5963) * $signed(input_fmap_217[7:0]) +
	( 13'sd 2403) * $signed(input_fmap_218[7:0]) +
	( 16'sd 31338) * $signed(input_fmap_219[7:0]) +
	( 16'sd 18321) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27469) * $signed(input_fmap_221[7:0]) +
	( 11'sd 799) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22434) * $signed(input_fmap_223[7:0]) +
	( 13'sd 2722) * $signed(input_fmap_224[7:0]) +
	( 14'sd 4389) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7138) * $signed(input_fmap_226[7:0]) +
	( 16'sd 25728) * $signed(input_fmap_227[7:0]) +
	( 10'sd 414) * $signed(input_fmap_228[7:0]) +
	( 15'sd 14415) * $signed(input_fmap_229[7:0]) +
	( 15'sd 13213) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3360) * $signed(input_fmap_231[7:0]) +
	( 14'sd 6599) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28256) * $signed(input_fmap_233[7:0]) +
	( 15'sd 9677) * $signed(input_fmap_234[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_235[7:0]) +
	( 14'sd 4701) * $signed(input_fmap_236[7:0]) +
	( 16'sd 25414) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23186) * $signed(input_fmap_238[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_239[7:0]) +
	( 16'sd 30578) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5667) * $signed(input_fmap_241[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28977) * $signed(input_fmap_243[7:0]) +
	( 16'sd 26055) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24427) * $signed(input_fmap_245[7:0]) +
	( 16'sd 26501) * $signed(input_fmap_246[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_247[7:0]) +
	( 16'sd 28874) * $signed(input_fmap_248[7:0]) +
	( 16'sd 26025) * $signed(input_fmap_249[7:0]) +
	( 12'sd 1186) * $signed(input_fmap_250[7:0]) +
	( 15'sd 9025) * $signed(input_fmap_251[7:0]) +
	( 15'sd 15821) * $signed(input_fmap_252[7:0]) +
	( 16'sd 30904) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26261) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24115) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_198;
assign conv_mac_198 = 
	( 16'sd 26559) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16366) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1733) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9271) * $signed(input_fmap_3[7:0]) +
	( 15'sd 10898) * $signed(input_fmap_4[7:0]) +
	( 11'sd 764) * $signed(input_fmap_5[7:0]) +
	( 14'sd 5233) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20707) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13521) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4874) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16713) * $signed(input_fmap_10[7:0]) +
	( 16'sd 30837) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23316) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8989) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32757) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31557) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30283) * $signed(input_fmap_16[7:0]) +
	( 14'sd 5769) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5599) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4547) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31388) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25988) * $signed(input_fmap_21[7:0]) +
	( 16'sd 17284) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30202) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30124) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22548) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30310) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30649) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24260) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19174) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15147) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27605) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10785) * $signed(input_fmap_33[7:0]) +
	( 16'sd 16443) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11219) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21425) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8423) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9295) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19185) * $signed(input_fmap_39[7:0]) +
	( 15'sd 9900) * $signed(input_fmap_40[7:0]) +
	( 10'sd 380) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16397) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2203) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6297) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16047) * $signed(input_fmap_45[7:0]) +
	( 16'sd 18841) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21445) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21247) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32115) * $signed(input_fmap_49[7:0]) +
	( 13'sd 3710) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28623) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32344) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16643) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17801) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24551) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16494) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29276) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19789) * $signed(input_fmap_58[7:0]) +
	( 15'sd 16216) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22824) * $signed(input_fmap_60[7:0]) +
	( 14'sd 8085) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6364) * $signed(input_fmap_62[7:0]) +
	( 16'sd 19655) * $signed(input_fmap_63[7:0]) +
	( 15'sd 8799) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10590) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25455) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31435) * $signed(input_fmap_67[7:0]) +
	( 15'sd 10635) * $signed(input_fmap_68[7:0]) +
	( 16'sd 22605) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6877) * $signed(input_fmap_70[7:0]) +
	( 11'sd 971) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19976) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24468) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15942) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3476) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32103) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29545) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14649) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31981) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1899) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8210) * $signed(input_fmap_82[7:0]) +
	( 15'sd 16227) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1093) * $signed(input_fmap_84[7:0]) +
	( 16'sd 20873) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9093) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24381) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11062) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1404) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3476) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16308) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4442) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12155) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7420) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4674) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30161) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17580) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6773) * $signed(input_fmap_102[7:0]) +
	( 15'sd 14170) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31677) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16898) * $signed(input_fmap_105[7:0]) +
	( 10'sd 337) * $signed(input_fmap_106[7:0]) +
	( 15'sd 9223) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12773) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26383) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22407) * $signed(input_fmap_110[7:0]) +
	( 14'sd 7184) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16034) * $signed(input_fmap_112[7:0]) +
	( 16'sd 23207) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7205) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24727) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20795) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23238) * $signed(input_fmap_117[7:0]) +
	( 16'sd 16651) * $signed(input_fmap_118[7:0]) +
	( 13'sd 3311) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8829) * $signed(input_fmap_120[7:0]) +
	( 15'sd 8355) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31440) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32479) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26607) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23121) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_128[7:0]) +
	( 13'sd 4077) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6226) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23396) * $signed(input_fmap_131[7:0]) +
	( 13'sd 3615) * $signed(input_fmap_132[7:0]) +
	( 16'sd 17245) * $signed(input_fmap_133[7:0]) +
	( 15'sd 10315) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23729) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30120) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9645) * $signed(input_fmap_137[7:0]) +
	( 16'sd 24797) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17559) * $signed(input_fmap_140[7:0]) +
	( 11'sd 905) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30203) * $signed(input_fmap_142[7:0]) +
	( 15'sd 9827) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19645) * $signed(input_fmap_144[7:0]) +
	( 16'sd 18586) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24267) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13988) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3407) * $signed(input_fmap_148[7:0]) +
	( 15'sd 10985) * $signed(input_fmap_149[7:0]) +
	( 16'sd 26150) * $signed(input_fmap_150[7:0]) +
	( 11'sd 592) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_152[7:0]) +
	( 16'sd 19820) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25788) * $signed(input_fmap_154[7:0]) +
	( 16'sd 26898) * $signed(input_fmap_155[7:0]) +
	( 14'sd 7320) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14160) * $signed(input_fmap_157[7:0]) +
	( 16'sd 16893) * $signed(input_fmap_158[7:0]) +
	( 15'sd 14495) * $signed(input_fmap_159[7:0]) +
	( 15'sd 10825) * $signed(input_fmap_160[7:0]) +
	( 16'sd 32619) * $signed(input_fmap_161[7:0]) +
	( 16'sd 17461) * $signed(input_fmap_162[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10036) * $signed(input_fmap_164[7:0]) +
	( 16'sd 24947) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18160) * $signed(input_fmap_166[7:0]) +
	( 13'sd 4011) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5225) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18966) * $signed(input_fmap_169[7:0]) +
	( 16'sd 19863) * $signed(input_fmap_170[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_171[7:0]) +
	( 16'sd 26634) * $signed(input_fmap_172[7:0]) +
	( 16'sd 16853) * $signed(input_fmap_173[7:0]) +
	( 15'sd 10574) * $signed(input_fmap_174[7:0]) +
	( 16'sd 18046) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21557) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22289) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2509) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3636) * $signed(input_fmap_179[7:0]) +
	( 15'sd 8226) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11686) * $signed(input_fmap_181[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_182[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9545) * $signed(input_fmap_184[7:0]) +
	( 16'sd 27122) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9815) * $signed(input_fmap_186[7:0]) +
	( 16'sd 26706) * $signed(input_fmap_187[7:0]) +
	( 16'sd 24485) * $signed(input_fmap_188[7:0]) +
	( 16'sd 20767) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4924) * $signed(input_fmap_190[7:0]) +
	( 15'sd 12628) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31667) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_193[7:0]) +
	( 13'sd 2208) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13791) * $signed(input_fmap_195[7:0]) +
	( 15'sd 11517) * $signed(input_fmap_196[7:0]) +
	( 16'sd 18659) * $signed(input_fmap_197[7:0]) +
	( 14'sd 4607) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28291) * $signed(input_fmap_199[7:0]) +
	( 16'sd 24748) * $signed(input_fmap_200[7:0]) +
	( 15'sd 16269) * $signed(input_fmap_201[7:0]) +
	( 16'sd 21342) * $signed(input_fmap_202[7:0]) +
	( 16'sd 18651) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29463) * $signed(input_fmap_205[7:0]) +
	( 16'sd 16411) * $signed(input_fmap_206[7:0]) +
	( 15'sd 15916) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15460) * $signed(input_fmap_208[7:0]) +
	( 16'sd 30986) * $signed(input_fmap_209[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28642) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1672) * $signed(input_fmap_212[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17010) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10901) * $signed(input_fmap_215[7:0]) +
	( 16'sd 26587) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30444) * $signed(input_fmap_217[7:0]) +
	( 15'sd 14135) * $signed(input_fmap_218[7:0]) +
	( 15'sd 11638) * $signed(input_fmap_219[7:0]) +
	( 14'sd 7753) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27863) * $signed(input_fmap_221[7:0]) +
	( 16'sd 21749) * $signed(input_fmap_222[7:0]) +
	( 15'sd 15809) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12253) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2476) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11676) * $signed(input_fmap_226[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4431) * $signed(input_fmap_228[7:0]) +
	( 16'sd 27815) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6181) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17176) * $signed(input_fmap_231[7:0]) +
	( 12'sd 1077) * $signed(input_fmap_232[7:0]) +
	( 15'sd 13724) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14915) * $signed(input_fmap_234[7:0]) +
	( 16'sd 30548) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2796) * $signed(input_fmap_236[7:0]) +
	( 14'sd 7979) * $signed(input_fmap_237[7:0]) +
	( 16'sd 24573) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22114) * $signed(input_fmap_239[7:0]) +
	( 13'sd 2655) * $signed(input_fmap_240[7:0]) +
	( 16'sd 27079) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15957) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2638) * $signed(input_fmap_243[7:0]) +
	( 16'sd 18496) * $signed(input_fmap_244[7:0]) +
	( 16'sd 29203) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10780) * $signed(input_fmap_246[7:0]) +
	( 15'sd 8662) * $signed(input_fmap_247[7:0]) +
	( 15'sd 14909) * $signed(input_fmap_248[7:0]) +
	( 16'sd 26558) * $signed(input_fmap_249[7:0]) +
	( 9'sd 196) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21613) * $signed(input_fmap_251[7:0]) +
	( 15'sd 15818) * $signed(input_fmap_252[7:0]) +
	( 15'sd 8321) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10611) * $signed(input_fmap_254[7:0]) +
	( 16'sd 29073) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_199;
assign conv_mac_199 = 
	( 15'sd 12040) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19991) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19445) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21446) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1637) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13883) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21593) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29182) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9862) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4518) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5609) * $signed(input_fmap_10[7:0]) +
	( 14'sd 7482) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24183) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31807) * $signed(input_fmap_13[7:0]) +
	( 16'sd 25171) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17913) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27768) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23565) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22411) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2882) * $signed(input_fmap_19[7:0]) +
	( 16'sd 30096) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16910) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23395) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19127) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21636) * $signed(input_fmap_24[7:0]) +
	( 16'sd 25911) * $signed(input_fmap_25[7:0]) +
	( 12'sd 1506) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20650) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1159) * $signed(input_fmap_28[7:0]) +
	( 16'sd 16420) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2157) * $signed(input_fmap_30[7:0]) +
	( 16'sd 26966) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18855) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15370) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27087) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16046) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22457) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11100) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2581) * $signed(input_fmap_38[7:0]) +
	( 15'sd 11959) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2521) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18705) * $signed(input_fmap_41[7:0]) +
	( 16'sd 20830) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11741) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26520) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23318) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12778) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1362) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7856) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8402) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31710) * $signed(input_fmap_51[7:0]) +
	( 15'sd 10393) * $signed(input_fmap_52[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6711) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9719) * $signed(input_fmap_55[7:0]) +
	( 16'sd 22806) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10507) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24125) * $signed(input_fmap_58[7:0]) +
	( 15'sd 8519) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32099) * $signed(input_fmap_60[7:0]) +
	( 14'sd 6522) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16731) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20259) * $signed(input_fmap_63[7:0]) +
	( 16'sd 32347) * $signed(input_fmap_64[7:0]) +
	( 16'sd 29665) * $signed(input_fmap_65[7:0]) +
	( 16'sd 19072) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5216) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14202) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25413) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10804) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30805) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14835) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4696) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22051) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26527) * $signed(input_fmap_78[7:0]) +
	( 16'sd 24063) * $signed(input_fmap_79[7:0]) +
	( 16'sd 28472) * $signed(input_fmap_80[7:0]) +
	( 11'sd 649) * $signed(input_fmap_81[7:0]) +
	( 16'sd 29636) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19604) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31949) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_85[7:0]) +
	( 14'sd 7097) * $signed(input_fmap_86[7:0]) +
	( 15'sd 11824) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30338) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9374) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3100) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17488) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5688) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2368) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24046) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17346) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30904) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21173) * $signed(input_fmap_98[7:0]) +
	( 16'sd 20398) * $signed(input_fmap_99[7:0]) +
	( 16'sd 29963) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23803) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1927) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2546) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16091) * $signed(input_fmap_104[7:0]) +
	( 15'sd 14227) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5114) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13076) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1157) * $signed(input_fmap_108[7:0]) +
	( 16'sd 25756) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4704) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18965) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23871) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3811) * $signed(input_fmap_113[7:0]) +
	( 13'sd 2236) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20494) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6095) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23029) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17720) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22664) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21992) * $signed(input_fmap_120[7:0]) +
	( 14'sd 8065) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26792) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18580) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1190) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2477) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3145) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18407) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30018) * $signed(input_fmap_128[7:0]) +
	( 16'sd 26670) * $signed(input_fmap_129[7:0]) +
	( 15'sd 8905) * $signed(input_fmap_130[7:0]) +
	( 16'sd 26944) * $signed(input_fmap_131[7:0]) +
	( 15'sd 15634) * $signed(input_fmap_132[7:0]) +
	( 12'sd 1544) * $signed(input_fmap_133[7:0]) +
	( 14'sd 6856) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18685) * $signed(input_fmap_135[7:0]) +
	( 16'sd 26898) * $signed(input_fmap_136[7:0]) +
	( 16'sd 32314) * $signed(input_fmap_137[7:0]) +
	( 16'sd 25432) * $signed(input_fmap_138[7:0]) +
	( 14'sd 4786) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9203) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5271) * $signed(input_fmap_141[7:0]) +
	( 16'sd 18365) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17338) * $signed(input_fmap_143[7:0]) +
	( 16'sd 25578) * $signed(input_fmap_144[7:0]) +
	( 16'sd 24024) * $signed(input_fmap_145[7:0]) +
	( 16'sd 28006) * $signed(input_fmap_146[7:0]) +
	( 14'sd 6118) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20903) * $signed(input_fmap_148[7:0]) +
	( 16'sd 20047) * $signed(input_fmap_149[7:0]) +
	( 15'sd 13426) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23247) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_152[7:0]) +
	( 15'sd 16224) * $signed(input_fmap_153[7:0]) +
	( 16'sd 26537) * $signed(input_fmap_154[7:0]) +
	( 15'sd 11282) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25681) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14906) * $signed(input_fmap_157[7:0]) +
	( 16'sd 29406) * $signed(input_fmap_158[7:0]) +
	( 15'sd 16068) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22792) * $signed(input_fmap_160[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24597) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27439) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13320) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_165[7:0]) +
	( 16'sd 21669) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26219) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17425) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20397) * $signed(input_fmap_169[7:0]) +
	( 10'sd 438) * $signed(input_fmap_170[7:0]) +
	( 16'sd 21666) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14925) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23226) * $signed(input_fmap_173[7:0]) +
	( 14'sd 5000) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21458) * $signed(input_fmap_175[7:0]) +
	( 15'sd 11976) * $signed(input_fmap_176[7:0]) +
	( 16'sd 21996) * $signed(input_fmap_177[7:0]) +
	( 16'sd 16902) * $signed(input_fmap_178[7:0]) +
	( 16'sd 24427) * $signed(input_fmap_179[7:0]) +
	( 12'sd 1133) * $signed(input_fmap_180[7:0]) +
	( 15'sd 13482) * $signed(input_fmap_181[7:0]) +
	( 15'sd 9849) * $signed(input_fmap_182[7:0]) +
	( 14'sd 7936) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26606) * $signed(input_fmap_184[7:0]) +
	( 16'sd 29697) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6198) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28925) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1491) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25429) * $signed(input_fmap_189[7:0]) +
	( 10'sd 490) * $signed(input_fmap_190[7:0]) +
	( 14'sd 8118) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27290) * $signed(input_fmap_192[7:0]) +
	( 13'sd 2350) * $signed(input_fmap_193[7:0]) +
	( 16'sd 22653) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22673) * $signed(input_fmap_195[7:0]) +
	( 10'sd 345) * $signed(input_fmap_196[7:0]) +
	( 16'sd 20103) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_198[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_199[7:0]) +
	( 16'sd 22185) * $signed(input_fmap_200[7:0]) +
	( 15'sd 16057) * $signed(input_fmap_201[7:0]) +
	( 16'sd 25707) * $signed(input_fmap_202[7:0]) +
	( 16'sd 18185) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11482) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11446) * $signed(input_fmap_205[7:0]) +
	( 14'sd 5733) * $signed(input_fmap_206[7:0]) +
	( 16'sd 27783) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6470) * $signed(input_fmap_208[7:0]) +
	( 16'sd 16681) * $signed(input_fmap_209[7:0]) +
	( 16'sd 22710) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3586) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12988) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28478) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14647) * $signed(input_fmap_214[7:0]) +
	( 16'sd 32261) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1069) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30670) * $signed(input_fmap_217[7:0]) +
	( 15'sd 11803) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15494) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19975) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6606) * $signed(input_fmap_221[7:0]) +
	( 16'sd 31758) * $signed(input_fmap_222[7:0]) +
	( 15'sd 13236) * $signed(input_fmap_223[7:0]) +
	( 15'sd 12159) * $signed(input_fmap_224[7:0]) +
	( 16'sd 16862) * $signed(input_fmap_225[7:0]) +
	( 16'sd 31201) * $signed(input_fmap_226[7:0]) +
	( 16'sd 28971) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8660) * $signed(input_fmap_228[7:0]) +
	( 16'sd 22321) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15828) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18424) * $signed(input_fmap_231[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_232[7:0]) +
	( 14'sd 7667) * $signed(input_fmap_233[7:0]) +
	( 13'sd 3477) * $signed(input_fmap_234[7:0]) +
	( 16'sd 24242) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12348) * $signed(input_fmap_236[7:0]) +
	( 14'sd 5102) * $signed(input_fmap_237[7:0]) +
	( 16'sd 30596) * $signed(input_fmap_238[7:0]) +
	( 16'sd 28845) * $signed(input_fmap_239[7:0]) +
	( 16'sd 16625) * $signed(input_fmap_240[7:0]) +
	( 16'sd 17905) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_243[7:0]) +
	( 15'sd 8794) * $signed(input_fmap_244[7:0]) +
	( 16'sd 17097) * $signed(input_fmap_245[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3389) * $signed(input_fmap_247[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12849) * $signed(input_fmap_250[7:0]) +
	( 15'sd 13208) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3033) * $signed(input_fmap_253[7:0]) +
	( 15'sd 16311) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10407) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_200;
assign conv_mac_200 = 
	( 11'sd 734) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15543) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17232) * $signed(input_fmap_2[7:0]) +
	( 13'sd 2645) * $signed(input_fmap_3[7:0]) +
	( 15'sd 8635) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19051) * $signed(input_fmap_5[7:0]) +
	( 16'sd 26144) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7464) * $signed(input_fmap_7[7:0]) +
	( 16'sd 26511) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15006) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9496) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19687) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2691) * $signed(input_fmap_12[7:0]) +
	( 11'sd 593) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27079) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18828) * $signed(input_fmap_15[7:0]) +
	( 14'sd 4141) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18228) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22534) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30381) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31112) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25222) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2217) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20489) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5271) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23820) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8546) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13091) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24241) * $signed(input_fmap_28[7:0]) +
	( 11'sd 579) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21704) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29988) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1432) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3914) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23972) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28487) * $signed(input_fmap_35[7:0]) +
	( 16'sd 28365) * $signed(input_fmap_36[7:0]) +
	( 16'sd 32393) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30458) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5831) * $signed(input_fmap_39[7:0]) +
	( 15'sd 12180) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28338) * $signed(input_fmap_42[7:0]) +
	( 15'sd 13451) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26176) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31417) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21338) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6196) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21898) * $signed(input_fmap_49[7:0]) +
	( 14'sd 4134) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32186) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27581) * $signed(input_fmap_52[7:0]) +
	( 16'sd 28479) * $signed(input_fmap_53[7:0]) +
	( 13'sd 2051) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28571) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2940) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20652) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3422) * $signed(input_fmap_58[7:0]) +
	( 16'sd 27116) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5292) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13465) * $signed(input_fmap_61[7:0]) +
	( 15'sd 10197) * $signed(input_fmap_62[7:0]) +
	( 16'sd 16579) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31179) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17944) * $signed(input_fmap_65[7:0]) +
	( 15'sd 13386) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8398) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5296) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8832) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12094) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6621) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28741) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21460) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19318) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14134) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8425) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11060) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4892) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14661) * $signed(input_fmap_80[7:0]) +
	( 15'sd 11413) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14977) * $signed(input_fmap_82[7:0]) +
	( 15'sd 10880) * $signed(input_fmap_83[7:0]) +
	( 15'sd 12500) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4137) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14957) * $signed(input_fmap_86[7:0]) +
	( 14'sd 4334) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11318) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30423) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10237) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8430) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_92[7:0]) +
	( 15'sd 13190) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21516) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27771) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18800) * $signed(input_fmap_96[7:0]) +
	( 10'sd 277) * $signed(input_fmap_97[7:0]) +
	( 16'sd 24683) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15433) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31226) * $signed(input_fmap_100[7:0]) +
	( 11'sd 655) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26407) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19221) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11333) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6074) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8329) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23546) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13720) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2938) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2690) * $signed(input_fmap_110[7:0]) +
	( 16'sd 18128) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26900) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19679) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19526) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13488) * $signed(input_fmap_115[7:0]) +
	( 11'sd 789) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4422) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18957) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20330) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17871) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19945) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13462) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20915) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16978) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5241) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19437) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15934) * $signed(input_fmap_127[7:0]) +
	( 16'sd 21369) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10282) * $signed(input_fmap_129[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_130[7:0]) +
	( 15'sd 12550) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18086) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22723) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25901) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23468) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25256) * $signed(input_fmap_136[7:0]) +
	( 16'sd 31186) * $signed(input_fmap_137[7:0]) +
	( 16'sd 24992) * $signed(input_fmap_138[7:0]) +
	( 14'sd 7047) * $signed(input_fmap_139[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29477) * $signed(input_fmap_141[7:0]) +
	( 16'sd 16520) * $signed(input_fmap_142[7:0]) +
	( 16'sd 24008) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28633) * $signed(input_fmap_144[7:0]) +
	( 16'sd 24496) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27790) * $signed(input_fmap_146[7:0]) +
	( 14'sd 7656) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4137) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15474) * $signed(input_fmap_149[7:0]) +
	( 15'sd 10732) * $signed(input_fmap_150[7:0]) +
	( 16'sd 25254) * $signed(input_fmap_151[7:0]) +
	( 15'sd 13475) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24626) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30154) * $signed(input_fmap_154[7:0]) +
	( 16'sd 32136) * $signed(input_fmap_155[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_156[7:0]) +
	( 15'sd 14192) * $signed(input_fmap_157[7:0]) +
	( 14'sd 7185) * $signed(input_fmap_158[7:0]) +
	( 16'sd 28013) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5757) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1981) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14414) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2292) * $signed(input_fmap_163[7:0]) +
	( 16'sd 31002) * $signed(input_fmap_164[7:0]) +
	( 14'sd 4421) * $signed(input_fmap_165[7:0]) +
	( 14'sd 5035) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31826) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26385) * $signed(input_fmap_168[7:0]) +
	( 16'sd 24639) * $signed(input_fmap_169[7:0]) +
	( 16'sd 19168) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7608) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1971) * $signed(input_fmap_172[7:0]) +
	( 16'sd 25412) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26441) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15328) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13276) * $signed(input_fmap_176[7:0]) +
	( 12'sd 1117) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3674) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15351) * $signed(input_fmap_180[7:0]) +
	( 15'sd 13008) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4258) * $signed(input_fmap_182[7:0]) +
	( 16'sd 22314) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9771) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11396) * $signed(input_fmap_185[7:0]) +
	( 15'sd 11707) * $signed(input_fmap_186[7:0]) +
	( 16'sd 17424) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23784) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26155) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5664) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14816) * $signed(input_fmap_191[7:0]) +
	( 14'sd 5391) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15136) * $signed(input_fmap_193[7:0]) +
	( 14'sd 5409) * $signed(input_fmap_194[7:0]) +
	( 16'sd 31624) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22415) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5775) * $signed(input_fmap_197[7:0]) +
	( 15'sd 11257) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24746) * $signed(input_fmap_199[7:0]) +
	( 16'sd 31886) * $signed(input_fmap_200[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_202[7:0]) +
	( 16'sd 29986) * $signed(input_fmap_203[7:0]) +
	( 16'sd 29641) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11117) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28775) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3025) * $signed(input_fmap_207[7:0]) +
	( 13'sd 2310) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13569) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1215) * $signed(input_fmap_210[7:0]) +
	( 11'sd 912) * $signed(input_fmap_211[7:0]) +
	( 15'sd 10706) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11098) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17648) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2386) * $signed(input_fmap_215[7:0]) +
	( 16'sd 21862) * $signed(input_fmap_216[7:0]) +
	( 16'sd 22839) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28268) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14781) * $signed(input_fmap_219[7:0]) +
	( 16'sd 32434) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1758) * $signed(input_fmap_221[7:0]) +
	( 14'sd 8018) * $signed(input_fmap_222[7:0]) +
	( 16'sd 29823) * $signed(input_fmap_223[7:0]) +
	( 13'sd 3495) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27930) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7121) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6155) * $signed(input_fmap_227[7:0]) +
	( 14'sd 5352) * $signed(input_fmap_228[7:0]) +
	( 11'sd 1009) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28791) * $signed(input_fmap_230[7:0]) +
	( 13'sd 2390) * $signed(input_fmap_231[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15308) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18254) * $signed(input_fmap_234[7:0]) +
	( 16'sd 28497) * $signed(input_fmap_235[7:0]) +
	( 14'sd 6772) * $signed(input_fmap_236[7:0]) +
	( 15'sd 13057) * $signed(input_fmap_237[7:0]) +
	( 16'sd 31386) * $signed(input_fmap_238[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18131) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15845) * $signed(input_fmap_241[7:0]) +
	( 15'sd 12053) * $signed(input_fmap_242[7:0]) +
	( 15'sd 10541) * $signed(input_fmap_243[7:0]) +
	( 13'sd 2536) * $signed(input_fmap_244[7:0]) +
	( 13'sd 3553) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30023) * $signed(input_fmap_246[7:0]) +
	( 16'sd 19387) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10603) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25422) * $signed(input_fmap_249[7:0]) +
	( 15'sd 11891) * $signed(input_fmap_250[7:0]) +
	( 16'sd 25918) * $signed(input_fmap_251[7:0]) +
	( 13'sd 3567) * $signed(input_fmap_252[7:0]) +
	( 13'sd 3445) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9441) * $signed(input_fmap_254[7:0]) +
	( 15'sd 9967) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_201;
assign conv_mac_201 = 
	( 16'sd 18795) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18117) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7446) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17665) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19682) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25998) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31432) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18055) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19723) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2318) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4722) * $signed(input_fmap_10[7:0]) +
	( 14'sd 4474) * $signed(input_fmap_11[7:0]) +
	( 16'sd 32454) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_14[7:0]) +
	( 16'sd 30638) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28422) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22567) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8528) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28219) * $signed(input_fmap_19[7:0]) +
	( 15'sd 13816) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3988) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4522) * $signed(input_fmap_22[7:0]) +
	( 16'sd 20324) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4130) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14256) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15340) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31665) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13787) * $signed(input_fmap_28[7:0]) +
	( 15'sd 8874) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29517) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32041) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29800) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2058) * $signed(input_fmap_33[7:0]) +
	( 14'sd 4379) * $signed(input_fmap_34[7:0]) +
	( 15'sd 16252) * $signed(input_fmap_35[7:0]) +
	( 16'sd 26856) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22525) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7621) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13837) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18422) * $signed(input_fmap_40[7:0]) +
	( 15'sd 14354) * $signed(input_fmap_41[7:0]) +
	( 16'sd 29559) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3953) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21607) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29795) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15658) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17904) * $signed(input_fmap_47[7:0]) +
	( 14'sd 8074) * $signed(input_fmap_48[7:0]) +
	( 11'sd 980) * $signed(input_fmap_49[7:0]) +
	( 16'sd 28061) * $signed(input_fmap_50[7:0]) +
	( 16'sd 28607) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25470) * $signed(input_fmap_52[7:0]) +
	( 16'sd 19668) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10745) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9786) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21044) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7818) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1091) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26689) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30484) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28268) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17190) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2222) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18282) * $signed(input_fmap_64[7:0]) +
	( 16'sd 18620) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3603) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11608) * $signed(input_fmap_67[7:0]) +
	( 16'sd 30839) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31078) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11037) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18113) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3891) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1029) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6822) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17681) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29041) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30024) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2726) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1897) * $signed(input_fmap_79[7:0]) +
	( 16'sd 32661) * $signed(input_fmap_80[7:0]) +
	( 15'sd 9906) * $signed(input_fmap_81[7:0]) +
	( 16'sd 25075) * $signed(input_fmap_82[7:0]) +
	( 15'sd 11764) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28330) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17162) * $signed(input_fmap_86[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_87[7:0]) +
	( 11'sd 959) * $signed(input_fmap_88[7:0]) +
	( 13'sd 3105) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22196) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11284) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12019) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3994) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30952) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28737) * $signed(input_fmap_95[7:0]) +
	( 13'sd 4036) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7257) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26227) * $signed(input_fmap_98[7:0]) +
	( 12'sd 2015) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5255) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29212) * $signed(input_fmap_101[7:0]) +
	( 11'sd 718) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19670) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17315) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31016) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4291) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27308) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28375) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13203) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21441) * $signed(input_fmap_110[7:0]) +
	( 16'sd 16989) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19900) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31440) * $signed(input_fmap_113[7:0]) +
	( 10'sd 339) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12485) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22821) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4372) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29488) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5480) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15298) * $signed(input_fmap_122[7:0]) +
	( 14'sd 8043) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11437) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27552) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17431) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6264) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13839) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5772) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30205) * $signed(input_fmap_130[7:0]) +
	( 16'sd 22245) * $signed(input_fmap_131[7:0]) +
	( 15'sd 13903) * $signed(input_fmap_132[7:0]) +
	( 14'sd 4988) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2657) * $signed(input_fmap_134[7:0]) +
	( 14'sd 4866) * $signed(input_fmap_135[7:0]) +
	( 15'sd 11253) * $signed(input_fmap_136[7:0]) +
	( 15'sd 8680) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29162) * $signed(input_fmap_138[7:0]) +
	( 16'sd 26027) * $signed(input_fmap_139[7:0]) +
	( 16'sd 18278) * $signed(input_fmap_140[7:0]) +
	( 13'sd 4078) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28042) * $signed(input_fmap_142[7:0]) +
	( 15'sd 9692) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_144[7:0]) +
	( 12'sd 1495) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1356) * $signed(input_fmap_146[7:0]) +
	( 15'sd 15744) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28140) * $signed(input_fmap_148[7:0]) +
	( 16'sd 20278) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18746) * $signed(input_fmap_150[7:0]) +
	( 16'sd 16943) * $signed(input_fmap_151[7:0]) +
	( 15'sd 11109) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23849) * $signed(input_fmap_153[7:0]) +
	( 16'sd 19142) * $signed(input_fmap_154[7:0]) +
	( 9'sd 180) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24150) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18264) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25104) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5459) * $signed(input_fmap_159[7:0]) +
	( 16'sd 16945) * $signed(input_fmap_160[7:0]) +
	( 15'sd 10196) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24816) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30995) * $signed(input_fmap_163[7:0]) +
	( 16'sd 18221) * $signed(input_fmap_164[7:0]) +
	( 16'sd 29118) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18839) * $signed(input_fmap_166[7:0]) +
	( 16'sd 16566) * $signed(input_fmap_167[7:0]) +
	( 15'sd 16382) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11731) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17493) * $signed(input_fmap_170[7:0]) +
	( 12'sd 1285) * $signed(input_fmap_171[7:0]) +
	( 16'sd 28269) * $signed(input_fmap_172[7:0]) +
	( 15'sd 14238) * $signed(input_fmap_173[7:0]) +
	( 16'sd 31535) * $signed(input_fmap_174[7:0]) +
	( 15'sd 11512) * $signed(input_fmap_175[7:0]) +
	( 16'sd 16466) * $signed(input_fmap_176[7:0]) +
	( 15'sd 9175) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32730) * $signed(input_fmap_178[7:0]) +
	( 15'sd 9039) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_180[7:0]) +
	( 16'sd 27018) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10462) * $signed(input_fmap_182[7:0]) +
	( 12'sd 1171) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9711) * $signed(input_fmap_184[7:0]) +
	( 15'sd 14514) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9220) * $signed(input_fmap_186[7:0]) +
	( 16'sd 23485) * $signed(input_fmap_187[7:0]) +
	( 16'sd 18266) * $signed(input_fmap_188[7:0]) +
	( 11'sd 653) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17000) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20802) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31785) * $signed(input_fmap_192[7:0]) +
	( 16'sd 17974) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12148) * $signed(input_fmap_194[7:0]) +
	( 15'sd 9424) * $signed(input_fmap_195[7:0]) +
	( 16'sd 21370) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25880) * $signed(input_fmap_197[7:0]) +
	( 11'sd 553) * $signed(input_fmap_198[7:0]) +
	( 16'sd 29406) * $signed(input_fmap_199[7:0]) +
	( 14'sd 7174) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22774) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11390) * $signed(input_fmap_202[7:0]) +
	( 13'sd 3256) * $signed(input_fmap_203[7:0]) +
	( 16'sd 26444) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2526) * $signed(input_fmap_206[7:0]) +
	( 15'sd 10871) * $signed(input_fmap_207[7:0]) +
	( 15'sd 13261) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13154) * $signed(input_fmap_209[7:0]) +
	( 16'sd 32433) * $signed(input_fmap_210[7:0]) +
	( 16'sd 18454) * $signed(input_fmap_211[7:0]) +
	( 10'sd 454) * $signed(input_fmap_212[7:0]) +
	( 16'sd 25407) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28206) * $signed(input_fmap_214[7:0]) +
	( 16'sd 28439) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11099) * $signed(input_fmap_216[7:0]) +
	( 15'sd 14925) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10613) * $signed(input_fmap_218[7:0]) +
	( 16'sd 23223) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21615) * $signed(input_fmap_220[7:0]) +
	( 16'sd 30190) * $signed(input_fmap_221[7:0]) +
	( 9'sd 128) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28353) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14760) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15523) * $signed(input_fmap_225[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6033) * $signed(input_fmap_227[7:0]) +
	( 16'sd 32634) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23426) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14130) * $signed(input_fmap_230[7:0]) +
	( 13'sd 2415) * $signed(input_fmap_231[7:0]) +
	( 14'sd 4607) * $signed(input_fmap_232[7:0]) +
	( 16'sd 20775) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18392) * $signed(input_fmap_234[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30623) * $signed(input_fmap_236[7:0]) +
	( 16'sd 32291) * $signed(input_fmap_237[7:0]) +
	( 15'sd 8569) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26518) * $signed(input_fmap_239[7:0]) +
	( 14'sd 6786) * $signed(input_fmap_240[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_241[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_242[7:0]) +
	( 14'sd 5564) * $signed(input_fmap_243[7:0]) +
	( 9'sd 215) * $signed(input_fmap_244[7:0]) +
	( 15'sd 15749) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15941) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13901) * $signed(input_fmap_247[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_248[7:0]) +
	( 16'sd 27268) * $signed(input_fmap_249[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_250[7:0]) +
	( 15'sd 8845) * $signed(input_fmap_251[7:0]) +
	( 15'sd 12500) * $signed(input_fmap_252[7:0]) +
	( 16'sd 23227) * $signed(input_fmap_253[7:0]) +
	( 16'sd 28709) * $signed(input_fmap_254[7:0]) +
	( 15'sd 15813) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_202;
assign conv_mac_202 = 
	( 16'sd 27674) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15104) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21197) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14405) * $signed(input_fmap_3[7:0]) +
	( 16'sd 29477) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8798) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9080) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3383) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11032) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25290) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10621) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10164) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28684) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14330) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10914) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3353) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8928) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27786) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23952) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27307) * $signed(input_fmap_20[7:0]) +
	( 16'sd 16676) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14238) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2179) * $signed(input_fmap_23[7:0]) +
	( 15'sd 9243) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3617) * $signed(input_fmap_25[7:0]) +
	( 16'sd 30002) * $signed(input_fmap_26[7:0]) +
	( 14'sd 8007) * $signed(input_fmap_27[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21692) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28679) * $signed(input_fmap_31[7:0]) +
	( 13'sd 3812) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2237) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26000) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3650) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12341) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30444) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1217) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9620) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2351) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4738) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_42[7:0]) +
	( 16'sd 16659) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15123) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20423) * $signed(input_fmap_45[7:0]) +
	( 16'sd 26750) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9901) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9240) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_49[7:0]) +
	( 16'sd 18444) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12799) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11443) * $signed(input_fmap_52[7:0]) +
	( 14'sd 8105) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18515) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24583) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4131) * $signed(input_fmap_56[7:0]) +
	( 16'sd 19978) * $signed(input_fmap_57[7:0]) +
	( 12'sd 1757) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22468) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29356) * $signed(input_fmap_60[7:0]) +
	( 15'sd 8944) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23263) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23140) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15990) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12337) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10215) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17877) * $signed(input_fmap_67[7:0]) +
	( 9'sd 243) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4190) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5659) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19367) * $signed(input_fmap_71[7:0]) +
	( 15'sd 10251) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27402) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32219) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15415) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12500) * $signed(input_fmap_76[7:0]) +
	( 15'sd 8958) * $signed(input_fmap_77[7:0]) +
	( 15'sd 16009) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21601) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5095) * $signed(input_fmap_80[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1247) * $signed(input_fmap_82[7:0]) +
	( 11'sd 793) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6882) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32567) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14168) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30420) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25652) * $signed(input_fmap_89[7:0]) +
	( 16'sd 21783) * $signed(input_fmap_90[7:0]) +
	( 13'sd 3753) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15373) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3694) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18663) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19339) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4111) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28498) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15479) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26357) * $signed(input_fmap_99[7:0]) +
	( 10'sd 268) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12917) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23607) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10527) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7100) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23612) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6675) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25281) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28615) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_110[7:0]) +
	( 15'sd 16281) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13805) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_113[7:0]) +
	( 15'sd 13786) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24148) * $signed(input_fmap_115[7:0]) +
	( 15'sd 8922) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20754) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_118[7:0]) +
	( 16'sd 26122) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29002) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9464) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24792) * $signed(input_fmap_122[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31418) * $signed(input_fmap_124[7:0]) +
	( 14'sd 5380) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15817) * $signed(input_fmap_126[7:0]) +
	( 16'sd 23305) * $signed(input_fmap_127[7:0]) +
	( 16'sd 30866) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10807) * $signed(input_fmap_129[7:0]) +
	( 16'sd 17100) * $signed(input_fmap_130[7:0]) +
	( 16'sd 22255) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8236) * $signed(input_fmap_132[7:0]) +
	( 15'sd 8639) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1223) * $signed(input_fmap_134[7:0]) +
	( 13'sd 3434) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7261) * $signed(input_fmap_136[7:0]) +
	( 14'sd 5059) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10243) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27579) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3011) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18391) * $signed(input_fmap_141[7:0]) +
	( 16'sd 20094) * $signed(input_fmap_142[7:0]) +
	( 15'sd 13172) * $signed(input_fmap_143[7:0]) +
	( 16'sd 32411) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28009) * $signed(input_fmap_145[7:0]) +
	( 15'sd 8442) * $signed(input_fmap_146[7:0]) +
	( 12'sd 1446) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11278) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17415) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18587) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14940) * $signed(input_fmap_151[7:0]) +
	( 16'sd 22482) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12000) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31551) * $signed(input_fmap_154[7:0]) +
	( 16'sd 16456) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15257) * $signed(input_fmap_156[7:0]) +
	( 15'sd 12561) * $signed(input_fmap_157[7:0]) +
	( 13'sd 3803) * $signed(input_fmap_158[7:0]) +
	( 8'sd 82) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18061) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28191) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29140) * $signed(input_fmap_162[7:0]) +
	( 15'sd 9874) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10324) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_165[7:0]) +
	( 16'sd 29294) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23534) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1803) * $signed(input_fmap_168[7:0]) +
	( 12'sd 1188) * $signed(input_fmap_169[7:0]) +
	( 16'sd 29644) * $signed(input_fmap_170[7:0]) +
	( 16'sd 28470) * $signed(input_fmap_171[7:0]) +
	( 16'sd 17527) * $signed(input_fmap_172[7:0]) +
	( 15'sd 13379) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16524) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21331) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29742) * $signed(input_fmap_177[7:0]) +
	( 16'sd 23198) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3593) * $signed(input_fmap_179[7:0]) +
	( 16'sd 22281) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15878) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6512) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12292) * $signed(input_fmap_183[7:0]) +
	( 16'sd 23462) * $signed(input_fmap_184[7:0]) +
	( 16'sd 19247) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26113) * $signed(input_fmap_186[7:0]) +
	( 15'sd 13207) * $signed(input_fmap_187[7:0]) +
	( 15'sd 14765) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5862) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4303) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19562) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15952) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27223) * $signed(input_fmap_193[7:0]) +
	( 15'sd 16061) * $signed(input_fmap_194[7:0]) +
	( 14'sd 6699) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24136) * $signed(input_fmap_196[7:0]) +
	( 15'sd 11587) * $signed(input_fmap_197[7:0]) +
	( 12'sd 1558) * $signed(input_fmap_198[7:0]) +
	( 16'sd 20840) * $signed(input_fmap_199[7:0]) +
	( 15'sd 8812) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18678) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31642) * $signed(input_fmap_202[7:0]) +
	( 15'sd 11627) * $signed(input_fmap_203[7:0]) +
	( 16'sd 21044) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29849) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27589) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11713) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7780) * $signed(input_fmap_209[7:0]) +
	( 14'sd 6057) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15896) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29092) * $signed(input_fmap_213[7:0]) +
	( 16'sd 29789) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7698) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28218) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25471) * $signed(input_fmap_217[7:0]) +
	( 11'sd 546) * $signed(input_fmap_218[7:0]) +
	( 16'sd 24044) * $signed(input_fmap_219[7:0]) +
	( 15'sd 8336) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27322) * $signed(input_fmap_221[7:0]) +
	( 16'sd 31727) * $signed(input_fmap_222[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_223[7:0]) +
	( 16'sd 21240) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3040) * $signed(input_fmap_225[7:0]) +
	( 13'sd 2575) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3303) * $signed(input_fmap_227[7:0]) +
	( 16'sd 28372) * $signed(input_fmap_228[7:0]) +
	( 12'sd 1504) * $signed(input_fmap_229[7:0]) +
	( 13'sd 2753) * $signed(input_fmap_230[7:0]) +
	( 13'sd 2838) * $signed(input_fmap_231[7:0]) +
	( 16'sd 25970) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10017) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19744) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3927) * $signed(input_fmap_235[7:0]) +
	( 16'sd 21707) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11093) * $signed(input_fmap_237[7:0]) +
	( 16'sd 24576) * $signed(input_fmap_238[7:0]) +
	( 16'sd 28963) * $signed(input_fmap_239[7:0]) +
	( 16'sd 24267) * $signed(input_fmap_240[7:0]) +
	( 15'sd 11847) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1062) * $signed(input_fmap_242[7:0]) +
	( 16'sd 18903) * $signed(input_fmap_243[7:0]) +
	( 15'sd 11559) * $signed(input_fmap_244[7:0]) +
	( 14'sd 6990) * $signed(input_fmap_245[7:0]) +
	( 15'sd 8283) * $signed(input_fmap_246[7:0]) +
	( 12'sd 1695) * $signed(input_fmap_247[7:0]) +
	( 11'sd 682) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2976) * $signed(input_fmap_249[7:0]) +
	( 16'sd 19724) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21176) * $signed(input_fmap_251[7:0]) +
	( 16'sd 31295) * $signed(input_fmap_252[7:0]) +
	( 16'sd 22212) * $signed(input_fmap_253[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26922) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_203;
assign conv_mac_203 = 
	( 14'sd 7298) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11416) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7707) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7266) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17927) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10264) * $signed(input_fmap_5[7:0]) +
	( 13'sd 2314) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28217) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18609) * $signed(input_fmap_8[7:0]) +
	( 13'sd 2335) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26814) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20024) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1224) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9218) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1377) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1782) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19475) * $signed(input_fmap_16[7:0]) +
	( 10'sd 305) * $signed(input_fmap_17[7:0]) +
	( 16'sd 22856) * $signed(input_fmap_18[7:0]) +
	( 16'sd 20932) * $signed(input_fmap_19[7:0]) +
	( 15'sd 15819) * $signed(input_fmap_20[7:0]) +
	( 16'sd 30670) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20129) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12220) * $signed(input_fmap_23[7:0]) +
	( 7'sd 32) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24062) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5515) * $signed(input_fmap_26[7:0]) +
	( 14'sd 4671) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13692) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3304) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12572) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27868) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9475) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27399) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24371) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15929) * $signed(input_fmap_35[7:0]) +
	( 16'sd 27809) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9720) * $signed(input_fmap_37[7:0]) +
	( 16'sd 20152) * $signed(input_fmap_38[7:0]) +
	( 16'sd 16950) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_40[7:0]) +
	( 16'sd 16519) * $signed(input_fmap_41[7:0]) +
	( 16'sd 24023) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25642) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11696) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28227) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9254) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27633) * $signed(input_fmap_47[7:0]) +
	( 16'sd 18961) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27655) * $signed(input_fmap_49[7:0]) +
	( 12'sd 1549) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26221) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6260) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30504) * $signed(input_fmap_53[7:0]) +
	( 14'sd 7561) * $signed(input_fmap_54[7:0]) +
	( 16'sd 16771) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18134) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20850) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31896) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28394) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19340) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16704) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29467) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2604) * $signed(input_fmap_63[7:0]) +
	( 16'sd 31434) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22652) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27510) * $signed(input_fmap_66[7:0]) +
	( 10'sd 278) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27524) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20679) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19752) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24869) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28380) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21430) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11460) * $signed(input_fmap_74[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_75[7:0]) +
	( 16'sd 22234) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13347) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13915) * $signed(input_fmap_78[7:0]) +
	( 12'sd 1444) * $signed(input_fmap_79[7:0]) +
	( 13'sd 4069) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25594) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9130) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5039) * $signed(input_fmap_83[7:0]) +
	( 16'sd 27550) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14615) * $signed(input_fmap_85[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5365) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28283) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7808) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12983) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28290) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30071) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3305) * $signed(input_fmap_93[7:0]) +
	( 14'sd 4531) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8027) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5413) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28152) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22290) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28057) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17667) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15376) * $signed(input_fmap_101[7:0]) +
	( 15'sd 13902) * $signed(input_fmap_102[7:0]) +
	( 16'sd 28048) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7219) * $signed(input_fmap_104[7:0]) +
	( 16'sd 20451) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28511) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11162) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19671) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19323) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23788) * $signed(input_fmap_111[7:0]) +
	( 16'sd 25619) * $signed(input_fmap_112[7:0]) +
	( 13'sd 3414) * $signed(input_fmap_113[7:0]) +
	( 14'sd 7999) * $signed(input_fmap_114[7:0]) +
	( 16'sd 16451) * $signed(input_fmap_115[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23469) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15363) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2696) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23128) * $signed(input_fmap_120[7:0]) +
	( 16'sd 28513) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12743) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15012) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11920) * $signed(input_fmap_124[7:0]) +
	( 16'sd 19403) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13680) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13904) * $signed(input_fmap_127[7:0]) +
	( 16'sd 27236) * $signed(input_fmap_128[7:0]) +
	( 16'sd 30632) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6842) * $signed(input_fmap_130[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14128) * $signed(input_fmap_132[7:0]) +
	( 15'sd 15243) * $signed(input_fmap_133[7:0]) +
	( 15'sd 8834) * $signed(input_fmap_134[7:0]) +
	( 16'sd 25476) * $signed(input_fmap_135[7:0]) +
	( 16'sd 16497) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12513) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28618) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30766) * $signed(input_fmap_140[7:0]) +
	( 14'sd 7189) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11168) * $signed(input_fmap_142[7:0]) +
	( 15'sd 15251) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31991) * $signed(input_fmap_144[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_145[7:0]) +
	( 16'sd 32607) * $signed(input_fmap_146[7:0]) +
	( 15'sd 15705) * $signed(input_fmap_147[7:0]) +
	( 13'sd 4094) * $signed(input_fmap_148[7:0]) +
	( 15'sd 9117) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18319) * $signed(input_fmap_150[7:0]) +
	( 16'sd 16554) * $signed(input_fmap_151[7:0]) +
	( 16'sd 28088) * $signed(input_fmap_152[7:0]) +
	( 16'sd 26101) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4101) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5201) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14454) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31100) * $signed(input_fmap_157[7:0]) +
	( 14'sd 6402) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6629) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4184) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29326) * $signed(input_fmap_162[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_163[7:0]) +
	( 16'sd 17858) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22938) * $signed(input_fmap_165[7:0]) +
	( 15'sd 13359) * $signed(input_fmap_166[7:0]) +
	( 15'sd 10882) * $signed(input_fmap_167[7:0]) +
	( 16'sd 27708) * $signed(input_fmap_168[7:0]) +
	( 16'sd 31001) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2561) * $signed(input_fmap_170[7:0]) +
	( 15'sd 9073) * $signed(input_fmap_171[7:0]) +
	( 15'sd 14657) * $signed(input_fmap_172[7:0]) +
	( 14'sd 7060) * $signed(input_fmap_173[7:0]) +
	( 16'sd 31766) * $signed(input_fmap_174[7:0]) +
	( 16'sd 20902) * $signed(input_fmap_175[7:0]) +
	( 14'sd 6779) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22036) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15013) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28252) * $signed(input_fmap_179[7:0]) +
	( 16'sd 26875) * $signed(input_fmap_180[7:0]) +
	( 15'sd 8232) * $signed(input_fmap_181[7:0]) +
	( 16'sd 25540) * $signed(input_fmap_182[7:0]) +
	( 16'sd 26774) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30726) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_185[7:0]) +
	( 14'sd 7392) * $signed(input_fmap_186[7:0]) +
	( 16'sd 23898) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12785) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30776) * $signed(input_fmap_189[7:0]) +
	( 15'sd 11479) * $signed(input_fmap_190[7:0]) +
	( 15'sd 11853) * $signed(input_fmap_191[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29134) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29389) * $signed(input_fmap_194[7:0]) +
	( 16'sd 16723) * $signed(input_fmap_195[7:0]) +
	( 16'sd 31870) * $signed(input_fmap_196[7:0]) +
	( 16'sd 30947) * $signed(input_fmap_197[7:0]) +
	( 15'sd 12026) * $signed(input_fmap_198[7:0]) +
	( 13'sd 3656) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20094) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9377) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17743) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2902) * $signed(input_fmap_203[7:0]) +
	( 16'sd 22085) * $signed(input_fmap_204[7:0]) +
	( 13'sd 3078) * $signed(input_fmap_205[7:0]) +
	( 7'sd 42) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12332) * $signed(input_fmap_207[7:0]) +
	( 16'sd 26060) * $signed(input_fmap_208[7:0]) +
	( 14'sd 6747) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1943) * $signed(input_fmap_210[7:0]) +
	( 16'sd 32348) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24443) * $signed(input_fmap_212[7:0]) +
	( 15'sd 9758) * $signed(input_fmap_213[7:0]) +
	( 16'sd 17642) * $signed(input_fmap_214[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_215[7:0]) +
	( 16'sd 22179) * $signed(input_fmap_216[7:0]) +
	( 11'sd 616) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_218[7:0]) +
	( 15'sd 11182) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_220[7:0]) +
	( 16'sd 17566) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18906) * $signed(input_fmap_222[7:0]) +
	( 16'sd 30129) * $signed(input_fmap_223[7:0]) +
	( 16'sd 16915) * $signed(input_fmap_224[7:0]) +
	( 16'sd 27026) * $signed(input_fmap_225[7:0]) +
	( 16'sd 32185) * $signed(input_fmap_226[7:0]) +
	( 16'sd 16733) * $signed(input_fmap_227[7:0]) +
	( 14'sd 6286) * $signed(input_fmap_228[7:0]) +
	( 16'sd 19266) * $signed(input_fmap_229[7:0]) +
	( 16'sd 16393) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20429) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14097) * $signed(input_fmap_232[7:0]) +
	( 16'sd 20866) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19920) * $signed(input_fmap_234[7:0]) +
	( 16'sd 16396) * $signed(input_fmap_235[7:0]) +
	( 14'sd 5246) * $signed(input_fmap_236[7:0]) +
	( 11'sd 581) * $signed(input_fmap_237[7:0]) +
	( 14'sd 4137) * $signed(input_fmap_238[7:0]) +
	( 15'sd 8865) * $signed(input_fmap_239[7:0]) +
	( 16'sd 27467) * $signed(input_fmap_240[7:0]) +
	( 16'sd 23041) * $signed(input_fmap_241[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13428) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19848) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30358) * $signed(input_fmap_245[7:0]) +
	( 16'sd 31007) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11832) * $signed(input_fmap_247[7:0]) +
	( 15'sd 10517) * $signed(input_fmap_248[7:0]) +
	( 16'sd 19955) * $signed(input_fmap_249[7:0]) +
	( 15'sd 8193) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7971) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13684) * $signed(input_fmap_252[7:0]) +
	( 16'sd 30568) * $signed(input_fmap_253[7:0]) +
	( 16'sd 24548) * $signed(input_fmap_254[7:0]) +
	( 16'sd 22546) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_204;
assign conv_mac_204 = 
	( 13'sd 2223) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5368) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31445) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24279) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25819) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20937) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25011) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9444) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11204) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25025) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6370) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3152) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24411) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15140) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31357) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32471) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17555) * $signed(input_fmap_17[7:0]) +
	( 15'sd 12486) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30698) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19772) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6652) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9267) * $signed(input_fmap_22[7:0]) +
	( 16'sd 25408) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8388) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21468) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15385) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28550) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6612) * $signed(input_fmap_28[7:0]) +
	( 16'sd 24330) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27443) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32565) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5824) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22777) * $signed(input_fmap_33[7:0]) +
	( 9'sd 229) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10326) * $signed(input_fmap_35[7:0]) +
	( 13'sd 2891) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18720) * $signed(input_fmap_37[7:0]) +
	( 12'sd 1635) * $signed(input_fmap_38[7:0]) +
	( 15'sd 15491) * $signed(input_fmap_39[7:0]) +
	( 15'sd 15963) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18872) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32323) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32399) * $signed(input_fmap_43[7:0]) +
	( 14'sd 7295) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21390) * $signed(input_fmap_45[7:0]) +
	( 16'sd 28204) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13212) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30323) * $signed(input_fmap_48[7:0]) +
	( 14'sd 7944) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29392) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19927) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19833) * $signed(input_fmap_52[7:0]) +
	( 16'sd 23619) * $signed(input_fmap_53[7:0]) +
	( 16'sd 19317) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5024) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4270) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14103) * $signed(input_fmap_57[7:0]) +
	( 16'sd 23971) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19425) * $signed(input_fmap_60[7:0]) +
	( 15'sd 9476) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11524) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3828) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15637) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31044) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23483) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8515) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5513) * $signed(input_fmap_68[7:0]) +
	( 16'sd 24005) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27990) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16537) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5074) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19009) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7065) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22451) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4793) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23956) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17531) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22047) * $signed(input_fmap_79[7:0]) +
	( 14'sd 6234) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13131) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24734) * $signed(input_fmap_82[7:0]) +
	( 15'sd 15876) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21072) * $signed(input_fmap_84[7:0]) +
	( 16'sd 30856) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22991) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8598) * $signed(input_fmap_87[7:0]) +
	( 16'sd 30252) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13277) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31389) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5426) * $signed(input_fmap_91[7:0]) +
	( 15'sd 12041) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22409) * $signed(input_fmap_93[7:0]) +
	( 16'sd 31320) * $signed(input_fmap_94[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24913) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7078) * $signed(input_fmap_97[7:0]) +
	( 16'sd 25367) * $signed(input_fmap_98[7:0]) +
	( 16'sd 16814) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16583) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28318) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18834) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13448) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23177) * $signed(input_fmap_104[7:0]) +
	( 14'sd 7879) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22824) * $signed(input_fmap_106[7:0]) +
	( 15'sd 12911) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14875) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23232) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31420) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3321) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26173) * $signed(input_fmap_112[7:0]) +
	( 16'sd 21575) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5068) * $signed(input_fmap_114[7:0]) +
	( 10'sd 264) * $signed(input_fmap_115[7:0]) +
	( 15'sd 16307) * $signed(input_fmap_116[7:0]) +
	( 14'sd 5521) * $signed(input_fmap_117[7:0]) +
	( 15'sd 15707) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30621) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12820) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3349) * $signed(input_fmap_121[7:0]) +
	( 14'sd 7630) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28467) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13065) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14236) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11860) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9453) * $signed(input_fmap_127[7:0]) +
	( 15'sd 14096) * $signed(input_fmap_128[7:0]) +
	( 16'sd 21769) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10934) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24896) * $signed(input_fmap_131[7:0]) +
	( 16'sd 31429) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31513) * $signed(input_fmap_133[7:0]) +
	( 15'sd 16315) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31515) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31828) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12624) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19154) * $signed(input_fmap_138[7:0]) +
	( 14'sd 4197) * $signed(input_fmap_139[7:0]) +
	( 13'sd 2299) * $signed(input_fmap_140[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_142[7:0]) +
	( 14'sd 4239) * $signed(input_fmap_143[7:0]) +
	( 14'sd 7010) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23204) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19543) * $signed(input_fmap_146[7:0]) +
	( 15'sd 10369) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23853) * $signed(input_fmap_149[7:0]) +
	( 15'sd 16153) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3868) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31948) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12993) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30445) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17161) * $signed(input_fmap_156[7:0]) +
	( 16'sd 32145) * $signed(input_fmap_157[7:0]) +
	( 16'sd 23177) * $signed(input_fmap_158[7:0]) +
	( 16'sd 22886) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11224) * $signed(input_fmap_160[7:0]) +
	( 13'sd 4039) * $signed(input_fmap_161[7:0]) +
	( 16'sd 31028) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8198) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25542) * $signed(input_fmap_164[7:0]) +
	( 16'sd 16911) * $signed(input_fmap_165[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17691) * $signed(input_fmap_167[7:0]) +
	( 16'sd 32020) * $signed(input_fmap_168[7:0]) +
	( 14'sd 6412) * $signed(input_fmap_169[7:0]) +
	( 10'sd 436) * $signed(input_fmap_170[7:0]) +
	( 14'sd 8120) * $signed(input_fmap_171[7:0]) +
	( 13'sd 2977) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12645) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11151) * $signed(input_fmap_174[7:0]) +
	( 16'sd 26666) * $signed(input_fmap_175[7:0]) +
	( 16'sd 23348) * $signed(input_fmap_176[7:0]) +
	( 16'sd 26515) * $signed(input_fmap_177[7:0]) +
	( 16'sd 16720) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20311) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6380) * $signed(input_fmap_180[7:0]) +
	( 16'sd 16842) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30012) * $signed(input_fmap_182[7:0]) +
	( 16'sd 21838) * $signed(input_fmap_183[7:0]) +
	( 16'sd 18003) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7391) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26904) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27199) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21856) * $signed(input_fmap_188[7:0]) +
	( 8'sd 82) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20515) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32643) * $signed(input_fmap_191[7:0]) +
	( 12'sd 1864) * $signed(input_fmap_192[7:0]) +
	( 15'sd 13919) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29653) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29309) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14402) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21101) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24257) * $signed(input_fmap_199[7:0]) +
	( 12'sd 1036) * $signed(input_fmap_200[7:0]) +
	( 14'sd 5574) * $signed(input_fmap_201[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_202[7:0]) +
	( 14'sd 6418) * $signed(input_fmap_203[7:0]) +
	( 16'sd 25848) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28386) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2398) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5597) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6501) * $signed(input_fmap_208[7:0]) +
	( 15'sd 12297) * $signed(input_fmap_209[7:0]) +
	( 14'sd 7600) * $signed(input_fmap_210[7:0]) +
	( 14'sd 7695) * $signed(input_fmap_211[7:0]) +
	( 13'sd 3926) * $signed(input_fmap_212[7:0]) +
	( 16'sd 31964) * $signed(input_fmap_213[7:0]) +
	( 11'sd 540) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6492) * $signed(input_fmap_215[7:0]) +
	( 14'sd 7095) * $signed(input_fmap_216[7:0]) +
	( 16'sd 25331) * $signed(input_fmap_217[7:0]) +
	( 16'sd 17538) * $signed(input_fmap_218[7:0]) +
	( 16'sd 16905) * $signed(input_fmap_219[7:0]) +
	( 15'sd 13260) * $signed(input_fmap_220[7:0]) +
	( 16'sd 20838) * $signed(input_fmap_221[7:0]) +
	( 16'sd 29753) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14598) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25523) * $signed(input_fmap_224[7:0]) +
	( 12'sd 1577) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10843) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9219) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31074) * $signed(input_fmap_228[7:0]) +
	( 14'sd 6573) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30475) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7727) * $signed(input_fmap_231[7:0]) +
	( 16'sd 19451) * $signed(input_fmap_232[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_233[7:0]) +
	( 11'sd 651) * $signed(input_fmap_234[7:0]) +
	( 15'sd 9096) * $signed(input_fmap_235[7:0]) +
	( 14'sd 4160) * $signed(input_fmap_236[7:0]) +
	( 16'sd 16558) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14553) * $signed(input_fmap_238[7:0]) +
	( 15'sd 11400) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23706) * $signed(input_fmap_240[7:0]) +
	( 15'sd 8526) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17949) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6014) * $signed(input_fmap_243[7:0]) +
	( 10'sd 418) * $signed(input_fmap_244[7:0]) +
	( 16'sd 26484) * $signed(input_fmap_245[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_246[7:0]) +
	( 16'sd 29825) * $signed(input_fmap_247[7:0]) +
	( 8'sd 100) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15067) * $signed(input_fmap_249[7:0]) +
	( 14'sd 6994) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12992) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26264) * $signed(input_fmap_252[7:0]) +
	( 16'sd 29152) * $signed(input_fmap_253[7:0]) +
	( 14'sd 6982) * $signed(input_fmap_254[7:0]) +
	( 15'sd 9665) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_205;
assign conv_mac_205 = 
	( 15'sd 13729) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27636) * $signed(input_fmap_1[7:0]) +
	( 15'sd 9102) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3413) * $signed(input_fmap_3[7:0]) +
	( 15'sd 9714) * $signed(input_fmap_4[7:0]) +
	( 15'sd 8831) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11026) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13570) * $signed(input_fmap_7[7:0]) +
	( 16'sd 20460) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13711) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7222) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6348) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12446) * $signed(input_fmap_12[7:0]) +
	( 14'sd 5489) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8561) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4942) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29184) * $signed(input_fmap_18[7:0]) +
	( 15'sd 8243) * $signed(input_fmap_19[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9985) * $signed(input_fmap_21[7:0]) +
	( 16'sd 16750) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8746) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5417) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24374) * $signed(input_fmap_25[7:0]) +
	( 16'sd 25236) * $signed(input_fmap_26[7:0]) +
	( 15'sd 14141) * $signed(input_fmap_27[7:0]) +
	( 15'sd 12229) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9606) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1663) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14226) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2294) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3785) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10759) * $signed(input_fmap_34[7:0]) +
	( 16'sd 30913) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6236) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11431) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22122) * $signed(input_fmap_38[7:0]) +
	( 13'sd 2243) * $signed(input_fmap_39[7:0]) +
	( 13'sd 2593) * $signed(input_fmap_40[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32192) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5880) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17645) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26956) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5467) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26911) * $signed(input_fmap_47[7:0]) +
	( 14'sd 7984) * $signed(input_fmap_48[7:0]) +
	( 16'sd 29575) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10324) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13119) * $signed(input_fmap_51[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3648) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31471) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19895) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6504) * $signed(input_fmap_57[7:0]) +
	( 15'sd 12593) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19796) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15393) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13764) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9654) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29070) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10907) * $signed(input_fmap_65[7:0]) +
	( 16'sd 18332) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22182) * $signed(input_fmap_67[7:0]) +
	( 16'sd 16944) * $signed(input_fmap_68[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_69[7:0]) +
	( 16'sd 29795) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16726) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25774) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10711) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15706) * $signed(input_fmap_74[7:0]) +
	( 16'sd 19110) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1100) * $signed(input_fmap_77[7:0]) +
	( 13'sd 4004) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11061) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30604) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2976) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8602) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28331) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15443) * $signed(input_fmap_84[7:0]) +
	( 13'sd 3799) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4652) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18637) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7604) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14450) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8753) * $signed(input_fmap_90[7:0]) +
	( 15'sd 12250) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11796) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_94[7:0]) +
	( 16'sd 27190) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3219) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3109) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9129) * $signed(input_fmap_99[7:0]) +
	( 16'sd 20635) * $signed(input_fmap_100[7:0]) +
	( 15'sd 11518) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16093) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31477) * $signed(input_fmap_103[7:0]) +
	( 16'sd 18482) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21836) * $signed(input_fmap_105[7:0]) +
	( 16'sd 16594) * $signed(input_fmap_106[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12837) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21321) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1305) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3234) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11746) * $signed(input_fmap_112[7:0]) +
	( 15'sd 14470) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32611) * $signed(input_fmap_114[7:0]) +
	( 16'sd 24037) * $signed(input_fmap_115[7:0]) +
	( 16'sd 25818) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2519) * $signed(input_fmap_117[7:0]) +
	( 16'sd 23427) * $signed(input_fmap_118[7:0]) +
	( 12'sd 1651) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29784) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17745) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31260) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5607) * $signed(input_fmap_123[7:0]) +
	( 16'sd 31316) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14850) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25882) * $signed(input_fmap_126[7:0]) +
	( 14'sd 4232) * $signed(input_fmap_127[7:0]) +
	( 16'sd 24971) * $signed(input_fmap_128[7:0]) +
	( 16'sd 18377) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_131[7:0]) +
	( 15'sd 9950) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12744) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2716) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27108) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15382) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25445) * $signed(input_fmap_137[7:0]) +
	( 16'sd 23461) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2977) * $signed(input_fmap_139[7:0]) +
	( 16'sd 22719) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13470) * $signed(input_fmap_141[7:0]) +
	( 16'sd 16896) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23812) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31884) * $signed(input_fmap_144[7:0]) +
	( 16'sd 30593) * $signed(input_fmap_145[7:0]) +
	( 14'sd 5386) * $signed(input_fmap_146[7:0]) +
	( 14'sd 7558) * $signed(input_fmap_147[7:0]) +
	( 15'sd 15126) * $signed(input_fmap_148[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_149[7:0]) +
	( 16'sd 29162) * $signed(input_fmap_150[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6831) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31009) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20686) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24136) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22452) * $signed(input_fmap_157[7:0]) +
	( 16'sd 27987) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26199) * $signed(input_fmap_159[7:0]) +
	( 16'sd 16537) * $signed(input_fmap_160[7:0]) +
	( 16'sd 17688) * $signed(input_fmap_161[7:0]) +
	( 16'sd 22351) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26491) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_164[7:0]) +
	( 15'sd 12623) * $signed(input_fmap_165[7:0]) +
	( 16'sd 22918) * $signed(input_fmap_166[7:0]) +
	( 15'sd 15469) * $signed(input_fmap_167[7:0]) +
	( 16'sd 17829) * $signed(input_fmap_168[7:0]) +
	( 9'sd 224) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11412) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_171[7:0]) +
	( 14'sd 4842) * $signed(input_fmap_172[7:0]) +
	( 15'sd 8587) * $signed(input_fmap_173[7:0]) +
	( 14'sd 8167) * $signed(input_fmap_174[7:0]) +
	( 16'sd 31306) * $signed(input_fmap_175[7:0]) +
	( 15'sd 13714) * $signed(input_fmap_176[7:0]) +
	( 15'sd 16109) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1730) * $signed(input_fmap_178[7:0]) +
	( 15'sd 11558) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21468) * $signed(input_fmap_180[7:0]) +
	( 16'sd 26411) * $signed(input_fmap_181[7:0]) +
	( 15'sd 8722) * $signed(input_fmap_182[7:0]) +
	( 11'sd 1013) * $signed(input_fmap_183[7:0]) +
	( 16'sd 25152) * $signed(input_fmap_184[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_185[7:0]) +
	( 16'sd 16841) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2666) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23614) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11676) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17846) * $signed(input_fmap_191[7:0]) +
	( 15'sd 13057) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10781) * $signed(input_fmap_193[7:0]) +
	( 16'sd 20036) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25957) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5848) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10474) * $signed(input_fmap_197[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28629) * $signed(input_fmap_199[7:0]) +
	( 16'sd 24224) * $signed(input_fmap_200[7:0]) +
	( 15'sd 11821) * $signed(input_fmap_201[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_202[7:0]) +
	( 14'sd 8135) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12763) * $signed(input_fmap_204[7:0]) +
	( 16'sd 17440) * $signed(input_fmap_205[7:0]) +
	( 15'sd 13396) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21054) * $signed(input_fmap_207[7:0]) +
	( 15'sd 11227) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13362) * $signed(input_fmap_209[7:0]) +
	( 16'sd 27459) * $signed(input_fmap_210[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_211[7:0]) +
	( 11'sd 607) * $signed(input_fmap_212[7:0]) +
	( 16'sd 20163) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31993) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9131) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5780) * $signed(input_fmap_216[7:0]) +
	( 16'sd 26084) * $signed(input_fmap_217[7:0]) +
	( 16'sd 24429) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19376) * $signed(input_fmap_219[7:0]) +
	( 14'sd 5641) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5913) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25856) * $signed(input_fmap_222[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30715) * $signed(input_fmap_224[7:0]) +
	( 15'sd 8341) * $signed(input_fmap_225[7:0]) +
	( 16'sd 25779) * $signed(input_fmap_226[7:0]) +
	( 16'sd 31726) * $signed(input_fmap_227[7:0]) +
	( 16'sd 23704) * $signed(input_fmap_228[7:0]) +
	( 15'sd 9742) * $signed(input_fmap_229[7:0]) +
	( 16'sd 16766) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20430) * $signed(input_fmap_231[7:0]) +
	( 12'sd 1929) * $signed(input_fmap_232[7:0]) +
	( 11'sd 721) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5791) * $signed(input_fmap_234[7:0]) +
	( 10'sd 309) * $signed(input_fmap_235[7:0]) +
	( 15'sd 16037) * $signed(input_fmap_236[7:0]) +
	( 16'sd 22899) * $signed(input_fmap_237[7:0]) +
	( 16'sd 31568) * $signed(input_fmap_238[7:0]) +
	( 16'sd 29743) * $signed(input_fmap_239[7:0]) +
	( 10'sd 344) * $signed(input_fmap_240[7:0]) +
	( 15'sd 8977) * $signed(input_fmap_241[7:0]) +
	( 15'sd 13477) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2736) * $signed(input_fmap_243[7:0]) +
	( 16'sd 29870) * $signed(input_fmap_244[7:0]) +
	( 11'sd 877) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1854) * $signed(input_fmap_246[7:0]) +
	( 15'sd 16175) * $signed(input_fmap_247[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21431) * $signed(input_fmap_249[7:0]) +
	( 15'sd 16381) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14561) * $signed(input_fmap_251[7:0]) +
	( 16'sd 25661) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17741) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31169) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20577) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_206;
assign conv_mac_206 = 
	( 16'sd 16959) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31462) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5100) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30330) * $signed(input_fmap_3[7:0]) +
	( 12'sd 1251) * $signed(input_fmap_4[7:0]) +
	( 11'sd 889) * $signed(input_fmap_5[7:0]) +
	( 16'sd 27320) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13138) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11523) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7792) * $signed(input_fmap_10[7:0]) +
	( 16'sd 20113) * $signed(input_fmap_11[7:0]) +
	( 15'sd 16157) * $signed(input_fmap_12[7:0]) +
	( 14'sd 6186) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1840) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9465) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28540) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4584) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4460) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1699) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20020) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25309) * $signed(input_fmap_21[7:0]) +
	( 13'sd 2531) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29316) * $signed(input_fmap_23[7:0]) +
	( 16'sd 31405) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21387) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_26[7:0]) +
	( 16'sd 32311) * $signed(input_fmap_27[7:0]) +
	( 9'sd 132) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5813) * $signed(input_fmap_29[7:0]) +
	( 12'sd 1702) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20468) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2740) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22222) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8422) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21188) * $signed(input_fmap_35[7:0]) +
	( 15'sd 15937) * $signed(input_fmap_36[7:0]) +
	( 16'sd 21129) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24564) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3998) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13604) * $signed(input_fmap_41[7:0]) +
	( 16'sd 22538) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19317) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20732) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23280) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13959) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19247) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12558) * $signed(input_fmap_49[7:0]) +
	( 15'sd 8461) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32182) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21405) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1470) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11806) * $signed(input_fmap_54[7:0]) +
	( 16'sd 28809) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28811) * $signed(input_fmap_56[7:0]) +
	( 16'sd 22846) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10934) * $signed(input_fmap_58[7:0]) +
	( 16'sd 28796) * $signed(input_fmap_59[7:0]) +
	( 16'sd 20449) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24850) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13629) * $signed(input_fmap_62[7:0]) +
	( 16'sd 17662) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13537) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10965) * $signed(input_fmap_65[7:0]) +
	( 15'sd 8937) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32123) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2987) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22374) * $signed(input_fmap_70[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1606) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10659) * $signed(input_fmap_73[7:0]) +
	( 16'sd 22889) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30703) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29768) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10933) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5116) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25622) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24305) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19444) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9955) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2233) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11262) * $signed(input_fmap_84[7:0]) +
	( 14'sd 7678) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20165) * $signed(input_fmap_87[7:0]) +
	( 16'sd 23622) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14651) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3041) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28649) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25135) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32085) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10247) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31552) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21261) * $signed(input_fmap_96[7:0]) +
	( 16'sd 32613) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10673) * $signed(input_fmap_98[7:0]) +
	( 16'sd 23529) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23759) * $signed(input_fmap_100[7:0]) +
	( 15'sd 13282) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29853) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2837) * $signed(input_fmap_103[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_104[7:0]) +
	( 16'sd 32679) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3940) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29348) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30309) * $signed(input_fmap_108[7:0]) +
	( 16'sd 17826) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12076) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22699) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_112[7:0]) +
	( 15'sd 13803) * $signed(input_fmap_113[7:0]) +
	( 11'sd 755) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2919) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4948) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24056) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5897) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22876) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1149) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15862) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29447) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3404) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9397) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22958) * $signed(input_fmap_125[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21830) * $signed(input_fmap_127[7:0]) +
	( 16'sd 18199) * $signed(input_fmap_128[7:0]) +
	( 15'sd 11282) * $signed(input_fmap_129[7:0]) +
	( 13'sd 2211) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14666) * $signed(input_fmap_131[7:0]) +
	( 15'sd 15955) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22076) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25615) * $signed(input_fmap_134[7:0]) +
	( 14'sd 4236) * $signed(input_fmap_135[7:0]) +
	( 16'sd 26559) * $signed(input_fmap_136[7:0]) +
	( 13'sd 3477) * $signed(input_fmap_137[7:0]) +
	( 15'sd 15707) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2941) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1438) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31867) * $signed(input_fmap_141[7:0]) +
	( 15'sd 12152) * $signed(input_fmap_142[7:0]) +
	( 16'sd 28699) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13418) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28809) * $signed(input_fmap_145[7:0]) +
	( 16'sd 26249) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21548) * $signed(input_fmap_147[7:0]) +
	( 16'sd 32321) * $signed(input_fmap_148[7:0]) +
	( 16'sd 16688) * $signed(input_fmap_149[7:0]) +
	( 16'sd 22570) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12258) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14239) * $signed(input_fmap_152[7:0]) +
	( 14'sd 7939) * $signed(input_fmap_153[7:0]) +
	( 16'sd 20762) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27333) * $signed(input_fmap_155[7:0]) +
	( 15'sd 9254) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31759) * $signed(input_fmap_157[7:0]) +
	( 16'sd 29086) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20310) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5720) * $signed(input_fmap_160[7:0]) +
	( 16'sd 30589) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10430) * $signed(input_fmap_162[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_163[7:0]) +
	( 16'sd 21057) * $signed(input_fmap_164[7:0]) +
	( 16'sd 17859) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19299) * $signed(input_fmap_166[7:0]) +
	( 16'sd 27046) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9023) * $signed(input_fmap_168[7:0]) +
	( 16'sd 23966) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_170[7:0]) +
	( 15'sd 12907) * $signed(input_fmap_171[7:0]) +
	( 16'sd 32375) * $signed(input_fmap_172[7:0]) +
	( 16'sd 27301) * $signed(input_fmap_173[7:0]) +
	( 14'sd 8057) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1312) * $signed(input_fmap_175[7:0]) +
	( 15'sd 15360) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18865) * $signed(input_fmap_177[7:0]) +
	( 16'sd 17817) * $signed(input_fmap_178[7:0]) +
	( 16'sd 26140) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6605) * $signed(input_fmap_180[7:0]) +
	( 16'sd 29760) * $signed(input_fmap_181[7:0]) +
	( 16'sd 32215) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5951) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26751) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17197) * $signed(input_fmap_185[7:0]) +
	( 16'sd 16806) * $signed(input_fmap_186[7:0]) +
	( 16'sd 29526) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12429) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5591) * $signed(input_fmap_189[7:0]) +
	( 13'sd 2222) * $signed(input_fmap_190[7:0]) +
	( 16'sd 27999) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_193[7:0]) +
	( 15'sd 16343) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17825) * $signed(input_fmap_195[7:0]) +
	( 15'sd 13620) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10166) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22790) * $signed(input_fmap_198[7:0]) +
	( 15'sd 13856) * $signed(input_fmap_199[7:0]) +
	( 16'sd 19609) * $signed(input_fmap_200[7:0]) +
	( 14'sd 7587) * $signed(input_fmap_201[7:0]) +
	( 13'sd 3371) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24506) * $signed(input_fmap_203[7:0]) +
	( 16'sd 29544) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5752) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28893) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18953) * $signed(input_fmap_207[7:0]) +
	( 16'sd 26143) * $signed(input_fmap_208[7:0]) +
	( 15'sd 15231) * $signed(input_fmap_209[7:0]) +
	( 16'sd 20609) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12262) * $signed(input_fmap_211[7:0]) +
	( 14'sd 7209) * $signed(input_fmap_212[7:0]) +
	( 14'sd 8146) * $signed(input_fmap_213[7:0]) +
	( 13'sd 2568) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1626) * $signed(input_fmap_215[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_216[7:0]) +
	( 15'sd 15110) * $signed(input_fmap_217[7:0]) +
	( 12'sd 1750) * $signed(input_fmap_218[7:0]) +
	( 12'sd 1838) * $signed(input_fmap_219[7:0]) +
	( 15'sd 8727) * $signed(input_fmap_220[7:0]) +
	( 16'sd 18045) * $signed(input_fmap_221[7:0]) +
	( 16'sd 29190) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17838) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13545) * $signed(input_fmap_224[7:0]) +
	( 14'sd 4662) * $signed(input_fmap_225[7:0]) +
	( 16'sd 19714) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24864) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1447) * $signed(input_fmap_228[7:0]) +
	( 15'sd 12826) * $signed(input_fmap_229[7:0]) +
	( 15'sd 11752) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_231[7:0]) +
	( 16'sd 21543) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15360) * $signed(input_fmap_233[7:0]) +
	( 13'sd 2617) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12676) * $signed(input_fmap_235[7:0]) +
	( 15'sd 13014) * $signed(input_fmap_236[7:0]) +
	( 16'sd 18071) * $signed(input_fmap_237[7:0]) +
	( 16'sd 17678) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5973) * $signed(input_fmap_239[7:0]) +
	( 16'sd 23924) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11529) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13954) * $signed(input_fmap_243[7:0]) +
	( 16'sd 21832) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24991) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28784) * $signed(input_fmap_246[7:0]) +
	( 16'sd 29321) * $signed(input_fmap_247[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14232) * $signed(input_fmap_249[7:0]) +
	( 15'sd 14632) * $signed(input_fmap_250[7:0]) +
	( 14'sd 5931) * $signed(input_fmap_251[7:0]) +
	( 15'sd 14522) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5728) * $signed(input_fmap_253[7:0]) +
	( 16'sd 19231) * $signed(input_fmap_254[7:0]) +
	( 16'sd 21531) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_207;
assign conv_mac_207 = 
	( 16'sd 30748) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31322) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26088) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23935) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16206) * $signed(input_fmap_4[7:0]) +
	( 15'sd 10228) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24616) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20411) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19964) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6307) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25584) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23727) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5185) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15497) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27065) * $signed(input_fmap_14[7:0]) +
	( 15'sd 11583) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25648) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13059) * $signed(input_fmap_17[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4996) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12238) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5403) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18762) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23210) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_24[7:0]) +
	( 16'sd 23425) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24993) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8334) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19948) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22941) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26237) * $signed(input_fmap_30[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6417) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21572) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7635) * $signed(input_fmap_34[7:0]) +
	( 16'sd 28088) * $signed(input_fmap_35[7:0]) +
	( 16'sd 16747) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8929) * $signed(input_fmap_37[7:0]) +
	( 16'sd 16614) * $signed(input_fmap_38[7:0]) +
	( 11'sd 528) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25688) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13128) * $signed(input_fmap_41[7:0]) +
	( 11'sd 976) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20993) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19944) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7095) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18077) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29014) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24678) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11974) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5800) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27779) * $signed(input_fmap_52[7:0]) +
	( 13'sd 2479) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11065) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29421) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19481) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25130) * $signed(input_fmap_57[7:0]) +
	( 16'sd 32391) * $signed(input_fmap_58[7:0]) +
	( 13'sd 2152) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13030) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24305) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8907) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24308) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22323) * $signed(input_fmap_64[7:0]) +
	( 16'sd 16809) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25525) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24686) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20227) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16864) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6867) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25741) * $signed(input_fmap_71[7:0]) +
	( 11'sd 614) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25161) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20097) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25921) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3197) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18872) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19213) * $signed(input_fmap_78[7:0]) +
	( 16'sd 28703) * $signed(input_fmap_79[7:0]) +
	( 14'sd 8189) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19716) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14391) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31778) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28930) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10239) * $signed(input_fmap_85[7:0]) +
	( 15'sd 10109) * $signed(input_fmap_86[7:0]) +
	( 16'sd 30327) * $signed(input_fmap_87[7:0]) +
	( 16'sd 20468) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9872) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31995) * $signed(input_fmap_90[7:0]) +
	( 15'sd 14175) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18101) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1666) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26356) * $signed(input_fmap_94[7:0]) +
	( 13'sd 3309) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31868) * $signed(input_fmap_96[7:0]) +
	( 14'sd 6037) * $signed(input_fmap_97[7:0]) +
	( 14'sd 6945) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3995) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28569) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6529) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16578) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31518) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31823) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13768) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13922) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14943) * $signed(input_fmap_107[7:0]) +
	( 15'sd 13474) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8711) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9950) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21130) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27271) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5846) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29021) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5721) * $signed(input_fmap_115[7:0]) +
	( 16'sd 16401) * $signed(input_fmap_116[7:0]) +
	( 14'sd 7783) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30253) * $signed(input_fmap_118[7:0]) +
	( 16'sd 20372) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22545) * $signed(input_fmap_120[7:0]) +
	( 12'sd 2004) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2886) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9399) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24814) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3520) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6288) * $signed(input_fmap_126[7:0]) +
	( 16'sd 25015) * $signed(input_fmap_127[7:0]) +
	( 15'sd 11883) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13592) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_130[7:0]) +
	( 13'sd 2342) * $signed(input_fmap_131[7:0]) +
	( 7'sd 51) * $signed(input_fmap_132[7:0]) +
	( 16'sd 20467) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19680) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28834) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25431) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9611) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18717) * $signed(input_fmap_139[7:0]) +
	( 16'sd 19169) * $signed(input_fmap_140[7:0]) +
	( 15'sd 13330) * $signed(input_fmap_141[7:0]) +
	( 15'sd 13213) * $signed(input_fmap_142[7:0]) +
	( 16'sd 21884) * $signed(input_fmap_143[7:0]) +
	( 15'sd 10305) * $signed(input_fmap_144[7:0]) +
	( 16'sd 24532) * $signed(input_fmap_145[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_147[7:0]) +
	( 15'sd 12835) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17284) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5181) * $signed(input_fmap_150[7:0]) +
	( 13'sd 2640) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24449) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31249) * $signed(input_fmap_153[7:0]) +
	( 15'sd 13823) * $signed(input_fmap_154[7:0]) +
	( 15'sd 14276) * $signed(input_fmap_155[7:0]) +
	( 15'sd 11808) * $signed(input_fmap_156[7:0]) +
	( 16'sd 18619) * $signed(input_fmap_157[7:0]) +
	( 16'sd 27333) * $signed(input_fmap_158[7:0]) +
	( 16'sd 28624) * $signed(input_fmap_159[7:0]) +
	( 13'sd 2776) * $signed(input_fmap_160[7:0]) +
	( 16'sd 29853) * $signed(input_fmap_161[7:0]) +
	( 16'sd 28474) * $signed(input_fmap_162[7:0]) +
	( 15'sd 10402) * $signed(input_fmap_163[7:0]) +
	( 16'sd 29804) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9160) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9947) * $signed(input_fmap_166[7:0]) +
	( 12'sd 1519) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29745) * $signed(input_fmap_168[7:0]) +
	( 16'sd 28435) * $signed(input_fmap_169[7:0]) +
	( 16'sd 32111) * $signed(input_fmap_170[7:0]) +
	( 16'sd 32125) * $signed(input_fmap_171[7:0]) +
	( 15'sd 8704) * $signed(input_fmap_172[7:0]) +
	( 16'sd 17692) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27284) * $signed(input_fmap_174[7:0]) +
	( 15'sd 15358) * $signed(input_fmap_175[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_176[7:0]) +
	( 15'sd 13466) * $signed(input_fmap_177[7:0]) +
	( 16'sd 20629) * $signed(input_fmap_178[7:0]) +
	( 15'sd 13535) * $signed(input_fmap_179[7:0]) +
	( 15'sd 13573) * $signed(input_fmap_180[7:0]) +
	( 15'sd 9783) * $signed(input_fmap_181[7:0]) +
	( 16'sd 17130) * $signed(input_fmap_182[7:0]) +
	( 16'sd 32564) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13430) * $signed(input_fmap_184[7:0]) +
	( 16'sd 30125) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9437) * $signed(input_fmap_186[7:0]) +
	( 12'sd 1113) * $signed(input_fmap_187[7:0]) +
	( 15'sd 15009) * $signed(input_fmap_188[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_189[7:0]) +
	( 15'sd 11170) * $signed(input_fmap_190[7:0]) +
	( 16'sd 16624) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29895) * $signed(input_fmap_192[7:0]) +
	( 12'sd 1269) * $signed(input_fmap_193[7:0]) +
	( 14'sd 4830) * $signed(input_fmap_194[7:0]) +
	( 15'sd 10985) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20304) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14527) * $signed(input_fmap_197[7:0]) +
	( 16'sd 18881) * $signed(input_fmap_198[7:0]) +
	( 16'sd 32068) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6227) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3104) * $signed(input_fmap_201[7:0]) +
	( 16'sd 28320) * $signed(input_fmap_202[7:0]) +
	( 16'sd 32287) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17732) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5152) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3298) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1127) * $signed(input_fmap_207[7:0]) +
	( 15'sd 9097) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11346) * $signed(input_fmap_209[7:0]) +
	( 14'sd 4115) * $signed(input_fmap_210[7:0]) +
	( 11'sd 561) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_212[7:0]) +
	( 16'sd 31091) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15183) * $signed(input_fmap_214[7:0]) +
	( 15'sd 15422) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18384) * $signed(input_fmap_216[7:0]) +
	( 13'sd 3623) * $signed(input_fmap_217[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_218[7:0]) +
	( 15'sd 8360) * $signed(input_fmap_219[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1406) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18197) * $signed(input_fmap_222[7:0]) +
	( 15'sd 13701) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13102) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13604) * $signed(input_fmap_225[7:0]) +
	( 16'sd 24455) * $signed(input_fmap_226[7:0]) +
	( 16'sd 24149) * $signed(input_fmap_227[7:0]) +
	( 16'sd 30434) * $signed(input_fmap_228[7:0]) +
	( 11'sd 955) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29007) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7335) * $signed(input_fmap_231[7:0]) +
	( 16'sd 27396) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10662) * $signed(input_fmap_233[7:0]) +
	( 12'sd 1204) * $signed(input_fmap_234[7:0]) +
	( 12'sd 1839) * $signed(input_fmap_235[7:0]) +
	( 16'sd 22177) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28735) * $signed(input_fmap_237[7:0]) +
	( 16'sd 31633) * $signed(input_fmap_238[7:0]) +
	( 13'sd 2637) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25661) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15707) * $signed(input_fmap_241[7:0]) +
	( 16'sd 28464) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13707) * $signed(input_fmap_243[7:0]) +
	( 16'sd 31432) * $signed(input_fmap_244[7:0]) +
	( 15'sd 11552) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23995) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18249) * $signed(input_fmap_247[7:0]) +
	( 15'sd 9975) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15947) * $signed(input_fmap_249[7:0]) +
	( 16'sd 31980) * $signed(input_fmap_250[7:0]) +
	( 16'sd 25832) * $signed(input_fmap_251[7:0]) +
	( 10'sd 348) * $signed(input_fmap_252[7:0]) +
	( 16'sd 19857) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2135) * $signed(input_fmap_254[7:0]) +
	( 16'sd 28636) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_208;
assign conv_mac_208 = 
	( 16'sd 20763) * $signed(input_fmap_0[7:0]) +
	( 15'sd 8452) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7629) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31272) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25381) * $signed(input_fmap_4[7:0]) +
	( 11'sd 714) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3261) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9360) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23589) * $signed(input_fmap_8[7:0]) +
	( 15'sd 16320) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12161) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19916) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23514) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11041) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10733) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28487) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6314) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6108) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29016) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28809) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26638) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24468) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31746) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18707) * $signed(input_fmap_23[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15678) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24911) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_27[7:0]) +
	( 15'sd 8923) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15649) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3038) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15864) * $signed(input_fmap_31[7:0]) +
	( 14'sd 7325) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12278) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14927) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6396) * $signed(input_fmap_35[7:0]) +
	( 14'sd 4678) * $signed(input_fmap_36[7:0]) +
	( 14'sd 4257) * $signed(input_fmap_37[7:0]) +
	( 16'sd 26658) * $signed(input_fmap_38[7:0]) +
	( 16'sd 18946) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25490) * $signed(input_fmap_40[7:0]) +
	( 13'sd 2612) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18094) * $signed(input_fmap_42[7:0]) +
	( 16'sd 28031) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9221) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20985) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5047) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_47[7:0]) +
	( 14'sd 8037) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20618) * $signed(input_fmap_49[7:0]) +
	( 9'sd 210) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25620) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3706) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12050) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18456) * $signed(input_fmap_54[7:0]) +
	( 13'sd 3670) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3745) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15476) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6643) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17550) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13830) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24663) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23619) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15464) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11955) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31224) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20174) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12487) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1196) * $signed(input_fmap_68[7:0]) +
	( 16'sd 32418) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16535) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8472) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26323) * $signed(input_fmap_72[7:0]) +
	( 16'sd 17470) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12228) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9640) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31736) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10880) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3329) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20421) * $signed(input_fmap_80[7:0]) +
	( 16'sd 24181) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9716) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6567) * $signed(input_fmap_84[7:0]) +
	( 15'sd 11055) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13573) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22180) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14920) * $signed(input_fmap_88[7:0]) +
	( 16'sd 26537) * $signed(input_fmap_89[7:0]) +
	( 15'sd 13625) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31982) * $signed(input_fmap_92[7:0]) +
	( 15'sd 12155) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3080) * $signed(input_fmap_94[7:0]) +
	( 16'sd 32478) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1570) * $signed(input_fmap_96[7:0]) +
	( 16'sd 23313) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_98[7:0]) +
	( 15'sd 16322) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_100[7:0]) +
	( 16'sd 18517) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32728) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2811) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17885) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4623) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5187) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32616) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7320) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12628) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24752) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18253) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11252) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15205) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20605) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9767) * $signed(input_fmap_116[7:0]) +
	( 15'sd 10312) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7442) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24134) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18924) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9165) * $signed(input_fmap_121[7:0]) +
	( 9'sd 176) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21098) * $signed(input_fmap_123[7:0]) +
	( 7'sd 45) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24536) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29609) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9700) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13346) * $signed(input_fmap_129[7:0]) +
	( 16'sd 18110) * $signed(input_fmap_130[7:0]) +
	( 16'sd 27613) * $signed(input_fmap_131[7:0]) +
	( 16'sd 23130) * $signed(input_fmap_132[7:0]) +
	( 16'sd 23027) * $signed(input_fmap_133[7:0]) +
	( 15'sd 8510) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27270) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7724) * $signed(input_fmap_136[7:0]) +
	( 14'sd 4246) * $signed(input_fmap_137[7:0]) +
	( 16'sd 21673) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11279) * $signed(input_fmap_139[7:0]) +
	( 14'sd 4934) * $signed(input_fmap_140[7:0]) +
	( 16'sd 30770) * $signed(input_fmap_141[7:0]) +
	( 16'sd 16858) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_143[7:0]) +
	( 15'sd 15281) * $signed(input_fmap_144[7:0]) +
	( 14'sd 5162) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14498) * $signed(input_fmap_146[7:0]) +
	( 16'sd 20419) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6550) * $signed(input_fmap_148[7:0]) +
	( 15'sd 14706) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9877) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14324) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7917) * $signed(input_fmap_152[7:0]) +
	( 16'sd 18665) * $signed(input_fmap_153[7:0]) +
	( 16'sd 18811) * $signed(input_fmap_154[7:0]) +
	( 12'sd 1581) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10849) * $signed(input_fmap_156[7:0]) +
	( 15'sd 9374) * $signed(input_fmap_157[7:0]) +
	( 16'sd 32310) * $signed(input_fmap_158[7:0]) +
	( 16'sd 21340) * $signed(input_fmap_159[7:0]) +
	( 12'sd 1738) * $signed(input_fmap_160[7:0]) +
	( 16'sd 29645) * $signed(input_fmap_161[7:0]) +
	( 14'sd 6875) * $signed(input_fmap_162[7:0]) +
	( 16'sd 29141) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19864) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22434) * $signed(input_fmap_165[7:0]) +
	( 15'sd 15562) * $signed(input_fmap_166[7:0]) +
	( 16'sd 21945) * $signed(input_fmap_167[7:0]) +
	( 15'sd 12746) * $signed(input_fmap_168[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9254) * $signed(input_fmap_170[7:0]) +
	( 12'sd 1153) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31064) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12717) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26913) * $signed(input_fmap_174[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21853) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7677) * $signed(input_fmap_177[7:0]) +
	( 16'sd 30983) * $signed(input_fmap_178[7:0]) +
	( 14'sd 5823) * $signed(input_fmap_179[7:0]) +
	( 14'sd 5852) * $signed(input_fmap_180[7:0]) +
	( 16'sd 24773) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5250) * $signed(input_fmap_182[7:0]) +
	( 16'sd 19490) * $signed(input_fmap_183[7:0]) +
	( 14'sd 4237) * $signed(input_fmap_184[7:0]) +
	( 16'sd 31411) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26138) * $signed(input_fmap_186[7:0]) +
	( 15'sd 15502) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29900) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3742) * $signed(input_fmap_189[7:0]) +
	( 16'sd 29839) * $signed(input_fmap_190[7:0]) +
	( 13'sd 2221) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31544) * $signed(input_fmap_192[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30626) * $signed(input_fmap_194[7:0]) +
	( 16'sd 32734) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12406) * $signed(input_fmap_196[7:0]) +
	( 14'sd 6816) * $signed(input_fmap_197[7:0]) +
	( 15'sd 11360) * $signed(input_fmap_198[7:0]) +
	( 16'sd 21958) * $signed(input_fmap_199[7:0]) +
	( 11'sd 808) * $signed(input_fmap_200[7:0]) +
	( 16'sd 31346) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31918) * $signed(input_fmap_202[7:0]) +
	( 15'sd 15936) * $signed(input_fmap_203[7:0]) +
	( 16'sd 23227) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12343) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27658) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29050) * $signed(input_fmap_207[7:0]) +
	( 15'sd 13542) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24819) * $signed(input_fmap_209[7:0]) +
	( 16'sd 17799) * $signed(input_fmap_210[7:0]) +
	( 11'sd 857) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19830) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23638) * $signed(input_fmap_213[7:0]) +
	( 15'sd 12682) * $signed(input_fmap_214[7:0]) +
	( 16'sd 20627) * $signed(input_fmap_215[7:0]) +
	( 16'sd 32117) * $signed(input_fmap_216[7:0]) +
	( 16'sd 21445) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22218) * $signed(input_fmap_218[7:0]) +
	( 16'sd 26628) * $signed(input_fmap_219[7:0]) +
	( 16'sd 32155) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6034) * $signed(input_fmap_221[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8233) * $signed(input_fmap_223[7:0]) +
	( 13'sd 2077) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5890) * $signed(input_fmap_225[7:0]) +
	( 16'sd 24021) * $signed(input_fmap_226[7:0]) +
	( 11'sd 754) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10543) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24860) * $signed(input_fmap_229[7:0]) +
	( 15'sd 8996) * $signed(input_fmap_230[7:0]) +
	( 15'sd 15346) * $signed(input_fmap_231[7:0]) +
	( 14'sd 7166) * $signed(input_fmap_232[7:0]) +
	( 16'sd 23865) * $signed(input_fmap_233[7:0]) +
	( 16'sd 21410) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14658) * $signed(input_fmap_235[7:0]) +
	( 13'sd 2845) * $signed(input_fmap_236[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28248) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19255) * $signed(input_fmap_239[7:0]) +
	( 15'sd 13300) * $signed(input_fmap_240[7:0]) +
	( 15'sd 15800) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11556) * $signed(input_fmap_242[7:0]) +
	( 16'sd 19494) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22737) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24512) * $signed(input_fmap_245[7:0]) +
	( 16'sd 30644) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21100) * $signed(input_fmap_247[7:0]) +
	( 15'sd 11614) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2520) * $signed(input_fmap_249[7:0]) +
	( 16'sd 20473) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27349) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28392) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6261) * $signed(input_fmap_253[7:0]) +
	( 11'sd 644) * $signed(input_fmap_254[7:0]) +
	( 13'sd 2137) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_209;
assign conv_mac_209 = 
	( 16'sd 17476) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27766) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27052) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23765) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5126) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27944) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30570) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28691) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15107) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30424) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28738) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28710) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27351) * $signed(input_fmap_13[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28884) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5240) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25218) * $signed(input_fmap_17[7:0]) +
	( 16'sd 28449) * $signed(input_fmap_18[7:0]) +
	( 7'sd 32) * $signed(input_fmap_19[7:0]) +
	( 14'sd 5296) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19279) * $signed(input_fmap_21[7:0]) +
	( 15'sd 10370) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7793) * $signed(input_fmap_23[7:0]) +
	( 15'sd 16101) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16555) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21455) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17527) * $signed(input_fmap_27[7:0]) +
	( 16'sd 20674) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11452) * $signed(input_fmap_29[7:0]) +
	( 15'sd 15088) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15723) * $signed(input_fmap_33[7:0]) +
	( 9'sd 198) * $signed(input_fmap_34[7:0]) +
	( 14'sd 7415) * $signed(input_fmap_35[7:0]) +
	( 15'sd 14066) * $signed(input_fmap_36[7:0]) +
	( 16'sd 28157) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3389) * $signed(input_fmap_38[7:0]) +
	( 16'sd 22904) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31983) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15071) * $signed(input_fmap_41[7:0]) +
	( 16'sd 21172) * $signed(input_fmap_42[7:0]) +
	( 16'sd 19031) * $signed(input_fmap_43[7:0]) +
	( 16'sd 30458) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20086) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7865) * $signed(input_fmap_46[7:0]) +
	( 15'sd 11015) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8515) * $signed(input_fmap_48[7:0]) +
	( 16'sd 20882) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17904) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31935) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15436) * $signed(input_fmap_52[7:0]) +
	( 12'sd 1803) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15223) * $signed(input_fmap_55[7:0]) +
	( 11'sd 534) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21178) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19238) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16558) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26950) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19625) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21012) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24438) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10853) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3065) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17856) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31188) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12236) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11487) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6447) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3189) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3091) * $signed(input_fmap_72[7:0]) +
	( 13'sd 3019) * $signed(input_fmap_73[7:0]) +
	( 16'sd 19180) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14208) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8402) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31350) * $signed(input_fmap_77[7:0]) +
	( 8'sd 80) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17148) * $signed(input_fmap_79[7:0]) +
	( 11'sd 679) * $signed(input_fmap_80[7:0]) +
	( 15'sd 16054) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11967) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18253) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16072) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4330) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20678) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1210) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1196) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32259) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19390) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16476) * $signed(input_fmap_91[7:0]) +
	( 16'sd 21503) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15302) * $signed(input_fmap_93[7:0]) +
	( 16'sd 30800) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16436) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15786) * $signed(input_fmap_96[7:0]) +
	( 16'sd 24665) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28590) * $signed(input_fmap_98[7:0]) +
	( 16'sd 25420) * $signed(input_fmap_99[7:0]) +
	( 16'sd 27233) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27585) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5065) * $signed(input_fmap_102[7:0]) +
	( 16'sd 22122) * $signed(input_fmap_103[7:0]) +
	( 16'sd 19216) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27071) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11743) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2940) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27340) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5414) * $signed(input_fmap_109[7:0]) +
	( 14'sd 4516) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10964) * $signed(input_fmap_111[7:0]) +
	( 15'sd 12090) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17543) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18494) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15156) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9150) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28036) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2499) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29077) * $signed(input_fmap_120[7:0]) +
	( 16'sd 18259) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5927) * $signed(input_fmap_122[7:0]) +
	( 11'sd 952) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24490) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16549) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3490) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17972) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4321) * $signed(input_fmap_128[7:0]) +
	( 16'sd 29551) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22530) * $signed(input_fmap_130[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_131[7:0]) +
	( 16'sd 16405) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21741) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_134[7:0]) +
	( 14'sd 5671) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2541) * $signed(input_fmap_136[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_137[7:0]) +
	( 15'sd 9332) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2924) * $signed(input_fmap_139[7:0]) +
	( 16'sd 20978) * $signed(input_fmap_140[7:0]) +
	( 16'sd 23945) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8249) * $signed(input_fmap_142[7:0]) +
	( 16'sd 24456) * $signed(input_fmap_143[7:0]) +
	( 14'sd 7225) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22337) * $signed(input_fmap_145[7:0]) +
	( 14'sd 6011) * $signed(input_fmap_146[7:0]) +
	( 16'sd 26661) * $signed(input_fmap_147[7:0]) +
	( 16'sd 28908) * $signed(input_fmap_148[7:0]) +
	( 15'sd 11766) * $signed(input_fmap_149[7:0]) +
	( 13'sd 3175) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23393) * $signed(input_fmap_151[7:0]) +
	( 15'sd 8902) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4270) * $signed(input_fmap_153[7:0]) +
	( 15'sd 16378) * $signed(input_fmap_154[7:0]) +
	( 15'sd 8941) * $signed(input_fmap_155[7:0]) +
	( 16'sd 30159) * $signed(input_fmap_156[7:0]) +
	( 15'sd 10672) * $signed(input_fmap_157[7:0]) +
	( 16'sd 19101) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_159[7:0]) +
	( 16'sd 29258) * $signed(input_fmap_160[7:0]) +
	( 14'sd 4706) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30526) * $signed(input_fmap_162[7:0]) +
	( 16'sd 25024) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1253) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30756) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3238) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24003) * $signed(input_fmap_167[7:0]) +
	( 14'sd 7441) * $signed(input_fmap_168[7:0]) +
	( 11'sd 678) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5056) * $signed(input_fmap_170[7:0]) +
	( 16'sd 28807) * $signed(input_fmap_171[7:0]) +
	( 16'sd 20780) * $signed(input_fmap_172[7:0]) +
	( 16'sd 21359) * $signed(input_fmap_173[7:0]) +
	( 16'sd 20164) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7124) * $signed(input_fmap_175[7:0]) +
	( 13'sd 3690) * $signed(input_fmap_176[7:0]) +
	( 2'sd 1) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14955) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6688) * $signed(input_fmap_179[7:0]) +
	( 15'sd 11923) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30687) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26888) * $signed(input_fmap_182[7:0]) +
	( 15'sd 12047) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15542) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9602) * $signed(input_fmap_186[7:0]) +
	( 10'sd 272) * $signed(input_fmap_187[7:0]) +
	( 16'sd 20097) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2070) * $signed(input_fmap_189[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20318) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27835) * $signed(input_fmap_192[7:0]) +
	( 14'sd 5290) * $signed(input_fmap_193[7:0]) +
	( 16'sd 17707) * $signed(input_fmap_194[7:0]) +
	( 16'sd 29647) * $signed(input_fmap_195[7:0]) +
	( 12'sd 1741) * $signed(input_fmap_196[7:0]) +
	( 15'sd 8425) * $signed(input_fmap_197[7:0]) +
	( 16'sd 26486) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16249) * $signed(input_fmap_199[7:0]) +
	( 15'sd 10815) * $signed(input_fmap_200[7:0]) +
	( 10'sd 506) * $signed(input_fmap_201[7:0]) +
	( 15'sd 12843) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21845) * $signed(input_fmap_203[7:0]) +
	( 16'sd 25986) * $signed(input_fmap_204[7:0]) +
	( 16'sd 26700) * $signed(input_fmap_205[7:0]) +
	( 15'sd 10747) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5499) * $signed(input_fmap_207[7:0]) +
	( 15'sd 9835) * $signed(input_fmap_208[7:0]) +
	( 14'sd 4992) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19773) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5446) * $signed(input_fmap_211[7:0]) +
	( 16'sd 31137) * $signed(input_fmap_212[7:0]) +
	( 15'sd 10380) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23293) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10655) * $signed(input_fmap_215[7:0]) +
	( 15'sd 13971) * $signed(input_fmap_216[7:0]) +
	( 16'sd 19099) * $signed(input_fmap_217[7:0]) +
	( 16'sd 18310) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5605) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30007) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19390) * $signed(input_fmap_221[7:0]) +
	( 16'sd 20656) * $signed(input_fmap_222[7:0]) +
	( 16'sd 26956) * $signed(input_fmap_223[7:0]) +
	( 11'sd 571) * $signed(input_fmap_224[7:0]) +
	( 15'sd 12190) * $signed(input_fmap_225[7:0]) +
	( 16'sd 20282) * $signed(input_fmap_226[7:0]) +
	( 16'sd 23105) * $signed(input_fmap_227[7:0]) +
	( 16'sd 21097) * $signed(input_fmap_228[7:0]) +
	( 16'sd 30514) * $signed(input_fmap_229[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20071) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8268) * $signed(input_fmap_232[7:0]) +
	( 14'sd 6585) * $signed(input_fmap_233[7:0]) +
	( 16'sd 28172) * $signed(input_fmap_234[7:0]) +
	( 14'sd 4509) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11303) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29179) * $signed(input_fmap_237[7:0]) +
	( 14'sd 8145) * $signed(input_fmap_238[7:0]) +
	( 13'sd 3414) * $signed(input_fmap_239[7:0]) +
	( 13'sd 3837) * $signed(input_fmap_240[7:0]) +
	( 15'sd 11984) * $signed(input_fmap_241[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_242[7:0]) +
	( 14'sd 8022) * $signed(input_fmap_243[7:0]) +
	( 15'sd 11242) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30888) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22013) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9252) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26025) * $signed(input_fmap_248[7:0]) +
	( 15'sd 10462) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32280) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21590) * $signed(input_fmap_251[7:0]) +
	( 16'sd 16765) * $signed(input_fmap_252[7:0]) +
	( 15'sd 8821) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2397) * $signed(input_fmap_254[7:0]) +
	( 14'sd 4832) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_210;
assign conv_mac_210 = 
	( 10'sd 264) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7140) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7144) * $signed(input_fmap_3[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_4[7:0]) +
	( 15'sd 9777) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20335) * $signed(input_fmap_6[7:0]) +
	( 16'sd 23277) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28046) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26749) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16801) * $signed(input_fmap_10[7:0]) +
	( 16'sd 28302) * $signed(input_fmap_11[7:0]) +
	( 15'sd 9546) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22516) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21842) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28214) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1897) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15577) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4727) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13133) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20070) * $signed(input_fmap_20[7:0]) +
	( 16'sd 19885) * $signed(input_fmap_21[7:0]) +
	( 15'sd 8575) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29864) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14456) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21575) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24871) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18000) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31318) * $signed(input_fmap_28[7:0]) +
	( 15'sd 16009) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18630) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4395) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22573) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16186) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30669) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9590) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12642) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9683) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4537) * $signed(input_fmap_38[7:0]) +
	( 16'sd 27991) * $signed(input_fmap_39[7:0]) +
	( 16'sd 28904) * $signed(input_fmap_40[7:0]) +
	( 15'sd 9519) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_42[7:0]) +
	( 11'sd 568) * $signed(input_fmap_43[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_44[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7999) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19696) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28515) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16542) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12072) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22488) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6758) * $signed(input_fmap_52[7:0]) +
	( 11'sd 538) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15058) * $signed(input_fmap_54[7:0]) +
	( 14'sd 5924) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13179) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15933) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18448) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20234) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32189) * $signed(input_fmap_60[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24546) * $signed(input_fmap_62[7:0]) +
	( 13'sd 3167) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5602) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19579) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32142) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17755) * $signed(input_fmap_67[7:0]) +
	( 12'sd 1755) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25211) * $signed(input_fmap_69[7:0]) +
	( 16'sd 32566) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27957) * $signed(input_fmap_71[7:0]) +
	( 10'sd 310) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1029) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24608) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31328) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15856) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16647) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9481) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8796) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21964) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30444) * $signed(input_fmap_81[7:0]) +
	( 16'sd 16863) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21134) * $signed(input_fmap_83[7:0]) +
	( 16'sd 26157) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23743) * $signed(input_fmap_85[7:0]) +
	( 15'sd 9908) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29306) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_88[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17505) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6882) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25272) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19537) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22930) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18813) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4668) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30549) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17689) * $signed(input_fmap_98[7:0]) +
	( 11'sd 978) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4237) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20551) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27228) * $signed(input_fmap_102[7:0]) +
	( 16'sd 26417) * $signed(input_fmap_103[7:0]) +
	( 10'sd 357) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24733) * $signed(input_fmap_105[7:0]) +
	( 16'sd 29175) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27492) * $signed(input_fmap_107[7:0]) +
	( 14'sd 6990) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20697) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14725) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29905) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31000) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29294) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15624) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9991) * $signed(input_fmap_116[7:0]) +
	( 16'sd 20911) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2707) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18297) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11392) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1552) * $signed(input_fmap_121[7:0]) +
	( 16'sd 23995) * $signed(input_fmap_122[7:0]) +
	( 16'sd 23974) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21360) * $signed(input_fmap_124[7:0]) +
	( 16'sd 18872) * $signed(input_fmap_125[7:0]) +
	( 13'sd 3585) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27324) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31184) * $signed(input_fmap_128[7:0]) +
	( 15'sd 11351) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12406) * $signed(input_fmap_130[7:0]) +
	( 16'sd 18105) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8237) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18227) * $signed(input_fmap_134[7:0]) +
	( 11'sd 907) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2302) * $signed(input_fmap_136[7:0]) +
	( 16'sd 20854) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31791) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14537) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29654) * $signed(input_fmap_140[7:0]) +
	( 16'sd 21810) * $signed(input_fmap_141[7:0]) +
	( 16'sd 29747) * $signed(input_fmap_142[7:0]) +
	( 15'sd 8987) * $signed(input_fmap_143[7:0]) +
	( 16'sd 26552) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21595) * $signed(input_fmap_145[7:0]) +
	( 15'sd 14779) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3904) * $signed(input_fmap_147[7:0]) +
	( 16'sd 18895) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7797) * $signed(input_fmap_149[7:0]) +
	( 16'sd 30937) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28808) * $signed(input_fmap_151[7:0]) +
	( 15'sd 12186) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31722) * $signed(input_fmap_153[7:0]) +
	( 16'sd 26501) * $signed(input_fmap_154[7:0]) +
	( 14'sd 6542) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15733) * $signed(input_fmap_156[7:0]) +
	( 16'sd 26630) * $signed(input_fmap_157[7:0]) +
	( 16'sd 29430) * $signed(input_fmap_158[7:0]) +
	( 16'sd 25962) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11608) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22857) * $signed(input_fmap_161[7:0]) +
	( 13'sd 3798) * $signed(input_fmap_162[7:0]) +
	( 15'sd 9506) * $signed(input_fmap_163[7:0]) +
	( 14'sd 7725) * $signed(input_fmap_164[7:0]) +
	( 15'sd 16037) * $signed(input_fmap_165[7:0]) +
	( 14'sd 4595) * $signed(input_fmap_166[7:0]) +
	( 15'sd 11148) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14473) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26185) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18263) * $signed(input_fmap_170[7:0]) +
	( 15'sd 9808) * $signed(input_fmap_171[7:0]) +
	( 14'sd 7863) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5755) * $signed(input_fmap_173[7:0]) +
	( 16'sd 27853) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5097) * $signed(input_fmap_175[7:0]) +
	( 16'sd 23482) * $signed(input_fmap_176[7:0]) +
	( 16'sd 24440) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1526) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20553) * $signed(input_fmap_179[7:0]) +
	( 13'sd 3038) * $signed(input_fmap_180[7:0]) +
	( 16'sd 19491) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26850) * $signed(input_fmap_182[7:0]) +
	( 13'sd 3067) * $signed(input_fmap_183[7:0]) +
	( 16'sd 31925) * $signed(input_fmap_184[7:0]) +
	( 14'sd 7146) * $signed(input_fmap_185[7:0]) +
	( 16'sd 30838) * $signed(input_fmap_186[7:0]) +
	( 15'sd 12240) * $signed(input_fmap_187[7:0]) +
	( 15'sd 13262) * $signed(input_fmap_188[7:0]) +
	( 16'sd 21926) * $signed(input_fmap_189[7:0]) +
	( 15'sd 11948) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24823) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24318) * $signed(input_fmap_192[7:0]) +
	( 10'sd 472) * $signed(input_fmap_193[7:0]) +
	( 15'sd 8962) * $signed(input_fmap_194[7:0]) +
	( 15'sd 9041) * $signed(input_fmap_195[7:0]) +
	( 15'sd 9469) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24940) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24033) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28850) * $signed(input_fmap_199[7:0]) +
	( 14'sd 7426) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22407) * $signed(input_fmap_201[7:0]) +
	( 16'sd 17860) * $signed(input_fmap_202[7:0]) +
	( 15'sd 9669) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12486) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5285) * $signed(input_fmap_205[7:0]) +
	( 13'sd 3978) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29397) * $signed(input_fmap_207[7:0]) +
	( 13'sd 3442) * $signed(input_fmap_208[7:0]) +
	( 15'sd 8413) * $signed(input_fmap_209[7:0]) +
	( 16'sd 26760) * $signed(input_fmap_210[7:0]) +
	( 14'sd 5599) * $signed(input_fmap_211[7:0]) +
	( 14'sd 7801) * $signed(input_fmap_212[7:0]) +
	( 11'sd 788) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7855) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_215[7:0]) +
	( 15'sd 10267) * $signed(input_fmap_216[7:0]) +
	( 16'sd 16994) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21907) * $signed(input_fmap_218[7:0]) +
	( 9'sd 190) * $signed(input_fmap_219[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23650) * $signed(input_fmap_221[7:0]) +
	( 11'sd 971) * $signed(input_fmap_222[7:0]) +
	( 16'sd 19488) * $signed(input_fmap_223[7:0]) +
	( 15'sd 11072) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2558) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27429) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20978) * $signed(input_fmap_227[7:0]) +
	( 14'sd 4533) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23488) * $signed(input_fmap_229[7:0]) +
	( 15'sd 13611) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7638) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14887) * $signed(input_fmap_232[7:0]) +
	( 15'sd 12193) * $signed(input_fmap_233[7:0]) +
	( 16'sd 28738) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19599) * $signed(input_fmap_235[7:0]) +
	( 14'sd 6185) * $signed(input_fmap_236[7:0]) +
	( 16'sd 22697) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27858) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21739) * $signed(input_fmap_239[7:0]) +
	( 16'sd 30477) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26508) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_242[7:0]) +
	( 12'sd 1362) * $signed(input_fmap_243[7:0]) +
	( 15'sd 9820) * $signed(input_fmap_244[7:0]) +
	( 12'sd 1140) * $signed(input_fmap_245[7:0]) +
	( 16'sd 29001) * $signed(input_fmap_246[7:0]) +
	( 16'sd 25952) * $signed(input_fmap_247[7:0]) +
	( 16'sd 22143) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24579) * $signed(input_fmap_249[7:0]) +
	( 16'sd 20777) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7484) * $signed(input_fmap_251[7:0]) +
	( 14'sd 7950) * $signed(input_fmap_252[7:0]) +
	( 16'sd 22748) * $signed(input_fmap_253[7:0]) +
	( 16'sd 16540) * $signed(input_fmap_254[7:0]) +
	( 15'sd 10066) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_211;
assign conv_mac_211 = 
	( 14'sd 5236) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4767) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8566) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15127) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13626) * $signed(input_fmap_4[7:0]) +
	( 10'sd 466) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20686) * $signed(input_fmap_7[7:0]) +
	( 15'sd 16219) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24755) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9911) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17233) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27083) * $signed(input_fmap_12[7:0]) +
	( 16'sd 27239) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17043) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2613) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22137) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31855) * $signed(input_fmap_17[7:0]) +
	( 16'sd 25215) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23345) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20744) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27728) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29468) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26036) * $signed(input_fmap_24[7:0]) +
	( 12'sd 1689) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23201) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7034) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19017) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_29[7:0]) +
	( 16'sd 21745) * $signed(input_fmap_30[7:0]) +
	( 16'sd 29613) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10889) * $signed(input_fmap_32[7:0]) +
	( 15'sd 15620) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12373) * $signed(input_fmap_34[7:0]) +
	( 13'sd 2594) * $signed(input_fmap_35[7:0]) +
	( 9'sd 224) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10099) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24334) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31279) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11660) * $signed(input_fmap_40[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9278) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2185) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23574) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21778) * $signed(input_fmap_45[7:0]) +
	( 11'sd 983) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26945) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9680) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24854) * $signed(input_fmap_49[7:0]) +
	( 14'sd 7001) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6921) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13783) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10537) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13650) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5770) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12767) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9807) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14799) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4513) * $signed(input_fmap_60[7:0]) +
	( 6'sd 19) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32242) * $signed(input_fmap_62[7:0]) +
	( 16'sd 28282) * $signed(input_fmap_63[7:0]) +
	( 14'sd 8154) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22196) * $signed(input_fmap_66[7:0]) +
	( 16'sd 23465) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11317) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29523) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13596) * $signed(input_fmap_70[7:0]) +
	( 15'sd 8769) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24276) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2747) * $signed(input_fmap_73[7:0]) +
	( 14'sd 4791) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31427) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_76[7:0]) +
	( 15'sd 12946) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2663) * $signed(input_fmap_78[7:0]) +
	( 16'sd 21131) * $signed(input_fmap_79[7:0]) +
	( 10'sd 316) * $signed(input_fmap_80[7:0]) +
	( 16'sd 26509) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_82[7:0]) +
	( 13'sd 4033) * $signed(input_fmap_83[7:0]) +
	( 15'sd 14399) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31421) * $signed(input_fmap_85[7:0]) +
	( 13'sd 2901) * $signed(input_fmap_86[7:0]) +
	( 7'sd 63) * $signed(input_fmap_87[7:0]) +
	( 15'sd 14888) * $signed(input_fmap_88[7:0]) +
	( 11'sd 799) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24957) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11744) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17777) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22844) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12753) * $signed(input_fmap_94[7:0]) +
	( 16'sd 21542) * $signed(input_fmap_95[7:0]) +
	( 13'sd 3244) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17464) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12347) * $signed(input_fmap_98[7:0]) +
	( 16'sd 17233) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31940) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7840) * $signed(input_fmap_101[7:0]) +
	( 11'sd 803) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9359) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20616) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1096) * $signed(input_fmap_105[7:0]) +
	( 14'sd 7102) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32255) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23468) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24975) * $signed(input_fmap_109[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11280) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30295) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24158) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25145) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15114) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29169) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20785) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32425) * $signed(input_fmap_119[7:0]) +
	( 14'sd 7137) * $signed(input_fmap_120[7:0]) +
	( 16'sd 24257) * $signed(input_fmap_121[7:0]) +
	( 12'sd 2017) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12086) * $signed(input_fmap_123[7:0]) +
	( 9'sd 217) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24841) * $signed(input_fmap_125[7:0]) +
	( 16'sd 32220) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12233) * $signed(input_fmap_127[7:0]) +
	( 16'sd 29044) * $signed(input_fmap_128[7:0]) +
	( 16'sd 32099) * $signed(input_fmap_129[7:0]) +
	( 16'sd 20068) * $signed(input_fmap_130[7:0]) +
	( 16'sd 30749) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10933) * $signed(input_fmap_132[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31986) * $signed(input_fmap_134[7:0]) +
	( 16'sd 22940) * $signed(input_fmap_135[7:0]) +
	( 16'sd 26405) * $signed(input_fmap_136[7:0]) +
	( 16'sd 23012) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19935) * $signed(input_fmap_138[7:0]) +
	( 15'sd 12856) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24195) * $signed(input_fmap_140[7:0]) +
	( 15'sd 15703) * $signed(input_fmap_141[7:0]) +
	( 14'sd 4947) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10680) * $signed(input_fmap_143[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_145[7:0]) +
	( 13'sd 4013) * $signed(input_fmap_146[7:0]) +
	( 16'sd 18972) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4604) * $signed(input_fmap_148[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27157) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17650) * $signed(input_fmap_151[7:0]) +
	( 16'sd 17375) * $signed(input_fmap_152[7:0]) +
	( 16'sd 30099) * $signed(input_fmap_153[7:0]) +
	( 15'sd 14751) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19565) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18405) * $signed(input_fmap_156[7:0]) +
	( 16'sd 24434) * $signed(input_fmap_157[7:0]) +
	( 16'sd 32277) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5499) * $signed(input_fmap_159[7:0]) +
	( 15'sd 16248) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23068) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24795) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15889) * $signed(input_fmap_163[7:0]) +
	( 15'sd 13624) * $signed(input_fmap_164[7:0]) +
	( 15'sd 11249) * $signed(input_fmap_165[7:0]) +
	( 16'sd 28856) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26941) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1138) * $signed(input_fmap_168[7:0]) +
	( 14'sd 7684) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31007) * $signed(input_fmap_170[7:0]) +
	( 16'sd 19725) * $signed(input_fmap_171[7:0]) +
	( 16'sd 23948) * $signed(input_fmap_172[7:0]) +
	( 16'sd 25765) * $signed(input_fmap_173[7:0]) +
	( 10'sd 307) * $signed(input_fmap_174[7:0]) +
	( 16'sd 22848) * $signed(input_fmap_175[7:0]) +
	( 16'sd 22278) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27672) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32693) * $signed(input_fmap_178[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_179[7:0]) +
	( 16'sd 25575) * $signed(input_fmap_180[7:0]) +
	( 16'sd 21208) * $signed(input_fmap_181[7:0]) +
	( 15'sd 16119) * $signed(input_fmap_182[7:0]) +
	( 15'sd 9694) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5503) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9843) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27508) * $signed(input_fmap_187[7:0]) +
	( 16'sd 16502) * $signed(input_fmap_188[7:0]) +
	( 16'sd 23914) * $signed(input_fmap_189[7:0]) +
	( 16'sd 21812) * $signed(input_fmap_190[7:0]) +
	( 15'sd 12443) * $signed(input_fmap_191[7:0]) +
	( 13'sd 2971) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6783) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18794) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5297) * $signed(input_fmap_195[7:0]) +
	( 16'sd 25688) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24880) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_198[7:0]) +
	( 16'sd 30485) * $signed(input_fmap_199[7:0]) +
	( 16'sd 28436) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27885) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18665) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5046) * $signed(input_fmap_203[7:0]) +
	( 15'sd 15955) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29680) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_206[7:0]) +
	( 16'sd 26173) * $signed(input_fmap_207[7:0]) +
	( 15'sd 13656) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23631) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3598) * $signed(input_fmap_210[7:0]) +
	( 16'sd 18912) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11592) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29996) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28849) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29911) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1162) * $signed(input_fmap_216[7:0]) +
	( 16'sd 31691) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28735) * $signed(input_fmap_218[7:0]) +
	( 16'sd 20229) * $signed(input_fmap_219[7:0]) +
	( 16'sd 18634) * $signed(input_fmap_220[7:0]) +
	( 11'sd 967) * $signed(input_fmap_221[7:0]) +
	( 15'sd 9486) * $signed(input_fmap_222[7:0]) +
	( 16'sd 30053) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1910) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26550) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18536) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3038) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24000) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26159) * $signed(input_fmap_229[7:0]) +
	( 15'sd 9205) * $signed(input_fmap_230[7:0]) +
	( 15'sd 10333) * $signed(input_fmap_231[7:0]) +
	( 16'sd 22886) * $signed(input_fmap_232[7:0]) +
	( 12'sd 1479) * $signed(input_fmap_233[7:0]) +
	( 15'sd 9693) * $signed(input_fmap_234[7:0]) +
	( 16'sd 21651) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23751) * $signed(input_fmap_236[7:0]) +
	( 15'sd 13126) * $signed(input_fmap_237[7:0]) +
	( 14'sd 7088) * $signed(input_fmap_238[7:0]) +
	( 16'sd 22027) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26498) * $signed(input_fmap_240[7:0]) +
	( 14'sd 8099) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11080) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28229) * $signed(input_fmap_243[7:0]) +
	( 16'sd 32178) * $signed(input_fmap_244[7:0]) +
	( 14'sd 4124) * $signed(input_fmap_245[7:0]) +
	( 16'sd 27658) * $signed(input_fmap_246[7:0]) +
	( 14'sd 4210) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32306) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24862) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12275) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15104) * $signed(input_fmap_251[7:0]) +
	( 15'sd 8312) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25026) * $signed(input_fmap_253[7:0]) +
	( 13'sd 3596) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24720) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_212;
assign conv_mac_212 = 
	( 11'sd 710) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10588) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16741) * $signed(input_fmap_2[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_3[7:0]) +
	( 16'sd 19012) * $signed(input_fmap_4[7:0]) +
	( 11'sd 564) * $signed(input_fmap_5[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_6[7:0]) +
	( 16'sd 17501) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13633) * $signed(input_fmap_8[7:0]) +
	( 15'sd 13160) * $signed(input_fmap_9[7:0]) +
	( 14'sd 6250) * $signed(input_fmap_10[7:0]) +
	( 16'sd 22275) * $signed(input_fmap_11[7:0]) +
	( 15'sd 10443) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19083) * $signed(input_fmap_13[7:0]) +
	( 13'sd 4073) * $signed(input_fmap_14[7:0]) +
	( 15'sd 13135) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_16[7:0]) +
	( 14'sd 4625) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10951) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29185) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19743) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2810) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21866) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1451) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17883) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18385) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31279) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12556) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26925) * $signed(input_fmap_30[7:0]) +
	( 16'sd 20325) * $signed(input_fmap_31[7:0]) +
	( 16'sd 30795) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3957) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13014) * $signed(input_fmap_34[7:0]) +
	( 14'sd 5595) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_36[7:0]) +
	( 11'sd 825) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_38[7:0]) +
	( 11'sd 764) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21637) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21598) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11538) * $signed(input_fmap_42[7:0]) +
	( 16'sd 30964) * $signed(input_fmap_43[7:0]) +
	( 16'sd 20619) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4995) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16366) * $signed(input_fmap_46[7:0]) +
	( 12'sd 2046) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21556) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5286) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1453) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32085) * $signed(input_fmap_52[7:0]) +
	( 16'sd 29648) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10739) * $signed(input_fmap_54[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10216) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8922) * $signed(input_fmap_57[7:0]) +
	( 15'sd 13418) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29848) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29819) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16758) * $signed(input_fmap_61[7:0]) +
	( 15'sd 16208) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18226) * $signed(input_fmap_63[7:0]) +
	( 12'sd 1054) * $signed(input_fmap_64[7:0]) +
	( 14'sd 5897) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32473) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11044) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18628) * $signed(input_fmap_68[7:0]) +
	( 15'sd 11366) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13276) * $signed(input_fmap_70[7:0]) +
	( 14'sd 8049) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13583) * $signed(input_fmap_72[7:0]) +
	( 15'sd 16093) * $signed(input_fmap_73[7:0]) +
	( 16'sd 25931) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4164) * $signed(input_fmap_75[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30029) * $signed(input_fmap_77[7:0]) +
	( 16'sd 27270) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4550) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20290) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16919) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23144) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2544) * $signed(input_fmap_84[7:0]) +
	( 15'sd 15266) * $signed(input_fmap_85[7:0]) +
	( 16'sd 21019) * $signed(input_fmap_86[7:0]) +
	( 13'sd 2857) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13322) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10411) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24256) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1368) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10793) * $signed(input_fmap_92[7:0]) +
	( 16'sd 27898) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32013) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28062) * $signed(input_fmap_95[7:0]) +
	( 16'sd 31231) * $signed(input_fmap_96[7:0]) +
	( 13'sd 2773) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8572) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30654) * $signed(input_fmap_99[7:0]) +
	( 13'sd 2213) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26597) * $signed(input_fmap_101[7:0]) +
	( 16'sd 31926) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21405) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1235) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28519) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6176) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28092) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8364) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8849) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9558) * $signed(input_fmap_110[7:0]) +
	( 13'sd 2828) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23578) * $signed(input_fmap_112[7:0]) +
	( 15'sd 16089) * $signed(input_fmap_113[7:0]) +
	( 14'sd 4262) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30129) * $signed(input_fmap_115[7:0]) +
	( 12'sd 2031) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3554) * $signed(input_fmap_117[7:0]) +
	( 15'sd 12068) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21514) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6795) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6171) * $signed(input_fmap_121[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10938) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27746) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20870) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25643) * $signed(input_fmap_126[7:0]) +
	( 11'sd 707) * $signed(input_fmap_127[7:0]) +
	( 16'sd 28240) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10490) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1589) * $signed(input_fmap_130[7:0]) +
	( 16'sd 29771) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10269) * $signed(input_fmap_132[7:0]) +
	( 16'sd 28086) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11573) * $signed(input_fmap_134[7:0]) +
	( 15'sd 14595) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30603) * $signed(input_fmap_136[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27644) * $signed(input_fmap_138[7:0]) +
	( 16'sd 25967) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1844) * $signed(input_fmap_140[7:0]) +
	( 15'sd 15727) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22416) * $signed(input_fmap_142[7:0]) +
	( 16'sd 19835) * $signed(input_fmap_143[7:0]) +
	( 16'sd 17285) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27785) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1815) * $signed(input_fmap_146[7:0]) +
	( 14'sd 4911) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26850) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21539) * $signed(input_fmap_150[7:0]) +
	( 16'sd 29262) * $signed(input_fmap_151[7:0]) +
	( 14'sd 6907) * $signed(input_fmap_152[7:0]) +
	( 16'sd 19183) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11579) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10982) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14907) * $signed(input_fmap_156[7:0]) +
	( 12'sd 1227) * $signed(input_fmap_157[7:0]) +
	( 15'sd 13762) * $signed(input_fmap_158[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_159[7:0]) +
	( 15'sd 12981) * $signed(input_fmap_160[7:0]) +
	( 15'sd 14472) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10342) * $signed(input_fmap_162[7:0]) +
	( 16'sd 18872) * $signed(input_fmap_163[7:0]) +
	( 16'sd 20894) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22174) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9086) * $signed(input_fmap_166[7:0]) +
	( 12'sd 1059) * $signed(input_fmap_167[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_168[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_169[7:0]) +
	( 15'sd 13503) * $signed(input_fmap_170[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9005) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19857) * $signed(input_fmap_173[7:0]) +
	( 16'sd 21048) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21890) * $signed(input_fmap_175[7:0]) +
	( 16'sd 19042) * $signed(input_fmap_176[7:0]) +
	( 16'sd 20647) * $signed(input_fmap_177[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_178[7:0]) +
	( 16'sd 17238) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32376) * $signed(input_fmap_180[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_181[7:0]) +
	( 16'sd 25950) * $signed(input_fmap_182[7:0]) +
	( 14'sd 7435) * $signed(input_fmap_183[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3303) * $signed(input_fmap_185[7:0]) +
	( 15'sd 8816) * $signed(input_fmap_186[7:0]) +
	( 14'sd 8150) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2852) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17519) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13362) * $signed(input_fmap_190[7:0]) +
	( 16'sd 16568) * $signed(input_fmap_191[7:0]) +
	( 16'sd 26470) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9828) * $signed(input_fmap_193[7:0]) +
	( 8'sd 115) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22613) * $signed(input_fmap_195[7:0]) +
	( 16'sd 29936) * $signed(input_fmap_196[7:0]) +
	( 15'sd 15592) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9210) * $signed(input_fmap_198[7:0]) +
	( 14'sd 4610) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20911) * $signed(input_fmap_200[7:0]) +
	( 16'sd 23368) * $signed(input_fmap_201[7:0]) +
	( 15'sd 9169) * $signed(input_fmap_202[7:0]) +
	( 15'sd 15138) * $signed(input_fmap_203[7:0]) +
	( 13'sd 4088) * $signed(input_fmap_204[7:0]) +
	( 16'sd 20714) * $signed(input_fmap_205[7:0]) +
	( 15'sd 10176) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5661) * $signed(input_fmap_207[7:0]) +
	( 13'sd 3257) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3778) * $signed(input_fmap_209[7:0]) +
	( 13'sd 2298) * $signed(input_fmap_210[7:0]) +
	( 16'sd 27077) * $signed(input_fmap_211[7:0]) +
	( 15'sd 10812) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2874) * $signed(input_fmap_213[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22404) * $signed(input_fmap_215[7:0]) +
	( 14'sd 7127) * $signed(input_fmap_216[7:0]) +
	( 15'sd 15803) * $signed(input_fmap_217[7:0]) +
	( 15'sd 11713) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14344) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1136) * $signed(input_fmap_220[7:0]) +
	( 14'sd 5629) * $signed(input_fmap_221[7:0]) +
	( 14'sd 4380) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8424) * $signed(input_fmap_223[7:0]) +
	( 16'sd 29601) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_225[7:0]) +
	( 14'sd 6593) * $signed(input_fmap_226[7:0]) +
	( 15'sd 9105) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22687) * $signed(input_fmap_228[7:0]) +
	( 15'sd 11029) * $signed(input_fmap_229[7:0]) +
	( 9'sd 254) * $signed(input_fmap_230[7:0]) +
	( 16'sd 22516) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14130) * $signed(input_fmap_232[7:0]) +
	( 14'sd 6225) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15070) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22292) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31983) * $signed(input_fmap_236[7:0]) +
	( 15'sd 14456) * $signed(input_fmap_237[7:0]) +
	( 16'sd 24906) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9815) * $signed(input_fmap_239[7:0]) +
	( 16'sd 31415) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18607) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13758) * $signed(input_fmap_243[7:0]) +
	( 10'sd 413) * $signed(input_fmap_244[7:0]) +
	( 14'sd 4307) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23385) * $signed(input_fmap_246[7:0]) +
	( 16'sd 26052) * $signed(input_fmap_247[7:0]) +
	( 16'sd 24719) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3746) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26409) * $signed(input_fmap_250[7:0]) +
	( 16'sd 30033) * $signed(input_fmap_251[7:0]) +
	( 16'sd 22823) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28322) * $signed(input_fmap_253[7:0]) +
	( 16'sd 22471) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5828) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_213;
assign conv_mac_213 = 
	( 15'sd 8999) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20847) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13902) * $signed(input_fmap_2[7:0]) +
	( 16'sd 17771) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27436) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23453) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6614) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1293) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30496) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19422) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31499) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14836) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19477) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14637) * $signed(input_fmap_14[7:0]) +
	( 15'sd 10017) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30872) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17673) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6330) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27394) * $signed(input_fmap_19[7:0]) +
	( 16'sd 25046) * $signed(input_fmap_20[7:0]) +
	( 13'sd 2470) * $signed(input_fmap_21[7:0]) +
	( 16'sd 28367) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10997) * $signed(input_fmap_23[7:0]) +
	( 16'sd 29567) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9679) * $signed(input_fmap_25[7:0]) +
	( 13'sd 3982) * $signed(input_fmap_26[7:0]) +
	( 16'sd 28355) * $signed(input_fmap_27[7:0]) +
	( 16'sd 25332) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2084) * $signed(input_fmap_29[7:0]) +
	( 16'sd 23508) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28036) * $signed(input_fmap_31[7:0]) +
	( 16'sd 22165) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2951) * $signed(input_fmap_33[7:0]) +
	( 16'sd 26269) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1732) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25939) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6226) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3578) * $signed(input_fmap_38[7:0]) +
	( 15'sd 9895) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21202) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24265) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8632) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16036) * $signed(input_fmap_43[7:0]) +
	( 16'sd 24769) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5110) * $signed(input_fmap_46[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32729) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18088) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5317) * $signed(input_fmap_50[7:0]) +
	( 14'sd 6082) * $signed(input_fmap_51[7:0]) +
	( 16'sd 21621) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20204) * $signed(input_fmap_53[7:0]) +
	( 15'sd 14730) * $signed(input_fmap_54[7:0]) +
	( 14'sd 7614) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13851) * $signed(input_fmap_56[7:0]) +
	( 12'sd 2014) * $signed(input_fmap_57[7:0]) +
	( 16'sd 31377) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23202) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32425) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24844) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12959) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2509) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6318) * $signed(input_fmap_64[7:0]) +
	( 14'sd 7733) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6829) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19262) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19294) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10899) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20587) * $signed(input_fmap_70[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7623) * $signed(input_fmap_72[7:0]) +
	( 16'sd 19292) * $signed(input_fmap_73[7:0]) +
	( 15'sd 14120) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25219) * $signed(input_fmap_75[7:0]) +
	( 14'sd 5912) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11906) * $signed(input_fmap_77[7:0]) +
	( 16'sd 23354) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3617) * $signed(input_fmap_79[7:0]) +
	( 15'sd 8512) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2901) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6237) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21425) * $signed(input_fmap_83[7:0]) +
	( 16'sd 21166) * $signed(input_fmap_84[7:0]) +
	( 16'sd 17419) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25640) * $signed(input_fmap_87[7:0]) +
	( 16'sd 26408) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28283) * $signed(input_fmap_89[7:0]) +
	( 15'sd 11452) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8764) * $signed(input_fmap_91[7:0]) +
	( 15'sd 10445) * $signed(input_fmap_92[7:0]) +
	( 16'sd 18873) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25372) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23867) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_96[7:0]) +
	( 16'sd 31131) * $signed(input_fmap_97[7:0]) +
	( 16'sd 29120) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21792) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6254) * $signed(input_fmap_100[7:0]) +
	( 15'sd 10585) * $signed(input_fmap_101[7:0]) +
	( 13'sd 2856) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1918) * $signed(input_fmap_103[7:0]) +
	( 13'sd 2849) * $signed(input_fmap_104[7:0]) +
	( 16'sd 23805) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5604) * $signed(input_fmap_106[7:0]) +
	( 16'sd 32304) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14781) * $signed(input_fmap_108[7:0]) +
	( 11'sd 916) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5128) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6152) * $signed(input_fmap_111[7:0]) +
	( 12'sd 1130) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25469) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27102) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9346) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15466) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28297) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30949) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27874) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15004) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27817) * $signed(input_fmap_121[7:0]) +
	( 11'sd 581) * $signed(input_fmap_122[7:0]) +
	( 16'sd 16588) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13185) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13287) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20114) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26346) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9535) * $signed(input_fmap_128[7:0]) +
	( 14'sd 4773) * $signed(input_fmap_129[7:0]) +
	( 16'sd 28343) * $signed(input_fmap_130[7:0]) +
	( 13'sd 3947) * $signed(input_fmap_131[7:0]) +
	( 15'sd 11069) * $signed(input_fmap_132[7:0]) +
	( 16'sd 30778) * $signed(input_fmap_133[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_134[7:0]) +
	( 15'sd 11749) * $signed(input_fmap_135[7:0]) +
	( 16'sd 32408) * $signed(input_fmap_136[7:0]) +
	( 14'sd 7262) * $signed(input_fmap_137[7:0]) +
	( 14'sd 6864) * $signed(input_fmap_138[7:0]) +
	( 14'sd 6748) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29238) * $signed(input_fmap_140[7:0]) +
	( 16'sd 27546) * $signed(input_fmap_141[7:0]) +
	( 16'sd 29352) * $signed(input_fmap_142[7:0]) +
	( 14'sd 6003) * $signed(input_fmap_143[7:0]) +
	( 15'sd 13018) * $signed(input_fmap_144[7:0]) +
	( 15'sd 14110) * $signed(input_fmap_145[7:0]) +
	( 16'sd 23821) * $signed(input_fmap_146[7:0]) +
	( 16'sd 24552) * $signed(input_fmap_147[7:0]) +
	( 12'sd 1239) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23341) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21235) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19248) * $signed(input_fmap_151[7:0]) +
	( 16'sd 17133) * $signed(input_fmap_152[7:0]) +
	( 15'sd 9347) * $signed(input_fmap_153[7:0]) +
	( 15'sd 13356) * $signed(input_fmap_154[7:0]) +
	( 14'sd 6129) * $signed(input_fmap_155[7:0]) +
	( 12'sd 1571) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15425) * $signed(input_fmap_157[7:0]) +
	( 15'sd 9770) * $signed(input_fmap_158[7:0]) +
	( 14'sd 7954) * $signed(input_fmap_159[7:0]) +
	( 16'sd 23629) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19439) * $signed(input_fmap_161[7:0]) +
	( 15'sd 15835) * $signed(input_fmap_162[7:0]) +
	( 14'sd 5166) * $signed(input_fmap_163[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_164[7:0]) +
	( 12'sd 1759) * $signed(input_fmap_165[7:0]) +
	( 15'sd 8856) * $signed(input_fmap_166[7:0]) +
	( 16'sd 32733) * $signed(input_fmap_167[7:0]) +
	( 16'sd 30841) * $signed(input_fmap_168[7:0]) +
	( 16'sd 20034) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14786) * $signed(input_fmap_170[7:0]) +
	( 11'sd 679) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12307) * $signed(input_fmap_172[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6592) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3124) * $signed(input_fmap_175[7:0]) +
	( 16'sd 32634) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6460) * $signed(input_fmap_177[7:0]) +
	( 15'sd 10790) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22373) * $signed(input_fmap_179[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_180[7:0]) +
	( 15'sd 13850) * $signed(input_fmap_181[7:0]) +
	( 11'sd 835) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5941) * $signed(input_fmap_183[7:0]) +
	( 16'sd 20565) * $signed(input_fmap_184[7:0]) +
	( 15'sd 8882) * $signed(input_fmap_185[7:0]) +
	( 15'sd 8387) * $signed(input_fmap_186[7:0]) +
	( 16'sd 30710) * $signed(input_fmap_187[7:0]) +
	( 10'sd 478) * $signed(input_fmap_188[7:0]) +
	( 15'sd 13082) * $signed(input_fmap_189[7:0]) +
	( 16'sd 31007) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19331) * $signed(input_fmap_191[7:0]) +
	( 13'sd 3010) * $signed(input_fmap_192[7:0]) +
	( 13'sd 3320) * $signed(input_fmap_193[7:0]) +
	( 16'sd 29330) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5889) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5691) * $signed(input_fmap_196[7:0]) +
	( 16'sd 19167) * $signed(input_fmap_197[7:0]) +
	( 12'sd 1478) * $signed(input_fmap_198[7:0]) +
	( 16'sd 17898) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5628) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18217) * $signed(input_fmap_201[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_202[7:0]) +
	( 15'sd 8940) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32744) * $signed(input_fmap_204[7:0]) +
	( 15'sd 16063) * $signed(input_fmap_205[7:0]) +
	( 16'sd 17610) * $signed(input_fmap_206[7:0]) +
	( 15'sd 15435) * $signed(input_fmap_207[7:0]) +
	( 15'sd 13929) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30050) * $signed(input_fmap_210[7:0]) +
	( 14'sd 7506) * $signed(input_fmap_211[7:0]) +
	( 16'sd 25540) * $signed(input_fmap_212[7:0]) +
	( 16'sd 30301) * $signed(input_fmap_213[7:0]) +
	( 15'sd 11802) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2319) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24985) * $signed(input_fmap_216[7:0]) +
	( 14'sd 6733) * $signed(input_fmap_217[7:0]) +
	( 15'sd 8503) * $signed(input_fmap_218[7:0]) +
	( 16'sd 22776) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26215) * $signed(input_fmap_220[7:0]) +
	( 15'sd 10858) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19939) * $signed(input_fmap_222[7:0]) +
	( 14'sd 7899) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7319) * $signed(input_fmap_224[7:0]) +
	( 16'sd 32665) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10821) * $signed(input_fmap_226[7:0]) +
	( 16'sd 32370) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10917) * $signed(input_fmap_228[7:0]) +
	( 16'sd 32514) * $signed(input_fmap_229[7:0]) +
	( 16'sd 22465) * $signed(input_fmap_230[7:0]) +
	( 16'sd 27711) * $signed(input_fmap_231[7:0]) +
	( 13'sd 2239) * $signed(input_fmap_232[7:0]) +
	( 15'sd 15981) * $signed(input_fmap_233[7:0]) +
	( 16'sd 28872) * $signed(input_fmap_234[7:0]) +
	( 16'sd 26362) * $signed(input_fmap_235[7:0]) +
	( 16'sd 19756) * $signed(input_fmap_236[7:0]) +
	( 16'sd 23094) * $signed(input_fmap_237[7:0]) +
	( 14'sd 6672) * $signed(input_fmap_238[7:0]) +
	( 14'sd 7750) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25189) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3483) * $signed(input_fmap_241[7:0]) +
	( 15'sd 12581) * $signed(input_fmap_242[7:0]) +
	( 15'sd 9959) * $signed(input_fmap_243[7:0]) +
	( 16'sd 31292) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12390) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23589) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15549) * $signed(input_fmap_247[7:0]) +
	( 16'sd 23943) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12497) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3869) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12308) * $signed(input_fmap_251[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27102) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2667) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24327) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_214;
assign conv_mac_214 = 
	( 13'sd 3027) * $signed(input_fmap_0[7:0]) +
	( 16'sd 25572) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16809) * $signed(input_fmap_2[7:0]) +
	( 16'sd 31151) * $signed(input_fmap_3[7:0]) +
	( 16'sd 30748) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25303) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6909) * $signed(input_fmap_6[7:0]) +
	( 14'sd 5551) * $signed(input_fmap_7[7:0]) +
	( 16'sd 25608) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31619) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1638) * $signed(input_fmap_10[7:0]) +
	( 15'sd 8628) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27315) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25942) * $signed(input_fmap_13[7:0]) +
	( 16'sd 28676) * $signed(input_fmap_14[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23197) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17320) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23793) * $signed(input_fmap_18[7:0]) +
	( 15'sd 11216) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8452) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15037) * $signed(input_fmap_21[7:0]) +
	( 16'sd 20093) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17668) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11562) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14563) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8600) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29039) * $signed(input_fmap_27[7:0]) +
	( 15'sd 9838) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18261) * $signed(input_fmap_29[7:0]) +
	( 11'sd 843) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27016) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15237) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29370) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11798) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24319) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10700) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18807) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25126) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5880) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18134) * $signed(input_fmap_40[7:0]) +
	( 15'sd 12838) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15929) * $signed(input_fmap_42[7:0]) +
	( 16'sd 17350) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1392) * $signed(input_fmap_45[7:0]) +
	( 15'sd 11322) * $signed(input_fmap_46[7:0]) +
	( 15'sd 10159) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8399) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27880) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19278) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23127) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9636) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10670) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8765) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25008) * $signed(input_fmap_55[7:0]) +
	( 16'sd 21953) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24217) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28846) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11187) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11282) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21788) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1401) * $signed(input_fmap_62[7:0]) +
	( 15'sd 14829) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10293) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20748) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11770) * $signed(input_fmap_66[7:0]) +
	( 16'sd 21614) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21833) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14636) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23247) * $signed(input_fmap_70[7:0]) +
	( 14'sd 4244) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19853) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27314) * $signed(input_fmap_73[7:0]) +
	( 16'sd 27397) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25953) * $signed(input_fmap_75[7:0]) +
	( 16'sd 16888) * $signed(input_fmap_76[7:0]) +
	( 14'sd 5915) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13929) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3733) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9739) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25898) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1711) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31213) * $signed(input_fmap_83[7:0]) +
	( 6'sd 22) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24318) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22249) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18818) * $signed(input_fmap_87[7:0]) +
	( 15'sd 8264) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2282) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20739) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28026) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19312) * $signed(input_fmap_92[7:0]) +
	( 14'sd 6959) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12779) * $signed(input_fmap_94[7:0]) +
	( 16'sd 26347) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22002) * $signed(input_fmap_96[7:0]) +
	( 15'sd 13051) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4857) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5954) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24596) * $signed(input_fmap_100[7:0]) +
	( 16'sd 22152) * $signed(input_fmap_101[7:0]) +
	( 16'sd 17093) * $signed(input_fmap_102[7:0]) +
	( 15'sd 12553) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27514) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4582) * $signed(input_fmap_105[7:0]) +
	( 16'sd 25339) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3938) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27936) * $signed(input_fmap_108[7:0]) +
	( 14'sd 7237) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24843) * $signed(input_fmap_110[7:0]) +
	( 15'sd 11073) * $signed(input_fmap_111[7:0]) +
	( 13'sd 2903) * $signed(input_fmap_112[7:0]) +
	( 10'sd 458) * $signed(input_fmap_113[7:0]) +
	( 16'sd 31677) * $signed(input_fmap_114[7:0]) +
	( 11'sd 751) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27705) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29426) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13867) * $signed(input_fmap_118[7:0]) +
	( 16'sd 23740) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10867) * $signed(input_fmap_120[7:0]) +
	( 13'sd 3821) * $signed(input_fmap_121[7:0]) +
	( 15'sd 10268) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7924) * $signed(input_fmap_123[7:0]) +
	( 16'sd 30150) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25591) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14713) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29120) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9923) * $signed(input_fmap_128[7:0]) +
	( 15'sd 9309) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12285) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15572) * $signed(input_fmap_131[7:0]) +
	( 15'sd 13971) * $signed(input_fmap_132[7:0]) +
	( 16'sd 17497) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25132) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27305) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17759) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27242) * $signed(input_fmap_137[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_138[7:0]) +
	( 16'sd 20160) * $signed(input_fmap_139[7:0]) +
	( 16'sd 32254) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18079) * $signed(input_fmap_141[7:0]) +
	( 16'sd 22456) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26543) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2829) * $signed(input_fmap_144[7:0]) +
	( 15'sd 11297) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18129) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_147[7:0]) +
	( 14'sd 5834) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15250) * $signed(input_fmap_149[7:0]) +
	( 16'sd 19832) * $signed(input_fmap_150[7:0]) +
	( 16'sd 20433) * $signed(input_fmap_151[7:0]) +
	( 15'sd 11886) * $signed(input_fmap_152[7:0]) +
	( 16'sd 16519) * $signed(input_fmap_153[7:0]) +
	( 11'sd 795) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20380) * $signed(input_fmap_155[7:0]) +
	( 15'sd 12531) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29753) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_158[7:0]) +
	( 14'sd 7013) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11304) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22849) * $signed(input_fmap_161[7:0]) +
	( 16'sd 30717) * $signed(input_fmap_162[7:0]) +
	( 16'sd 19898) * $signed(input_fmap_163[7:0]) +
	( 15'sd 15029) * $signed(input_fmap_164[7:0]) +
	( 16'sd 31457) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18217) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7988) * $signed(input_fmap_167[7:0]) +
	( 16'sd 23898) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21655) * $signed(input_fmap_169[7:0]) +
	( 11'sd 516) * $signed(input_fmap_170[7:0]) +
	( 16'sd 26125) * $signed(input_fmap_171[7:0]) +
	( 16'sd 32255) * $signed(input_fmap_172[7:0]) +
	( 16'sd 30195) * $signed(input_fmap_173[7:0]) +
	( 13'sd 3672) * $signed(input_fmap_174[7:0]) +
	( 15'sd 12692) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7174) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15414) * $signed(input_fmap_177[7:0]) +
	( 15'sd 12312) * $signed(input_fmap_178[7:0]) +
	( 14'sd 4370) * $signed(input_fmap_179[7:0]) +
	( 14'sd 5512) * $signed(input_fmap_180[7:0]) +
	( 16'sd 27852) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19375) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17405) * $signed(input_fmap_183[7:0]) +
	( 13'sd 3269) * $signed(input_fmap_184[7:0]) +
	( 16'sd 18870) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9378) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4645) * $signed(input_fmap_187[7:0]) +
	( 16'sd 21146) * $signed(input_fmap_188[7:0]) +
	( 16'sd 31778) * $signed(input_fmap_189[7:0]) +
	( 16'sd 22401) * $signed(input_fmap_190[7:0]) +
	( 16'sd 27424) * $signed(input_fmap_191[7:0]) +
	( 10'sd 324) * $signed(input_fmap_192[7:0]) +
	( 16'sd 18872) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26304) * $signed(input_fmap_194[7:0]) +
	( 16'sd 26439) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15760) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25283) * $signed(input_fmap_197[7:0]) +
	( 15'sd 8592) * $signed(input_fmap_198[7:0]) +
	( 16'sd 26285) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29131) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16945) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31610) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19158) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14092) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28224) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12749) * $signed(input_fmap_206[7:0]) +
	( 15'sd 8824) * $signed(input_fmap_207[7:0]) +
	( 16'sd 20425) * $signed(input_fmap_208[7:0]) +
	( 14'sd 4236) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1616) * $signed(input_fmap_210[7:0]) +
	( 16'sd 19840) * $signed(input_fmap_211[7:0]) +
	( 16'sd 31242) * $signed(input_fmap_212[7:0]) +
	( 16'sd 25265) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28322) * $signed(input_fmap_214[7:0]) +
	( 15'sd 13871) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4225) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30598) * $signed(input_fmap_217[7:0]) +
	( 15'sd 14759) * $signed(input_fmap_218[7:0]) +
	( 16'sd 23997) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25607) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15785) * $signed(input_fmap_221[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_222[7:0]) +
	( 14'sd 4827) * $signed(input_fmap_223[7:0]) +
	( 9'sd 179) * $signed(input_fmap_224[7:0]) +
	( 14'sd 7475) * $signed(input_fmap_225[7:0]) +
	( 16'sd 19527) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20971) * $signed(input_fmap_227[7:0]) +
	( 15'sd 14545) * $signed(input_fmap_228[7:0]) +
	( 15'sd 11754) * $signed(input_fmap_229[7:0]) +
	( 13'sd 3922) * $signed(input_fmap_230[7:0]) +
	( 16'sd 32467) * $signed(input_fmap_231[7:0]) +
	( 16'sd 30752) * $signed(input_fmap_232[7:0]) +
	( 16'sd 22157) * $signed(input_fmap_233[7:0]) +
	( 15'sd 11922) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22264) * $signed(input_fmap_235[7:0]) +
	( 16'sd 17656) * $signed(input_fmap_236[7:0]) +
	( 14'sd 7627) * $signed(input_fmap_237[7:0]) +
	( 16'sd 21298) * $signed(input_fmap_238[7:0]) +
	( 15'sd 14348) * $signed(input_fmap_239[7:0]) +
	( 16'sd 17554) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23382) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22473) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30873) * $signed(input_fmap_244[7:0]) +
	( 15'sd 12015) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28588) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_247[7:0]) +
	( 16'sd 27632) * $signed(input_fmap_248[7:0]) +
	( 16'sd 18107) * $signed(input_fmap_249[7:0]) +
	( 15'sd 10538) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19161) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30384) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27181) * $signed(input_fmap_253[7:0]) +
	( 16'sd 27039) * $signed(input_fmap_254[7:0]) +
	( 15'sd 13764) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_215;
assign conv_mac_215 = 
	( 16'sd 18033) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30738) * $signed(input_fmap_1[7:0]) +
	( 11'sd 892) * $signed(input_fmap_2[7:0]) +
	( 16'sd 23471) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_4[7:0]) +
	( 15'sd 16154) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21371) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19288) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7449) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5838) * $signed(input_fmap_9[7:0]) +
	( 16'sd 16598) * $signed(input_fmap_10[7:0]) +
	( 9'sd 149) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7878) * $signed(input_fmap_12[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1944) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15949) * $signed(input_fmap_15[7:0]) +
	( 16'sd 27514) * $signed(input_fmap_16[7:0]) +
	( 15'sd 15041) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21363) * $signed(input_fmap_18[7:0]) +
	( 12'sd 1765) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9110) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13716) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11731) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15821) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22646) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17896) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18634) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29662) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4638) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12970) * $signed(input_fmap_29[7:0]) +
	( 13'sd 4031) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18015) * $signed(input_fmap_31[7:0]) +
	( 16'sd 25600) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19941) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22019) * $signed(input_fmap_35[7:0]) +
	( 11'sd 629) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1273) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13215) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4547) * $signed(input_fmap_39[7:0]) +
	( 16'sd 22830) * $signed(input_fmap_40[7:0]) +
	( 16'sd 19820) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12655) * $signed(input_fmap_42[7:0]) +
	( 15'sd 14504) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15626) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28707) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31603) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20806) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19274) * $signed(input_fmap_49[7:0]) +
	( 15'sd 14656) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1421) * $signed(input_fmap_51[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_52[7:0]) +
	( 11'sd 535) * $signed(input_fmap_53[7:0]) +
	( 16'sd 31347) * $signed(input_fmap_54[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30729) * $signed(input_fmap_56[7:0]) +
	( 12'sd 1173) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10102) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7411) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18718) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31952) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17317) * $signed(input_fmap_62[7:0]) +
	( 16'sd 22088) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17605) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19279) * $signed(input_fmap_65[7:0]) +
	( 12'sd 1313) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5382) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4271) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1545) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11144) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7276) * $signed(input_fmap_71[7:0]) +
	( 16'sd 19143) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24223) * $signed(input_fmap_73[7:0]) +
	( 15'sd 12215) * $signed(input_fmap_74[7:0]) +
	( 11'sd 674) * $signed(input_fmap_75[7:0]) +
	( 16'sd 23684) * $signed(input_fmap_76[7:0]) +
	( 16'sd 31391) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24263) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29133) * $signed(input_fmap_80[7:0]) +
	( 16'sd 29378) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22891) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18118) * $signed(input_fmap_83[7:0]) +
	( 16'sd 17319) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6372) * $signed(input_fmap_85[7:0]) +
	( 16'sd 24722) * $signed(input_fmap_86[7:0]) +
	( 15'sd 10229) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1270) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12578) * $signed(input_fmap_89[7:0]) +
	( 14'sd 7037) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11516) * $signed(input_fmap_91[7:0]) +
	( 12'sd 1759) * $signed(input_fmap_92[7:0]) +
	( 10'sd 500) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28685) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18369) * $signed(input_fmap_95[7:0]) +
	( 15'sd 14600) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17986) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10587) * $signed(input_fmap_98[7:0]) +
	( 13'sd 3593) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32546) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23831) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16336) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10927) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24188) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21787) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5437) * $signed(input_fmap_106[7:0]) +
	( 8'sd 66) * $signed(input_fmap_107[7:0]) +
	( 15'sd 16244) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32426) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11636) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32605) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19209) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26943) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9015) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20125) * $signed(input_fmap_115[7:0]) +
	( 16'sd 28429) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16673) * $signed(input_fmap_117[7:0]) +
	( 16'sd 28631) * $signed(input_fmap_118[7:0]) +
	( 15'sd 9314) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15526) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19975) * $signed(input_fmap_121[7:0]) +
	( 13'sd 2624) * $signed(input_fmap_122[7:0]) +
	( 15'sd 16273) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20885) * $signed(input_fmap_125[7:0]) +
	( 5'sd 10) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30939) * $signed(input_fmap_127[7:0]) +
	( 16'sd 24528) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1157) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12499) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23899) * $signed(input_fmap_131[7:0]) +
	( 16'sd 32404) * $signed(input_fmap_132[7:0]) +
	( 15'sd 8895) * $signed(input_fmap_133[7:0]) +
	( 16'sd 16875) * $signed(input_fmap_134[7:0]) +
	( 16'sd 28597) * $signed(input_fmap_135[7:0]) +
	( 16'sd 27426) * $signed(input_fmap_136[7:0]) +
	( 15'sd 15185) * $signed(input_fmap_137[7:0]) +
	( 15'sd 8205) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8251) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30679) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3520) * $signed(input_fmap_141[7:0]) +
	( 16'sd 17392) * $signed(input_fmap_142[7:0]) +
	( 15'sd 10330) * $signed(input_fmap_143[7:0]) +
	( 14'sd 8133) * $signed(input_fmap_144[7:0]) +
	( 16'sd 31128) * $signed(input_fmap_145[7:0]) +
	( 16'sd 19875) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20124) * $signed(input_fmap_148[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_149[7:0]) +
	( 15'sd 15600) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28311) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14894) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23329) * $signed(input_fmap_153[7:0]) +
	( 15'sd 15048) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30503) * $signed(input_fmap_155[7:0]) +
	( 15'sd 14948) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11404) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20342) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2492) * $signed(input_fmap_159[7:0]) +
	( 13'sd 3570) * $signed(input_fmap_160[7:0]) +
	( 15'sd 12376) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14895) * $signed(input_fmap_162[7:0]) +
	( 16'sd 28738) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8682) * $signed(input_fmap_164[7:0]) +
	( 15'sd 14985) * $signed(input_fmap_165[7:0]) +
	( 16'sd 21179) * $signed(input_fmap_166[7:0]) +
	( 7'sd 53) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14342) * $signed(input_fmap_168[7:0]) +
	( 13'sd 3559) * $signed(input_fmap_169[7:0]) +
	( 12'sd 1809) * $signed(input_fmap_170[7:0]) +
	( 11'sd 810) * $signed(input_fmap_171[7:0]) +
	( 16'sd 16639) * $signed(input_fmap_172[7:0]) +
	( 16'sd 28571) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6521) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17170) * $signed(input_fmap_175[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_176[7:0]) +
	( 16'sd 26099) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_178[7:0]) +
	( 16'sd 26802) * $signed(input_fmap_179[7:0]) +
	( 15'sd 11852) * $signed(input_fmap_180[7:0]) +
	( 15'sd 14229) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4303) * $signed(input_fmap_182[7:0]) +
	( 11'sd 663) * $signed(input_fmap_183[7:0]) +
	( 12'sd 1201) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18846) * $signed(input_fmap_186[7:0]) +
	( 16'sd 24788) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29191) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20387) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14698) * $signed(input_fmap_191[7:0]) +
	( 14'sd 4393) * $signed(input_fmap_192[7:0]) +
	( 14'sd 8000) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18138) * $signed(input_fmap_194[7:0]) +
	( 15'sd 10199) * $signed(input_fmap_195[7:0]) +
	( 11'sd 668) * $signed(input_fmap_196[7:0]) +
	( 16'sd 17640) * $signed(input_fmap_197[7:0]) +
	( 15'sd 13222) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14985) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5114) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6184) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19284) * $signed(input_fmap_202[7:0]) +
	( 14'sd 4966) * $signed(input_fmap_203[7:0]) +
	( 16'sd 18524) * $signed(input_fmap_204[7:0]) +
	( 16'sd 17321) * $signed(input_fmap_205[7:0]) +
	( 16'sd 25439) * $signed(input_fmap_206[7:0]) +
	( 16'sd 19005) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4792) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11311) * $signed(input_fmap_209[7:0]) +
	( 15'sd 13930) * $signed(input_fmap_210[7:0]) +
	( 16'sd 25318) * $signed(input_fmap_211[7:0]) +
	( 16'sd 27339) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11537) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31638) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9008) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4918) * $signed(input_fmap_216[7:0]) +
	( 15'sd 8211) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30413) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5574) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19018) * $signed(input_fmap_220[7:0]) +
	( 13'sd 3200) * $signed(input_fmap_221[7:0]) +
	( 12'sd 1403) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24956) * $signed(input_fmap_223[7:0]) +
	( 16'sd 31250) * $signed(input_fmap_224[7:0]) +
	( 14'sd 6416) * $signed(input_fmap_225[7:0]) +
	( 8'sd 91) * $signed(input_fmap_226[7:0]) +
	( 16'sd 25187) * $signed(input_fmap_227[7:0]) +
	( 16'sd 29965) * $signed(input_fmap_228[7:0]) +
	( 10'sd 418) * $signed(input_fmap_229[7:0]) +
	( 16'sd 16475) * $signed(input_fmap_230[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29491) * $signed(input_fmap_232[7:0]) +
	( 14'sd 4188) * $signed(input_fmap_233[7:0]) +
	( 12'sd 1959) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19816) * $signed(input_fmap_235[7:0]) +
	( 15'sd 9885) * $signed(input_fmap_236[7:0]) +
	( 16'sd 31942) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3938) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20284) * $signed(input_fmap_239[7:0]) +
	( 15'sd 15332) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5917) * $signed(input_fmap_241[7:0]) +
	( 14'sd 7777) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7564) * $signed(input_fmap_243[7:0]) +
	( 16'sd 29390) * $signed(input_fmap_244[7:0]) +
	( 16'sd 26345) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9877) * $signed(input_fmap_246[7:0]) +
	( 14'sd 7543) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1592) * $signed(input_fmap_248[7:0]) +
	( 15'sd 8941) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32690) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_251[7:0]) +
	( 16'sd 28511) * $signed(input_fmap_252[7:0]) +
	( 16'sd 31759) * $signed(input_fmap_253[7:0]) +
	( 14'sd 7351) * $signed(input_fmap_254[7:0]) +
	( 16'sd 32210) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_216;
assign conv_mac_216 = 
	( 15'sd 11432) * $signed(input_fmap_0[7:0]) +
	( 14'sd 6516) * $signed(input_fmap_1[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25510) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3719) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30863) * $signed(input_fmap_6[7:0]) +
	( 16'sd 26234) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1771) * $signed(input_fmap_8[7:0]) +
	( 13'sd 4088) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9887) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9690) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1548) * $signed(input_fmap_13[7:0]) +
	( 16'sd 29638) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6179) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19989) * $signed(input_fmap_16[7:0]) +
	( 16'sd 16984) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29939) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_19[7:0]) +
	( 16'sd 24880) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3360) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6919) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7387) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30802) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21230) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21255) * $signed(input_fmap_26[7:0]) +
	( 14'sd 7873) * $signed(input_fmap_27[7:0]) +
	( 14'sd 7506) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13977) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26810) * $signed(input_fmap_30[7:0]) +
	( 16'sd 19177) * $signed(input_fmap_31[7:0]) +
	( 16'sd 32404) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27201) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3579) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16637) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32337) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19353) * $signed(input_fmap_37[7:0]) +
	( 16'sd 19881) * $signed(input_fmap_38[7:0]) +
	( 16'sd 31941) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20494) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11910) * $signed(input_fmap_41[7:0]) +
	( 16'sd 32480) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24978) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3872) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21011) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2443) * $signed(input_fmap_46[7:0]) +
	( 13'sd 2233) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3311) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18321) * $signed(input_fmap_49[7:0]) +
	( 13'sd 2622) * $signed(input_fmap_50[7:0]) +
	( 16'sd 22111) * $signed(input_fmap_51[7:0]) +
	( 14'sd 4151) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25719) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6234) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8848) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12667) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23660) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28335) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32345) * $signed(input_fmap_59[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16878) * $signed(input_fmap_61[7:0]) +
	( 16'sd 32613) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10636) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17819) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23024) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23323) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13802) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24068) * $signed(input_fmap_68[7:0]) +
	( 16'sd 28706) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22256) * $signed(input_fmap_70[7:0]) +
	( 16'sd 21728) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11620) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7101) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11840) * $signed(input_fmap_74[7:0]) +
	( 16'sd 22805) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13030) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18481) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13072) * $signed(input_fmap_78[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19055) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1180) * $signed(input_fmap_81[7:0]) +
	( 15'sd 11813) * $signed(input_fmap_82[7:0]) +
	( 15'sd 12664) * $signed(input_fmap_83[7:0]) +
	( 15'sd 8210) * $signed(input_fmap_84[7:0]) +
	( 15'sd 9484) * $signed(input_fmap_85[7:0]) +
	( 16'sd 17806) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31735) * $signed(input_fmap_87[7:0]) +
	( 16'sd 16935) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29516) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3196) * $signed(input_fmap_90[7:0]) +
	( 16'sd 32058) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20769) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17297) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23057) * $signed(input_fmap_94[7:0]) +
	( 11'sd 723) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1547) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7822) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4601) * $signed(input_fmap_98[7:0]) +
	( 8'sd 107) * $signed(input_fmap_99[7:0]) +
	( 16'sd 22348) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31122) * $signed(input_fmap_101[7:0]) +
	( 14'sd 7154) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8272) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25958) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6378) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6965) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2974) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32474) * $signed(input_fmap_108[7:0]) +
	( 16'sd 20887) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3555) * $signed(input_fmap_110[7:0]) +
	( 15'sd 10577) * $signed(input_fmap_111[7:0]) +
	( 15'sd 8490) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4495) * $signed(input_fmap_113[7:0]) +
	( 16'sd 18785) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2124) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13139) * $signed(input_fmap_117[7:0]) +
	( 16'sd 31008) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24146) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15912) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1652) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3815) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30366) * $signed(input_fmap_123[7:0]) +
	( 15'sd 13005) * $signed(input_fmap_124[7:0]) +
	( 16'sd 31881) * $signed(input_fmap_125[7:0]) +
	( 15'sd 13946) * $signed(input_fmap_126[7:0]) +
	( 12'sd 1779) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13881) * $signed(input_fmap_128[7:0]) +
	( 11'sd 572) * $signed(input_fmap_129[7:0]) +
	( 16'sd 26802) * $signed(input_fmap_130[7:0]) +
	( 15'sd 12482) * $signed(input_fmap_131[7:0]) +
	( 13'sd 3700) * $signed(input_fmap_132[7:0]) +
	( 16'sd 20174) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31344) * $signed(input_fmap_134[7:0]) +
	( 16'sd 22177) * $signed(input_fmap_135[7:0]) +
	( 11'sd 876) * $signed(input_fmap_136[7:0]) +
	( 15'sd 14161) * $signed(input_fmap_137[7:0]) +
	( 16'sd 30923) * $signed(input_fmap_138[7:0]) +
	( 16'sd 26107) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30581) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24784) * $signed(input_fmap_141[7:0]) +
	( 13'sd 3056) * $signed(input_fmap_142[7:0]) +
	( 13'sd 2969) * $signed(input_fmap_143[7:0]) +
	( 13'sd 3982) * $signed(input_fmap_144[7:0]) +
	( 15'sd 13995) * $signed(input_fmap_145[7:0]) +
	( 16'sd 28651) * $signed(input_fmap_146[7:0]) +
	( 15'sd 12447) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26155) * $signed(input_fmap_148[7:0]) +
	( 15'sd 11805) * $signed(input_fmap_149[7:0]) +
	( 16'sd 26101) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28135) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2565) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1110) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6023) * $signed(input_fmap_154[7:0]) +
	( 16'sd 17185) * $signed(input_fmap_155[7:0]) +
	( 14'sd 5480) * $signed(input_fmap_156[7:0]) +
	( 13'sd 3765) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11423) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2270) * $signed(input_fmap_159[7:0]) +
	( 12'sd 1414) * $signed(input_fmap_160[7:0]) +
	( 15'sd 15880) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2892) * $signed(input_fmap_162[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3203) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2249) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_166[7:0]) +
	( 16'sd 28694) * $signed(input_fmap_167[7:0]) +
	( 15'sd 8271) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27685) * $signed(input_fmap_169[7:0]) +
	( 10'sd 478) * $signed(input_fmap_170[7:0]) +
	( 16'sd 24016) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3120) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23188) * $signed(input_fmap_173[7:0]) +
	( 16'sd 29177) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1057) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20719) * $signed(input_fmap_176[7:0]) +
	( 14'sd 5899) * $signed(input_fmap_177[7:0]) +
	( 16'sd 19375) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2344) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29854) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25772) * $signed(input_fmap_181[7:0]) +
	( 10'sd 350) * $signed(input_fmap_182[7:0]) +
	( 16'sd 30601) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26397) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1630) * $signed(input_fmap_185[7:0]) +
	( 16'sd 30985) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4374) * $signed(input_fmap_187[7:0]) +
	( 16'sd 24776) * $signed(input_fmap_188[7:0]) +
	( 16'sd 29946) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30445) * $signed(input_fmap_190[7:0]) +
	( 16'sd 18864) * $signed(input_fmap_191[7:0]) +
	( 11'sd 780) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20329) * $signed(input_fmap_193[7:0]) +
	( 15'sd 12536) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17876) * $signed(input_fmap_195[7:0]) +
	( 16'sd 20287) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5369) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2710) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10910) * $signed(input_fmap_199[7:0]) +
	( 10'sd 299) * $signed(input_fmap_200[7:0]) +
	( 8'sd 93) * $signed(input_fmap_201[7:0]) +
	( 16'sd 32636) * $signed(input_fmap_202[7:0]) +
	( 16'sd 26305) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14932) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31411) * $signed(input_fmap_205[7:0]) +
	( 15'sd 11216) * $signed(input_fmap_206[7:0]) +
	( 16'sd 17988) * $signed(input_fmap_207[7:0]) +
	( 16'sd 21443) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11547) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18262) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28315) * $signed(input_fmap_211[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5206) * $signed(input_fmap_213[7:0]) +
	( 13'sd 2385) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9670) * $signed(input_fmap_215[7:0]) +
	( 16'sd 21168) * $signed(input_fmap_216[7:0]) +
	( 14'sd 7143) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21380) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10258) * $signed(input_fmap_219[7:0]) +
	( 16'sd 26080) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25808) * $signed(input_fmap_221[7:0]) +
	( 16'sd 22161) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28822) * $signed(input_fmap_223[7:0]) +
	( 16'sd 31974) * $signed(input_fmap_224[7:0]) +
	( 16'sd 30076) * $signed(input_fmap_225[7:0]) +
	( 16'sd 17641) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2484) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31202) * $signed(input_fmap_228[7:0]) +
	( 13'sd 2887) * $signed(input_fmap_229[7:0]) +
	( 16'sd 22573) * $signed(input_fmap_230[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_231[7:0]) +
	( 16'sd 23670) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10977) * $signed(input_fmap_233[7:0]) +
	( 16'sd 31030) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7978) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27918) * $signed(input_fmap_236[7:0]) +
	( 14'sd 4623) * $signed(input_fmap_237[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_238[7:0]) +
	( 11'sd 517) * $signed(input_fmap_239[7:0]) +
	( 11'sd 904) * $signed(input_fmap_240[7:0]) +
	( 16'sd 22804) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29318) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2081) * $signed(input_fmap_243[7:0]) +
	( 16'sd 16603) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19053) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1268) * $signed(input_fmap_246[7:0]) +
	( 14'sd 8067) * $signed(input_fmap_247[7:0]) +
	( 16'sd 31341) * $signed(input_fmap_248[7:0]) +
	( 16'sd 29531) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25520) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6688) * $signed(input_fmap_251[7:0]) +
	( 16'sd 21855) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17270) * $signed(input_fmap_253[7:0]) +
	( 16'sd 32239) * $signed(input_fmap_254[7:0]) +
	( 16'sd 29281) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_217;
assign conv_mac_217 = 
	( 13'sd 2340) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19934) * $signed(input_fmap_1[7:0]) +
	( 16'sd 16506) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6982) * $signed(input_fmap_3[7:0]) +
	( 15'sd 16247) * $signed(input_fmap_4[7:0]) +
	( 16'sd 32003) * $signed(input_fmap_5[7:0]) +
	( 15'sd 11091) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14344) * $signed(input_fmap_7[7:0]) +
	( 16'sd 22527) * $signed(input_fmap_8[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28414) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29836) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8602) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20271) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12886) * $signed(input_fmap_14[7:0]) +
	( 15'sd 16217) * $signed(input_fmap_15[7:0]) +
	( 16'sd 24531) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29392) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6374) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9182) * $signed(input_fmap_20[7:0]) +
	( 14'sd 6669) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5778) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11996) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7808) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31458) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15532) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22070) * $signed(input_fmap_27[7:0]) +
	( 14'sd 8151) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9340) * $signed(input_fmap_29[7:0]) +
	( 10'sd 379) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24418) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29778) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10431) * $signed(input_fmap_33[7:0]) +
	( 15'sd 12071) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32321) * $signed(input_fmap_35[7:0]) +
	( 16'sd 17078) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29509) * $signed(input_fmap_37[7:0]) +
	( 16'sd 27504) * $signed(input_fmap_38[7:0]) +
	( 15'sd 10581) * $signed(input_fmap_39[7:0]) +
	( 16'sd 32077) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18944) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26200) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18907) * $signed(input_fmap_43[7:0]) +
	( 16'sd 18213) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15861) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23495) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8003) * $signed(input_fmap_47[7:0]) +
	( 15'sd 9347) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24070) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20809) * $signed(input_fmap_50[7:0]) +
	( 16'sd 20078) * $signed(input_fmap_51[7:0]) +
	( 16'sd 27852) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24859) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12440) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20190) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25378) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17560) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25197) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7131) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12367) * $signed(input_fmap_61[7:0]) +
	( 15'sd 15383) * $signed(input_fmap_62[7:0]) +
	( 14'sd 8102) * $signed(input_fmap_63[7:0]) +
	( 16'sd 23868) * $signed(input_fmap_64[7:0]) +
	( 14'sd 8089) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14536) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24917) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11054) * $signed(input_fmap_68[7:0]) +
	( 14'sd 6369) * $signed(input_fmap_69[7:0]) +
	( 15'sd 11227) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3539) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23868) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1562) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5241) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14684) * $signed(input_fmap_75[7:0]) +
	( 14'sd 6894) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21245) * $signed(input_fmap_78[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_79[7:0]) +
	( 15'sd 14129) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25551) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_82[7:0]) +
	( 16'sd 29725) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16380) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1906) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14486) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8419) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22751) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1557) * $signed(input_fmap_89[7:0]) +
	( 12'sd 1619) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17947) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19523) * $signed(input_fmap_92[7:0]) +
	( 16'sd 28853) * $signed(input_fmap_93[7:0]) +
	( 14'sd 6486) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10976) * $signed(input_fmap_95[7:0]) +
	( 16'sd 27170) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18614) * $signed(input_fmap_97[7:0]) +
	( 16'sd 20346) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24733) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6784) * $signed(input_fmap_101[7:0]) +
	( 6'sd 22) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_103[7:0]) +
	( 16'sd 23376) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15266) * $signed(input_fmap_105[7:0]) +
	( 14'sd 5514) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14090) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28934) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32740) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19070) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1565) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3302) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22515) * $signed(input_fmap_113[7:0]) +
	( 16'sd 20236) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15619) * $signed(input_fmap_115[7:0]) +
	( 15'sd 15975) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6534) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4967) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22683) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20444) * $signed(input_fmap_120[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28171) * $signed(input_fmap_122[7:0]) +
	( 14'sd 7107) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5859) * $signed(input_fmap_124[7:0]) +
	( 13'sd 3600) * $signed(input_fmap_125[7:0]) +
	( 16'sd 23020) * $signed(input_fmap_126[7:0]) +
	( 16'sd 20933) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13957) * $signed(input_fmap_128[7:0]) +
	( 14'sd 6824) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31950) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14767) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1702) * $signed(input_fmap_132[7:0]) +
	( 15'sd 13974) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3903) * $signed(input_fmap_134[7:0]) +
	( 16'sd 20241) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1471) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13344) * $signed(input_fmap_137[7:0]) +
	( 9'sd 241) * $signed(input_fmap_138[7:0]) +
	( 16'sd 24151) * $signed(input_fmap_139[7:0]) +
	( 13'sd 3498) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29087) * $signed(input_fmap_141[7:0]) +
	( 12'sd 1556) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1724) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_144[7:0]) +
	( 11'sd 908) * $signed(input_fmap_145[7:0]) +
	( 16'sd 31511) * $signed(input_fmap_146[7:0]) +
	( 13'sd 2545) * $signed(input_fmap_147[7:0]) +
	( 13'sd 3709) * $signed(input_fmap_148[7:0]) +
	( 15'sd 9674) * $signed(input_fmap_149[7:0]) +
	( 15'sd 14016) * $signed(input_fmap_150[7:0]) +
	( 16'sd 28369) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30732) * $signed(input_fmap_152[7:0]) +
	( 16'sd 20163) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11756) * $signed(input_fmap_154[7:0]) +
	( 15'sd 9706) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20980) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29740) * $signed(input_fmap_157[7:0]) +
	( 14'sd 6221) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2759) * $signed(input_fmap_159[7:0]) +
	( 15'sd 11401) * $signed(input_fmap_160[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_161[7:0]) +
	( 16'sd 28059) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3919) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1078) * $signed(input_fmap_164[7:0]) +
	( 16'sd 30217) * $signed(input_fmap_165[7:0]) +
	( 9'sd 188) * $signed(input_fmap_166[7:0]) +
	( 16'sd 23321) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1956) * $signed(input_fmap_168[7:0]) +
	( 16'sd 19022) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11698) * $signed(input_fmap_170[7:0]) +
	( 16'sd 28803) * $signed(input_fmap_171[7:0]) +
	( 15'sd 8284) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1729) * $signed(input_fmap_173[7:0]) +
	( 16'sd 29757) * $signed(input_fmap_174[7:0]) +
	( 16'sd 16745) * $signed(input_fmap_175[7:0]) +
	( 15'sd 16377) * $signed(input_fmap_176[7:0]) +
	( 16'sd 28830) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14190) * $signed(input_fmap_178[7:0]) +
	( 16'sd 20996) * $signed(input_fmap_179[7:0]) +
	( 6'sd 22) * $signed(input_fmap_180[7:0]) +
	( 13'sd 2545) * $signed(input_fmap_181[7:0]) +
	( 16'sd 31687) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17382) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14960) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6577) * $signed(input_fmap_185[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_186[7:0]) +
	( 16'sd 30437) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17120) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2063) * $signed(input_fmap_189[7:0]) +
	( 13'sd 3261) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26301) * $signed(input_fmap_191[7:0]) +
	( 13'sd 2409) * $signed(input_fmap_192[7:0]) +
	( 15'sd 10753) * $signed(input_fmap_193[7:0]) +
	( 12'sd 1779) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1470) * $signed(input_fmap_195[7:0]) +
	( 15'sd 13192) * $signed(input_fmap_196[7:0]) +
	( 15'sd 13423) * $signed(input_fmap_197[7:0]) +
	( 14'sd 7233) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23395) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13290) * $signed(input_fmap_200[7:0]) +
	( 16'sd 25219) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31203) * $signed(input_fmap_202[7:0]) +
	( 13'sd 4083) * $signed(input_fmap_203[7:0]) +
	( 15'sd 9249) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18682) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_206[7:0]) +
	( 16'sd 22024) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15182) * $signed(input_fmap_208[7:0]) +
	( 16'sd 22458) * $signed(input_fmap_209[7:0]) +
	( 14'sd 7217) * $signed(input_fmap_210[7:0]) +
	( 16'sd 22130) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29685) * $signed(input_fmap_212[7:0]) +
	( 16'sd 27820) * $signed(input_fmap_213[7:0]) +
	( 16'sd 29462) * $signed(input_fmap_214[7:0]) +
	( 15'sd 15179) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4563) * $signed(input_fmap_216[7:0]) +
	( 16'sd 16777) * $signed(input_fmap_217[7:0]) +
	( 16'sd 21370) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19910) * $signed(input_fmap_219[7:0]) +
	( 16'sd 17568) * $signed(input_fmap_220[7:0]) +
	( 11'sd 961) * $signed(input_fmap_221[7:0]) +
	( 16'sd 20016) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12753) * $signed(input_fmap_223[7:0]) +
	( 15'sd 9980) * $signed(input_fmap_224[7:0]) +
	( 15'sd 10481) * $signed(input_fmap_225[7:0]) +
	( 16'sd 28729) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13203) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_228[7:0]) +
	( 16'sd 26049) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29786) * $signed(input_fmap_230[7:0]) +
	( 15'sd 11859) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9705) * $signed(input_fmap_232[7:0]) +
	( 13'sd 2875) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4801) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7053) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27999) * $signed(input_fmap_236[7:0]) +
	( 16'sd 25736) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27911) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31274) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10026) * $signed(input_fmap_240[7:0]) +
	( 14'sd 4443) * $signed(input_fmap_241[7:0]) +
	( 13'sd 2437) * $signed(input_fmap_242[7:0]) +
	( 16'sd 31903) * $signed(input_fmap_243[7:0]) +
	( 14'sd 4868) * $signed(input_fmap_244[7:0]) +
	( 15'sd 9266) * $signed(input_fmap_245[7:0]) +
	( 13'sd 3444) * $signed(input_fmap_246[7:0]) +
	( 15'sd 16051) * $signed(input_fmap_247[7:0]) +
	( 12'sd 1578) * $signed(input_fmap_248[7:0]) +
	( 16'sd 23956) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22077) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15547) * $signed(input_fmap_251[7:0]) +
	( 11'sd 873) * $signed(input_fmap_252[7:0]) +
	( 15'sd 14599) * $signed(input_fmap_253[7:0]) +
	( 15'sd 10939) * $signed(input_fmap_254[7:0]) +
	( 14'sd 7562) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_218;
assign conv_mac_218 = 
	( 14'sd 7414) * $signed(input_fmap_0[7:0]) +
	( 15'sd 15037) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3807) * $signed(input_fmap_2[7:0]) +
	( 16'sd 22245) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_4[7:0]) +
	( 16'sd 20948) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9125) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3307) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4923) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6367) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21306) * $signed(input_fmap_10[7:0]) +
	( 12'sd 1683) * $signed(input_fmap_11[7:0]) +
	( 16'sd 18236) * $signed(input_fmap_12[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17940) * $signed(input_fmap_14[7:0]) +
	( 15'sd 8827) * $signed(input_fmap_15[7:0]) +
	( 15'sd 15579) * $signed(input_fmap_16[7:0]) +
	( 16'sd 31402) * $signed(input_fmap_17[7:0]) +
	( 16'sd 21901) * $signed(input_fmap_18[7:0]) +
	( 16'sd 30589) * $signed(input_fmap_19[7:0]) +
	( 13'sd 3284) * $signed(input_fmap_20[7:0]) +
	( 16'sd 27442) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7833) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14810) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25159) * $signed(input_fmap_24[7:0]) +
	( 15'sd 10303) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28268) * $signed(input_fmap_26[7:0]) +
	( 15'sd 11261) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30598) * $signed(input_fmap_28[7:0]) +
	( 13'sd 2786) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31644) * $signed(input_fmap_30[7:0]) +
	( 15'sd 14591) * $signed(input_fmap_31[7:0]) +
	( 16'sd 27818) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24737) * $signed(input_fmap_33[7:0]) +
	( 15'sd 13701) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16972) * $signed(input_fmap_35[7:0]) +
	( 14'sd 8151) * $signed(input_fmap_36[7:0]) +
	( 16'sd 17625) * $signed(input_fmap_37[7:0]) +
	( 11'sd 797) * $signed(input_fmap_38[7:0]) +
	( 15'sd 16253) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_40[7:0]) +
	( 15'sd 10438) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9637) * $signed(input_fmap_42[7:0]) +
	( 14'sd 7082) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13322) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14788) * $signed(input_fmap_45[7:0]) +
	( 16'sd 27316) * $signed(input_fmap_46[7:0]) +
	( 9'sd 225) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19606) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23069) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27785) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29000) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14448) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25016) * $signed(input_fmap_53[7:0]) +
	( 15'sd 8963) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25144) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_56[7:0]) +
	( 15'sd 15296) * $signed(input_fmap_57[7:0]) +
	( 16'sd 30299) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17359) * $signed(input_fmap_59[7:0]) +
	( 16'sd 32248) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27026) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28332) * $signed(input_fmap_62[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17288) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12178) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6663) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17159) * $signed(input_fmap_67[7:0]) +
	( 15'sd 15891) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2741) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19265) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2527) * $signed(input_fmap_71[7:0]) +
	( 16'sd 24916) * $signed(input_fmap_72[7:0]) +
	( 15'sd 12245) * $signed(input_fmap_73[7:0]) +
	( 16'sd 24387) * $signed(input_fmap_74[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20721) * $signed(input_fmap_76[7:0]) +
	( 14'sd 6536) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18403) * $signed(input_fmap_78[7:0]) +
	( 15'sd 9388) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13583) * $signed(input_fmap_80[7:0]) +
	( 16'sd 27502) * $signed(input_fmap_81[7:0]) +
	( 14'sd 5306) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21152) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5993) * $signed(input_fmap_84[7:0]) +
	( 16'sd 16521) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29806) * $signed(input_fmap_86[7:0]) +
	( 16'sd 20026) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25500) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20797) * $signed(input_fmap_89[7:0]) +
	( 16'sd 19011) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31596) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24556) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30374) * $signed(input_fmap_93[7:0]) +
	( 16'sd 17158) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20895) * $signed(input_fmap_95[7:0]) +
	( 14'sd 7781) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27253) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3165) * $signed(input_fmap_98[7:0]) +
	( 14'sd 4822) * $signed(input_fmap_99[7:0]) +
	( 11'sd 1008) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3913) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12894) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6034) * $signed(input_fmap_103[7:0]) +
	( 14'sd 4157) * $signed(input_fmap_104[7:0]) +
	( 16'sd 16597) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21376) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25802) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10535) * $signed(input_fmap_108[7:0]) +
	( 16'sd 22365) * $signed(input_fmap_109[7:0]) +
	( 16'sd 28493) * $signed(input_fmap_110[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_111[7:0]) +
	( 16'sd 26419) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15449) * $signed(input_fmap_113[7:0]) +
	( 10'sd 466) * $signed(input_fmap_114[7:0]) +
	( 14'sd 6571) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26014) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26286) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29178) * $signed(input_fmap_118[7:0]) +
	( 15'sd 11857) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11039) * $signed(input_fmap_120[7:0]) +
	( 16'sd 31687) * $signed(input_fmap_121[7:0]) +
	( 10'sd 408) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12470) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12338) * $signed(input_fmap_124[7:0]) +
	( 15'sd 14887) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12695) * $signed(input_fmap_126[7:0]) +
	( 15'sd 9722) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9641) * $signed(input_fmap_128[7:0]) +
	( 15'sd 10413) * $signed(input_fmap_129[7:0]) +
	( 12'sd 1686) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_131[7:0]) +
	( 14'sd 6575) * $signed(input_fmap_132[7:0]) +
	( 16'sd 23623) * $signed(input_fmap_133[7:0]) +
	( 16'sd 26912) * $signed(input_fmap_134[7:0]) +
	( 15'sd 14165) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21408) * $signed(input_fmap_136[7:0]) +
	( 15'sd 8885) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27321) * $signed(input_fmap_138[7:0]) +
	( 16'sd 18066) * $signed(input_fmap_139[7:0]) +
	( 16'sd 29524) * $signed(input_fmap_140[7:0]) +
	( 16'sd 16419) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8305) * $signed(input_fmap_142[7:0]) +
	( 16'sd 27404) * $signed(input_fmap_143[7:0]) +
	( 14'sd 7315) * $signed(input_fmap_144[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_145[7:0]) +
	( 16'sd 22684) * $signed(input_fmap_146[7:0]) +
	( 16'sd 27498) * $signed(input_fmap_147[7:0]) +
	( 15'sd 14803) * $signed(input_fmap_148[7:0]) +
	( 12'sd 1818) * $signed(input_fmap_149[7:0]) +
	( 15'sd 11271) * $signed(input_fmap_150[7:0]) +
	( 16'sd 32363) * $signed(input_fmap_151[7:0]) +
	( 16'sd 32179) * $signed(input_fmap_152[7:0]) +
	( 15'sd 9780) * $signed(input_fmap_153[7:0]) +
	( 12'sd 1694) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19210) * $signed(input_fmap_155[7:0]) +
	( 16'sd 24317) * $signed(input_fmap_156[7:0]) +
	( 16'sd 20530) * $signed(input_fmap_157[7:0]) +
	( 15'sd 13491) * $signed(input_fmap_158[7:0]) +
	( 16'sd 25941) * $signed(input_fmap_159[7:0]) +
	( 10'sd 328) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19400) * $signed(input_fmap_161[7:0]) +
	( 15'sd 8852) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26942) * $signed(input_fmap_163[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_164[7:0]) +
	( 13'sd 4068) * $signed(input_fmap_165[7:0]) +
	( 16'sd 27247) * $signed(input_fmap_166[7:0]) +
	( 15'sd 12132) * $signed(input_fmap_167[7:0]) +
	( 14'sd 7639) * $signed(input_fmap_168[7:0]) +
	( 15'sd 14843) * $signed(input_fmap_169[7:0]) +
	( 15'sd 10734) * $signed(input_fmap_170[7:0]) +
	( 16'sd 22409) * $signed(input_fmap_171[7:0]) +
	( 11'sd 595) * $signed(input_fmap_172[7:0]) +
	( 16'sd 26822) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14736) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7670) * $signed(input_fmap_175[7:0]) +
	( 11'sd 968) * $signed(input_fmap_176[7:0]) +
	( 15'sd 8432) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22915) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25017) * $signed(input_fmap_179[7:0]) +
	( 14'sd 7479) * $signed(input_fmap_180[7:0]) +
	( 11'sd 564) * $signed(input_fmap_181[7:0]) +
	( 16'sd 32604) * $signed(input_fmap_182[7:0]) +
	( 14'sd 5085) * $signed(input_fmap_183[7:0]) +
	( 16'sd 30385) * $signed(input_fmap_184[7:0]) +
	( 15'sd 16163) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_186[7:0]) +
	( 16'sd 27186) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4952) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30897) * $signed(input_fmap_189[7:0]) +
	( 16'sd 24187) * $signed(input_fmap_190[7:0]) +
	( 16'sd 25607) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22433) * $signed(input_fmap_192[7:0]) +
	( 14'sd 6584) * $signed(input_fmap_193[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_194[7:0]) +
	( 16'sd 20170) * $signed(input_fmap_195[7:0]) +
	( 16'sd 29928) * $signed(input_fmap_196[7:0]) +
	( 16'sd 23047) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9695) * $signed(input_fmap_198[7:0]) +
	( 16'sd 32732) * $signed(input_fmap_199[7:0]) +
	( 16'sd 24171) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22514) * $signed(input_fmap_201[7:0]) +
	( 16'sd 16739) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19098) * $signed(input_fmap_203[7:0]) +
	( 15'sd 10723) * $signed(input_fmap_204[7:0]) +
	( 15'sd 14432) * $signed(input_fmap_205[7:0]) +
	( 14'sd 6139) * $signed(input_fmap_206[7:0]) +
	( 16'sd 20726) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8542) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3443) * $signed(input_fmap_209[7:0]) +
	( 14'sd 8091) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26149) * $signed(input_fmap_211[7:0]) +
	( 15'sd 8608) * $signed(input_fmap_212[7:0]) +
	( 15'sd 14698) * $signed(input_fmap_213[7:0]) +
	( 15'sd 14081) * $signed(input_fmap_214[7:0]) +
	( 16'sd 24470) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18911) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9133) * $signed(input_fmap_217[7:0]) +
	( 15'sd 16081) * $signed(input_fmap_218[7:0]) +
	( 15'sd 13198) * $signed(input_fmap_219[7:0]) +
	( 13'sd 3500) * $signed(input_fmap_220[7:0]) +
	( 13'sd 2316) * $signed(input_fmap_221[7:0]) +
	( 16'sd 26329) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28477) * $signed(input_fmap_223[7:0]) +
	( 16'sd 19013) * $signed(input_fmap_224[7:0]) +
	( 16'sd 29865) * $signed(input_fmap_225[7:0]) +
	( 15'sd 13620) * $signed(input_fmap_226[7:0]) +
	( 12'sd 1396) * $signed(input_fmap_227[7:0]) +
	( 15'sd 8445) * $signed(input_fmap_228[7:0]) +
	( 16'sd 18826) * $signed(input_fmap_229[7:0]) +
	( 16'sd 23304) * $signed(input_fmap_230[7:0]) +
	( 16'sd 22938) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_232[7:0]) +
	( 15'sd 12306) * $signed(input_fmap_233[7:0]) +
	( 16'sd 16446) * $signed(input_fmap_234[7:0]) +
	( 16'sd 17625) * $signed(input_fmap_235[7:0]) +
	( 16'sd 26814) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2911) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28095) * $signed(input_fmap_238[7:0]) +
	( 14'sd 6704) * $signed(input_fmap_239[7:0]) +
	( 16'sd 28676) * $signed(input_fmap_240[7:0]) +
	( 16'sd 28417) * $signed(input_fmap_241[7:0]) +
	( 16'sd 16656) * $signed(input_fmap_242[7:0]) +
	( 16'sd 18589) * $signed(input_fmap_243[7:0]) +
	( 15'sd 15864) * $signed(input_fmap_244[7:0]) +
	( 14'sd 7504) * $signed(input_fmap_245[7:0]) +
	( 13'sd 2061) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21670) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15262) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3173) * $signed(input_fmap_250[7:0]) +
	( 15'sd 10826) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26732) * $signed(input_fmap_252[7:0]) +
	( 16'sd 22696) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2435) * $signed(input_fmap_254[7:0]) +
	( 16'sd 29683) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_219;
assign conv_mac_219 = 
	( 14'sd 5437) * $signed(input_fmap_0[7:0]) +
	( 15'sd 11791) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2447) * $signed(input_fmap_2[7:0]) +
	( 14'sd 4608) * $signed(input_fmap_3[7:0]) +
	( 15'sd 15772) * $signed(input_fmap_4[7:0]) +
	( 16'sd 25989) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1425) * $signed(input_fmap_6[7:0]) +
	( 13'sd 3271) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12810) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15745) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9559) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26554) * $signed(input_fmap_11[7:0]) +
	( 16'sd 17725) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15862) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15866) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22487) * $signed(input_fmap_15[7:0]) +
	( 14'sd 6004) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21392) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4318) * $signed(input_fmap_18[7:0]) +
	( 16'sd 22301) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23546) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26334) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23120) * $signed(input_fmap_22[7:0]) +
	( 16'sd 19457) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7440) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31835) * $signed(input_fmap_25[7:0]) +
	( 16'sd 17395) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9125) * $signed(input_fmap_27[7:0]) +
	( 16'sd 27991) * $signed(input_fmap_28[7:0]) +
	( 14'sd 4419) * $signed(input_fmap_29[7:0]) +
	( 16'sd 27409) * $signed(input_fmap_30[7:0]) +
	( 13'sd 2609) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18356) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13880) * $signed(input_fmap_33[7:0]) +
	( 16'sd 27234) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13496) * $signed(input_fmap_35[7:0]) +
	( 15'sd 8245) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11221) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24224) * $signed(input_fmap_38[7:0]) +
	( 16'sd 26341) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20989) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24347) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23045) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10647) * $signed(input_fmap_43[7:0]) +
	( 14'sd 4809) * $signed(input_fmap_44[7:0]) +
	( 16'sd 24874) * $signed(input_fmap_45[7:0]) +
	( 16'sd 31795) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26700) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30330) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5178) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27538) * $signed(input_fmap_50[7:0]) +
	( 16'sd 24675) * $signed(input_fmap_51[7:0]) +
	( 16'sd 30365) * $signed(input_fmap_52[7:0]) +
	( 11'sd 1019) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29729) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17932) * $signed(input_fmap_55[7:0]) +
	( 16'sd 30437) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6506) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10773) * $signed(input_fmap_58[7:0]) +
	( 10'sd 491) * $signed(input_fmap_59[7:0]) +
	( 16'sd 18503) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27256) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2435) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12083) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24327) * $signed(input_fmap_64[7:0]) +
	( 16'sd 24487) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32675) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14939) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29842) * $signed(input_fmap_68[7:0]) +
	( 9'sd 207) * $signed(input_fmap_69[7:0]) +
	( 16'sd 25110) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16025) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11303) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11341) * $signed(input_fmap_73[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23170) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19480) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19689) * $signed(input_fmap_77[7:0]) +
	( 16'sd 30466) * $signed(input_fmap_78[7:0]) +
	( 15'sd 8412) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30051) * $signed(input_fmap_80[7:0]) +
	( 10'sd 303) * $signed(input_fmap_81[7:0]) +
	( 15'sd 13150) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9137) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2231) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18635) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28694) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19653) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16107) * $signed(input_fmap_88[7:0]) +
	( 12'sd 1489) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12406) * $signed(input_fmap_90[7:0]) +
	( 12'sd 1525) * $signed(input_fmap_91[7:0]) +
	( 16'sd 25956) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26078) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13736) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23431) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20870) * $signed(input_fmap_96[7:0]) +
	( 13'sd 3824) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9645) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29047) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31624) * $signed(input_fmap_100[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16415) * $signed(input_fmap_102[7:0]) +
	( 13'sd 2084) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27494) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26671) * $signed(input_fmap_105[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11661) * $signed(input_fmap_107[7:0]) +
	( 14'sd 7416) * $signed(input_fmap_108[7:0]) +
	( 15'sd 12434) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29729) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17250) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13736) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19880) * $signed(input_fmap_113[7:0]) +
	( 16'sd 25283) * $signed(input_fmap_114[7:0]) +
	( 14'sd 8054) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9120) * $signed(input_fmap_116[7:0]) +
	( 11'sd 802) * $signed(input_fmap_117[7:0]) +
	( 15'sd 11258) * $signed(input_fmap_118[7:0]) +
	( 14'sd 6527) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9037) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25678) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11086) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21991) * $signed(input_fmap_124[7:0]) +
	( 15'sd 12981) * $signed(input_fmap_125[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10235) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2071) * $signed(input_fmap_128[7:0]) +
	( 11'sd 895) * $signed(input_fmap_129[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_130[7:0]) +
	( 16'sd 27317) * $signed(input_fmap_131[7:0]) +
	( 16'sd 19974) * $signed(input_fmap_132[7:0]) +
	( 11'sd 665) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1478) * $signed(input_fmap_134[7:0]) +
	( 16'sd 24250) * $signed(input_fmap_135[7:0]) +
	( 16'sd 27693) * $signed(input_fmap_136[7:0]) +
	( 13'sd 2709) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11680) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27146) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17847) * $signed(input_fmap_140[7:0]) +
	( 13'sd 4039) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11553) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20978) * $signed(input_fmap_143[7:0]) +
	( 12'sd 1534) * $signed(input_fmap_144[7:0]) +
	( 13'sd 2797) * $signed(input_fmap_145[7:0]) +
	( 16'sd 18699) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17875) * $signed(input_fmap_147[7:0]) +
	( 16'sd 19213) * $signed(input_fmap_148[7:0]) +
	( 15'sd 13158) * $signed(input_fmap_149[7:0]) +
	( 16'sd 29190) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24687) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21025) * $signed(input_fmap_152[7:0]) +
	( 16'sd 27468) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23831) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_155[7:0]) +
	( 16'sd 27860) * $signed(input_fmap_156[7:0]) +
	( 16'sd 21296) * $signed(input_fmap_157[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_158[7:0]) +
	( 16'sd 29075) * $signed(input_fmap_159[7:0]) +
	( 15'sd 10741) * $signed(input_fmap_160[7:0]) +
	( 16'sd 28964) * $signed(input_fmap_161[7:0]) +
	( 16'sd 25744) * $signed(input_fmap_162[7:0]) +
	( 14'sd 6334) * $signed(input_fmap_163[7:0]) +
	( 11'sd 549) * $signed(input_fmap_164[7:0]) +
	( 13'sd 3819) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19469) * $signed(input_fmap_166[7:0]) +
	( 15'sd 14684) * $signed(input_fmap_167[7:0]) +
	( 16'sd 32089) * $signed(input_fmap_168[7:0]) +
	( 16'sd 17291) * $signed(input_fmap_169[7:0]) +
	( 13'sd 3108) * $signed(input_fmap_170[7:0]) +
	( 15'sd 11120) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6931) * $signed(input_fmap_172[7:0]) +
	( 15'sd 8782) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11201) * $signed(input_fmap_174[7:0]) +
	( 15'sd 13707) * $signed(input_fmap_175[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_176[7:0]) +
	( 16'sd 20474) * $signed(input_fmap_177[7:0]) +
	( 15'sd 12414) * $signed(input_fmap_178[7:0]) +
	( 14'sd 7600) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32650) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28438) * $signed(input_fmap_181[7:0]) +
	( 15'sd 9357) * $signed(input_fmap_182[7:0]) +
	( 16'sd 16994) * $signed(input_fmap_183[7:0]) +
	( 16'sd 20856) * $signed(input_fmap_184[7:0]) +
	( 15'sd 9057) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12259) * $signed(input_fmap_186[7:0]) +
	( 15'sd 14847) * $signed(input_fmap_187[7:0]) +
	( 14'sd 8132) * $signed(input_fmap_188[7:0]) +
	( 16'sd 31822) * $signed(input_fmap_189[7:0]) +
	( 16'sd 23424) * $signed(input_fmap_190[7:0]) +
	( 12'sd 1883) * $signed(input_fmap_191[7:0]) +
	( 16'sd 26488) * $signed(input_fmap_192[7:0]) +
	( 16'sd 19224) * $signed(input_fmap_193[7:0]) +
	( 16'sd 25415) * $signed(input_fmap_194[7:0]) +
	( 16'sd 31397) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24068) * $signed(input_fmap_196[7:0]) +
	( 14'sd 7482) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27750) * $signed(input_fmap_198[7:0]) +
	( 15'sd 9080) * $signed(input_fmap_199[7:0]) +
	( 13'sd 2583) * $signed(input_fmap_200[7:0]) +
	( 16'sd 24079) * $signed(input_fmap_201[7:0]) +
	( 16'sd 25685) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13263) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2625) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2415) * $signed(input_fmap_205[7:0]) +
	( 16'sd 23437) * $signed(input_fmap_206[7:0]) +
	( 16'sd 19459) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18636) * $signed(input_fmap_208[7:0]) +
	( 14'sd 5122) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11314) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10279) * $signed(input_fmap_211[7:0]) +
	( 14'sd 5235) * $signed(input_fmap_212[7:0]) +
	( 14'sd 4543) * $signed(input_fmap_213[7:0]) +
	( 16'sd 27779) * $signed(input_fmap_214[7:0]) +
	( 16'sd 29670) * $signed(input_fmap_215[7:0]) +
	( 16'sd 22638) * $signed(input_fmap_216[7:0]) +
	( 15'sd 8491) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26264) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3537) * $signed(input_fmap_219[7:0]) +
	( 16'sd 28573) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28472) * $signed(input_fmap_221[7:0]) +
	( 16'sd 29091) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14000) * $signed(input_fmap_223[7:0]) +
	( 16'sd 22027) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2272) * $signed(input_fmap_225[7:0]) +
	( 16'sd 18103) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14801) * $signed(input_fmap_227[7:0]) +
	( 15'sd 9157) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20982) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18836) * $signed(input_fmap_230[7:0]) +
	( 15'sd 12391) * $signed(input_fmap_231[7:0]) +
	( 15'sd 13136) * $signed(input_fmap_232[7:0]) +
	( 14'sd 7190) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13121) * $signed(input_fmap_234[7:0]) +
	( 15'sd 13774) * $signed(input_fmap_235[7:0]) +
	( 16'sd 16979) * $signed(input_fmap_236[7:0]) +
	( 16'sd 30981) * $signed(input_fmap_237[7:0]) +
	( 16'sd 23802) * $signed(input_fmap_238[7:0]) +
	( 14'sd 4580) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1526) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_241[7:0]) +
	( 16'sd 20358) * $signed(input_fmap_242[7:0]) +
	( 11'sd 527) * $signed(input_fmap_243[7:0]) +
	( 15'sd 12146) * $signed(input_fmap_244[7:0]) +
	( 11'sd 551) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10726) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3422) * $signed(input_fmap_247[7:0]) +
	( 15'sd 16179) * $signed(input_fmap_248[7:0]) +
	( 16'sd 23770) * $signed(input_fmap_249[7:0]) +
	( 16'sd 23098) * $signed(input_fmap_250[7:0]) +
	( 16'sd 24562) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10819) * $signed(input_fmap_252[7:0]) +
	( 15'sd 10232) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23896) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23637) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_220;
assign conv_mac_220 = 
	( 16'sd 26670) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23016) * $signed(input_fmap_1[7:0]) +
	( 15'sd 11842) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8834) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5727) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14029) * $signed(input_fmap_5[7:0]) +
	( 15'sd 13221) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20375) * $signed(input_fmap_7[7:0]) +
	( 15'sd 14944) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3805) * $signed(input_fmap_9[7:0]) +
	( 16'sd 29116) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23485) * $signed(input_fmap_11[7:0]) +
	( 15'sd 14308) * $signed(input_fmap_12[7:0]) +
	( 16'sd 29276) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22708) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14921) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19656) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30924) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26967) * $signed(input_fmap_18[7:0]) +
	( 15'sd 14526) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22602) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15359) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25469) * $signed(input_fmap_22[7:0]) +
	( 16'sd 16540) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24858) * $signed(input_fmap_24[7:0]) +
	( 16'sd 21346) * $signed(input_fmap_25[7:0]) +
	( 14'sd 5025) * $signed(input_fmap_26[7:0]) +
	( 16'sd 31224) * $signed(input_fmap_27[7:0]) +
	( 16'sd 22513) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1817) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29294) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28189) * $signed(input_fmap_31[7:0]) +
	( 15'sd 13372) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4837) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21326) * $signed(input_fmap_34[7:0]) +
	( 16'sd 16901) * $signed(input_fmap_35[7:0]) +
	( 11'sd 707) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7012) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7973) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29908) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20384) * $signed(input_fmap_40[7:0]) +
	( 14'sd 6292) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14692) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17056) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4753) * $signed(input_fmap_45[7:0]) +
	( 15'sd 13953) * $signed(input_fmap_46[7:0]) +
	( 14'sd 6582) * $signed(input_fmap_47[7:0]) +
	( 15'sd 12837) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30487) * $signed(input_fmap_49[7:0]) +
	( 15'sd 13744) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32729) * $signed(input_fmap_51[7:0]) +
	( 15'sd 14037) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20184) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21819) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11363) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23505) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29830) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2742) * $signed(input_fmap_58[7:0]) +
	( 16'sd 29997) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25614) * $signed(input_fmap_60[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_61[7:0]) +
	( 11'sd 937) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9587) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21754) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_65[7:0]) +
	( 14'sd 4218) * $signed(input_fmap_66[7:0]) +
	( 16'sd 19690) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23762) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1087) * $signed(input_fmap_69[7:0]) +
	( 16'sd 18706) * $signed(input_fmap_70[7:0]) +
	( 15'sd 16357) * $signed(input_fmap_71[7:0]) +
	( 11'sd 717) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4918) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8546) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29902) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30961) * $signed(input_fmap_76[7:0]) +
	( 16'sd 29639) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5776) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_79[7:0]) +
	( 16'sd 29195) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6670) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30010) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1924) * $signed(input_fmap_83[7:0]) +
	( 16'sd 20805) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18760) * $signed(input_fmap_85[7:0]) +
	( 11'sd 615) * $signed(input_fmap_86[7:0]) +
	( 15'sd 13340) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7135) * $signed(input_fmap_88[7:0]) +
	( 16'sd 30886) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29166) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30702) * $signed(input_fmap_91[7:0]) +
	( 14'sd 7648) * $signed(input_fmap_92[7:0]) +
	( 15'sd 14611) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32219) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24420) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10440) * $signed(input_fmap_96[7:0]) +
	( 14'sd 5694) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_98[7:0]) +
	( 15'sd 15858) * $signed(input_fmap_99[7:0]) +
	( 14'sd 6359) * $signed(input_fmap_100[7:0]) +
	( 16'sd 26039) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9622) * $signed(input_fmap_102[7:0]) +
	( 14'sd 6001) * $signed(input_fmap_103[7:0]) +
	( 15'sd 9886) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13076) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9119) * $signed(input_fmap_106[7:0]) +
	( 13'sd 3623) * $signed(input_fmap_107[7:0]) +
	( 16'sd 24714) * $signed(input_fmap_108[7:0]) +
	( 15'sd 8884) * $signed(input_fmap_109[7:0]) +
	( 16'sd 31682) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19117) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13595) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1406) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12514) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27047) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6762) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4300) * $signed(input_fmap_117[7:0]) +
	( 14'sd 5674) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27170) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25172) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4358) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2219) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2865) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27158) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29810) * $signed(input_fmap_126[7:0]) +
	( 16'sd 30071) * $signed(input_fmap_127[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_128[7:0]) +
	( 15'sd 16176) * $signed(input_fmap_129[7:0]) +
	( 16'sd 30969) * $signed(input_fmap_130[7:0]) +
	( 11'sd 993) * $signed(input_fmap_131[7:0]) +
	( 16'sd 27079) * $signed(input_fmap_132[7:0]) +
	( 16'sd 16848) * $signed(input_fmap_133[7:0]) +
	( 16'sd 25664) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18724) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8410) * $signed(input_fmap_136[7:0]) +
	( 13'sd 2069) * $signed(input_fmap_137[7:0]) +
	( 15'sd 8591) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21897) * $signed(input_fmap_139[7:0]) +
	( 16'sd 18336) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22796) * $signed(input_fmap_141[7:0]) +
	( 13'sd 2051) * $signed(input_fmap_142[7:0]) +
	( 13'sd 2598) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31835) * $signed(input_fmap_144[7:0]) +
	( 13'sd 3419) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15455) * $signed(input_fmap_146[7:0]) +
	( 9'sd 217) * $signed(input_fmap_147[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7992) * $signed(input_fmap_149[7:0]) +
	( 16'sd 17606) * $signed(input_fmap_150[7:0]) +
	( 14'sd 8077) * $signed(input_fmap_151[7:0]) +
	( 14'sd 5544) * $signed(input_fmap_152[7:0]) +
	( 14'sd 6512) * $signed(input_fmap_153[7:0]) +
	( 13'sd 3855) * $signed(input_fmap_154[7:0]) +
	( 15'sd 8911) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20315) * $signed(input_fmap_156[7:0]) +
	( 16'sd 31628) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25966) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3368) * $signed(input_fmap_159[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_160[7:0]) +
	( 15'sd 16349) * $signed(input_fmap_161[7:0]) +
	( 16'sd 20861) * $signed(input_fmap_162[7:0]) +
	( 14'sd 5146) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_164[7:0]) +
	( 16'sd 20444) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30644) * $signed(input_fmap_166[7:0]) +
	( 14'sd 6816) * $signed(input_fmap_167[7:0]) +
	( 13'sd 2256) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12455) * $signed(input_fmap_169[7:0]) +
	( 15'sd 16275) * $signed(input_fmap_170[7:0]) +
	( 16'sd 29863) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31134) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1112) * $signed(input_fmap_173[7:0]) +
	( 16'sd 23515) * $signed(input_fmap_174[7:0]) +
	( 16'sd 26533) * $signed(input_fmap_175[7:0]) +
	( 15'sd 14941) * $signed(input_fmap_176[7:0]) +
	( 13'sd 3488) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22621) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28583) * $signed(input_fmap_179[7:0]) +
	( 16'sd 31988) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25958) * $signed(input_fmap_181[7:0]) +
	( 15'sd 14177) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2403) * $signed(input_fmap_183[7:0]) +
	( 16'sd 29379) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11298) * $signed(input_fmap_185[7:0]) +
	( 14'sd 5384) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11526) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32171) * $signed(input_fmap_188[7:0]) +
	( 16'sd 20139) * $signed(input_fmap_189[7:0]) +
	( 15'sd 12875) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24764) * $signed(input_fmap_191[7:0]) +
	( 16'sd 17830) * $signed(input_fmap_192[7:0]) +
	( 15'sd 14224) * $signed(input_fmap_193[7:0]) +
	( 15'sd 10350) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22927) * $signed(input_fmap_195[7:0]) +
	( 16'sd 23961) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21596) * $signed(input_fmap_197[7:0]) +
	( 14'sd 6935) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16153) * $signed(input_fmap_199[7:0]) +
	( 16'sd 21208) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16557) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18733) * $signed(input_fmap_202[7:0]) +
	( 16'sd 26111) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4388) * $signed(input_fmap_204[7:0]) +
	( 14'sd 7335) * $signed(input_fmap_205[7:0]) +
	( 16'sd 25919) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13923) * $signed(input_fmap_207[7:0]) +
	( 15'sd 10329) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18438) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15751) * $signed(input_fmap_210[7:0]) +
	( 16'sd 29155) * $signed(input_fmap_211[7:0]) +
	( 14'sd 7167) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29288) * $signed(input_fmap_213[7:0]) +
	( 16'sd 21403) * $signed(input_fmap_214[7:0]) +
	( 15'sd 13232) * $signed(input_fmap_215[7:0]) +
	( 16'sd 30030) * $signed(input_fmap_216[7:0]) +
	( 16'sd 28066) * $signed(input_fmap_217[7:0]) +
	( 16'sd 23040) * $signed(input_fmap_218[7:0]) +
	( 15'sd 13421) * $signed(input_fmap_219[7:0]) +
	( 14'sd 8014) * $signed(input_fmap_220[7:0]) +
	( 15'sd 14128) * $signed(input_fmap_221[7:0]) +
	( 16'sd 21066) * $signed(input_fmap_222[7:0]) +
	( 15'sd 9318) * $signed(input_fmap_223[7:0]) +
	( 14'sd 4790) * $signed(input_fmap_224[7:0]) +
	( 15'sd 16149) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7622) * $signed(input_fmap_226[7:0]) +
	( 16'sd 18250) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26742) * $signed(input_fmap_228[7:0]) +
	( 16'sd 29095) * $signed(input_fmap_229[7:0]) +
	( 16'sd 23460) * $signed(input_fmap_230[7:0]) +
	( 16'sd 21302) * $signed(input_fmap_231[7:0]) +
	( 11'sd 983) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28605) * $signed(input_fmap_233[7:0]) +
	( 16'sd 16405) * $signed(input_fmap_234[7:0]) +
	( 16'sd 31429) * $signed(input_fmap_235[7:0]) +
	( 16'sd 19986) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11109) * $signed(input_fmap_237[7:0]) +
	( 16'sd 29904) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31026) * $signed(input_fmap_239[7:0]) +
	( 16'sd 24546) * $signed(input_fmap_240[7:0]) +
	( 15'sd 14442) * $signed(input_fmap_241[7:0]) +
	( 16'sd 16492) * $signed(input_fmap_242[7:0]) +
	( 15'sd 9697) * $signed(input_fmap_243[7:0]) +
	( 15'sd 10288) * $signed(input_fmap_244[7:0]) +
	( 15'sd 13320) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_246[7:0]) +
	( 16'sd 22177) * $signed(input_fmap_247[7:0]) +
	( 16'sd 23661) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_249[7:0]) +
	( 14'sd 8038) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19394) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10574) * $signed(input_fmap_252[7:0]) +
	( 16'sd 22095) * $signed(input_fmap_253[7:0]) +
	( 16'sd 17887) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23559) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_221;
assign conv_mac_221 = 
	( 15'sd 12488) * $signed(input_fmap_0[7:0]) +
	( 16'sd 19579) * $signed(input_fmap_1[7:0]) +
	( 16'sd 19498) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30737) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25197) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14698) * $signed(input_fmap_5[7:0]) +
	( 14'sd 6740) * $signed(input_fmap_6[7:0]) +
	( 16'sd 21942) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24492) * $signed(input_fmap_8[7:0]) +
	( 13'sd 3722) * $signed(input_fmap_9[7:0]) +
	( 15'sd 14328) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_11[7:0]) +
	( 14'sd 4406) * $signed(input_fmap_12[7:0]) +
	( 13'sd 2239) * $signed(input_fmap_13[7:0]) +
	( 10'sd 383) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6920) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10561) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2571) * $signed(input_fmap_17[7:0]) +
	( 16'sd 24851) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9784) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17123) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31088) * $signed(input_fmap_21[7:0]) +
	( 14'sd 4529) * $signed(input_fmap_22[7:0]) +
	( 16'sd 28441) * $signed(input_fmap_23[7:0]) +
	( 16'sd 25139) * $signed(input_fmap_24[7:0]) +
	( 9'sd 222) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22699) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13338) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4354) * $signed(input_fmap_28[7:0]) +
	( 15'sd 11279) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4969) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7222) * $signed(input_fmap_31[7:0]) +
	( 16'sd 26138) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13349) * $signed(input_fmap_33[7:0]) +
	( 13'sd 2526) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26485) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1506) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3602) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22533) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5483) * $signed(input_fmap_39[7:0]) +
	( 11'sd 802) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11913) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5920) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8470) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19996) * $signed(input_fmap_44[7:0]) +
	( 13'sd 3285) * $signed(input_fmap_45[7:0]) +
	( 14'sd 6532) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13446) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31758) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25879) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31978) * $signed(input_fmap_51[7:0]) +
	( 14'sd 6734) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6310) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10765) * $signed(input_fmap_55[7:0]) +
	( 16'sd 28665) * $signed(input_fmap_56[7:0]) +
	( 16'sd 31042) * $signed(input_fmap_57[7:0]) +
	( 15'sd 8614) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19060) * $signed(input_fmap_59[7:0]) +
	( 15'sd 15182) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31581) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4780) * $signed(input_fmap_62[7:0]) +
	( 15'sd 12785) * $signed(input_fmap_63[7:0]) +
	( 16'sd 22100) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10110) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9471) * $signed(input_fmap_66[7:0]) +
	( 16'sd 17065) * $signed(input_fmap_67[7:0]) +
	( 16'sd 20431) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26824) * $signed(input_fmap_69[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_70[7:0]) +
	( 16'sd 18326) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4638) * $signed(input_fmap_72[7:0]) +
	( 15'sd 15879) * $signed(input_fmap_73[7:0]) +
	( 15'sd 15685) * $signed(input_fmap_74[7:0]) +
	( 16'sd 31306) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12298) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23319) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7877) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13717) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31507) * $signed(input_fmap_80[7:0]) +
	( 16'sd 31553) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3203) * $signed(input_fmap_83[7:0]) +
	( 16'sd 19607) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1351) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14332) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27925) * $signed(input_fmap_88[7:0]) +
	( 14'sd 8165) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3614) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8204) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22058) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15755) * $signed(input_fmap_93[7:0]) +
	( 15'sd 10740) * $signed(input_fmap_94[7:0]) +
	( 16'sd 18014) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19460) * $signed(input_fmap_96[7:0]) +
	( 16'sd 29676) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30302) * $signed(input_fmap_98[7:0]) +
	( 16'sd 26668) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18480) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6612) * $signed(input_fmap_101[7:0]) +
	( 15'sd 10788) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25959) * $signed(input_fmap_103[7:0]) +
	( 15'sd 10136) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1979) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22695) * $signed(input_fmap_106[7:0]) +
	( 16'sd 27871) * $signed(input_fmap_107[7:0]) +
	( 16'sd 18375) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11612) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22717) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13425) * $signed(input_fmap_111[7:0]) +
	( 16'sd 19656) * $signed(input_fmap_112[7:0]) +
	( 12'sd 1715) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9745) * $signed(input_fmap_114[7:0]) +
	( 15'sd 14763) * $signed(input_fmap_115[7:0]) +
	( 16'sd 17757) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13047) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25203) * $signed(input_fmap_118[7:0]) +
	( 16'sd 25246) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11566) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17768) * $signed(input_fmap_121[7:0]) +
	( 15'sd 16004) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6864) * $signed(input_fmap_123[7:0]) +
	( 15'sd 15531) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20273) * $signed(input_fmap_125[7:0]) +
	( 14'sd 5701) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3063) * $signed(input_fmap_127[7:0]) +
	( 12'sd 1276) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1099) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14116) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19540) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14434) * $signed(input_fmap_132[7:0]) +
	( 13'sd 3714) * $signed(input_fmap_133[7:0]) +
	( 16'sd 17668) * $signed(input_fmap_134[7:0]) +
	( 13'sd 2626) * $signed(input_fmap_135[7:0]) +
	( 16'sd 16627) * $signed(input_fmap_136[7:0]) +
	( 12'sd 1555) * $signed(input_fmap_137[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_138[7:0]) +
	( 8'sd 121) * $signed(input_fmap_139[7:0]) +
	( 16'sd 16955) * $signed(input_fmap_140[7:0]) +
	( 16'sd 17888) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30966) * $signed(input_fmap_142[7:0]) +
	( 15'sd 11923) * $signed(input_fmap_143[7:0]) +
	( 15'sd 12354) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23928) * $signed(input_fmap_145[7:0]) +
	( 16'sd 17202) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13589) * $signed(input_fmap_147[7:0]) +
	( 15'sd 9085) * $signed(input_fmap_148[7:0]) +
	( 14'sd 7413) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31214) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24535) * $signed(input_fmap_151[7:0]) +
	( 15'sd 13751) * $signed(input_fmap_152[7:0]) +
	( 15'sd 13510) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11149) * $signed(input_fmap_154[7:0]) +
	( 15'sd 9302) * $signed(input_fmap_155[7:0]) +
	( 16'sd 21508) * $signed(input_fmap_156[7:0]) +
	( 12'sd 1952) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20799) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2823) * $signed(input_fmap_159[7:0]) +
	( 15'sd 13754) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22066) * $signed(input_fmap_161[7:0]) +
	( 16'sd 32719) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20716) * $signed(input_fmap_163[7:0]) +
	( 15'sd 14608) * $signed(input_fmap_164[7:0]) +
	( 16'sd 25381) * $signed(input_fmap_165[7:0]) +
	( 16'sd 28707) * $signed(input_fmap_166[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1243) * $signed(input_fmap_168[7:0]) +
	( 16'sd 29360) * $signed(input_fmap_169[7:0]) +
	( 12'sd 1270) * $signed(input_fmap_170[7:0]) +
	( 16'sd 30280) * $signed(input_fmap_171[7:0]) +
	( 16'sd 24458) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5718) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16646) * $signed(input_fmap_174[7:0]) +
	( 16'sd 31942) * $signed(input_fmap_175[7:0]) +
	( 16'sd 17281) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6006) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22456) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3736) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28284) * $signed(input_fmap_180[7:0]) +
	( 14'sd 4796) * $signed(input_fmap_181[7:0]) +
	( 15'sd 15869) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17177) * $signed(input_fmap_183[7:0]) +
	( 14'sd 5944) * $signed(input_fmap_184[7:0]) +
	( 16'sd 16844) * $signed(input_fmap_185[7:0]) +
	( 15'sd 14352) * $signed(input_fmap_186[7:0]) +
	( 15'sd 12442) * $signed(input_fmap_187[7:0]) +
	( 16'sd 26179) * $signed(input_fmap_188[7:0]) +
	( 16'sd 20868) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27663) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5582) * $signed(input_fmap_191[7:0]) +
	( 14'sd 7933) * $signed(input_fmap_192[7:0]) +
	( 16'sd 24994) * $signed(input_fmap_193[7:0]) +
	( 15'sd 11414) * $signed(input_fmap_194[7:0]) +
	( 16'sd 16825) * $signed(input_fmap_195[7:0]) +
	( 16'sd 24106) * $signed(input_fmap_196[7:0]) +
	( 16'sd 23945) * $signed(input_fmap_197[7:0]) +
	( 16'sd 22516) * $signed(input_fmap_198[7:0]) +
	( 15'sd 16296) * $signed(input_fmap_199[7:0]) +
	( 16'sd 24414) * $signed(input_fmap_200[7:0]) +
	( 16'sd 27236) * $signed(input_fmap_201[7:0]) +
	( 15'sd 8458) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19020) * $signed(input_fmap_203[7:0]) +
	( 11'sd 528) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30337) * $signed(input_fmap_205[7:0]) +
	( 15'sd 8292) * $signed(input_fmap_206[7:0]) +
	( 16'sd 32701) * $signed(input_fmap_207[7:0]) +
	( 12'sd 1702) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13064) * $signed(input_fmap_209[7:0]) +
	( 16'sd 25032) * $signed(input_fmap_210[7:0]) +
	( 16'sd 25620) * $signed(input_fmap_211[7:0]) +
	( 15'sd 10325) * $signed(input_fmap_212[7:0]) +
	( 16'sd 22588) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23798) * $signed(input_fmap_214[7:0]) +
	( 16'sd 26437) * $signed(input_fmap_215[7:0]) +
	( 16'sd 20054) * $signed(input_fmap_216[7:0]) +
	( 14'sd 4298) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30264) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12965) * $signed(input_fmap_219[7:0]) +
	( 16'sd 25451) * $signed(input_fmap_220[7:0]) +
	( 14'sd 7381) * $signed(input_fmap_221[7:0]) +
	( 16'sd 22933) * $signed(input_fmap_222[7:0]) +
	( 16'sd 18007) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17849) * $signed(input_fmap_224[7:0]) +
	( 15'sd 14256) * $signed(input_fmap_225[7:0]) +
	( 15'sd 9442) * $signed(input_fmap_226[7:0]) +
	( 14'sd 6453) * $signed(input_fmap_227[7:0]) +
	( 16'sd 17643) * $signed(input_fmap_228[7:0]) +
	( 14'sd 7607) * $signed(input_fmap_229[7:0]) +
	( 11'sd 669) * $signed(input_fmap_230[7:0]) +
	( 15'sd 8826) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29639) * $signed(input_fmap_232[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_233[7:0]) +
	( 16'sd 25388) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7780) * $signed(input_fmap_235[7:0]) +
	( 14'sd 6119) * $signed(input_fmap_236[7:0]) +
	( 16'sd 27547) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27747) * $signed(input_fmap_238[7:0]) +
	( 15'sd 10777) * $signed(input_fmap_239[7:0]) +
	( 15'sd 10534) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26333) * $signed(input_fmap_241[7:0]) +
	( 14'sd 6896) * $signed(input_fmap_242[7:0]) +
	( 12'sd 1513) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24718) * $signed(input_fmap_244[7:0]) +
	( 16'sd 16703) * $signed(input_fmap_245[7:0]) +
	( 13'sd 3192) * $signed(input_fmap_246[7:0]) +
	( 14'sd 4253) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26515) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17170) * $signed(input_fmap_249[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_250[7:0]) +
	( 16'sd 32310) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27724) * $signed(input_fmap_252[7:0]) +
	( 15'sd 15650) * $signed(input_fmap_253[7:0]) +
	( 15'sd 15175) * $signed(input_fmap_254[7:0]) +
	( 15'sd 15889) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_222;
assign conv_mac_222 = 
	( 13'sd 3218) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14501) * $signed(input_fmap_1[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15994) * $signed(input_fmap_3[7:0]) +
	( 16'sd 26695) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11615) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30166) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18122) * $signed(input_fmap_7[7:0]) +
	( 16'sd 19489) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1917) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20007) * $signed(input_fmap_10[7:0]) +
	( 16'sd 29739) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3125) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_13[7:0]) +
	( 15'sd 8436) * $signed(input_fmap_14[7:0]) +
	( 16'sd 31930) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28858) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11904) * $signed(input_fmap_17[7:0]) +
	( 16'sd 27109) * $signed(input_fmap_18[7:0]) +
	( 16'sd 32651) * $signed(input_fmap_19[7:0]) +
	( 16'sd 19474) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21975) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16080) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4792) * $signed(input_fmap_23[7:0]) +
	( 15'sd 11360) * $signed(input_fmap_24[7:0]) +
	( 13'sd 2295) * $signed(input_fmap_25[7:0]) +
	( 14'sd 7473) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21276) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17807) * $signed(input_fmap_28[7:0]) +
	( 16'sd 31636) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3525) * $signed(input_fmap_30[7:0]) +
	( 15'sd 13297) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2378) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18558) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5238) * $signed(input_fmap_34[7:0]) +
	( 11'sd 559) * $signed(input_fmap_35[7:0]) +
	( 16'sd 25691) * $signed(input_fmap_36[7:0]) +
	( 16'sd 18747) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2271) * $signed(input_fmap_38[7:0]) +
	( 11'sd 758) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13527) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30397) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25273) * $signed(input_fmap_43[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1365) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5327) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8859) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30138) * $signed(input_fmap_49[7:0]) +
	( 16'sd 22467) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17867) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26756) * $signed(input_fmap_52[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25503) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17895) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_57[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16687) * $signed(input_fmap_59[7:0]) +
	( 15'sd 13669) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11296) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1494) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1532) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17625) * $signed(input_fmap_64[7:0]) +
	( 15'sd 8857) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11675) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16934) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9973) * $signed(input_fmap_68[7:0]) +
	( 16'sd 16510) * $signed(input_fmap_69[7:0]) +
	( 13'sd 2398) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2430) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4569) * $signed(input_fmap_72[7:0]) +
	( 15'sd 9414) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13573) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13692) * $signed(input_fmap_75[7:0]) +
	( 11'sd 690) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18931) * $signed(input_fmap_77[7:0]) +
	( 16'sd 19807) * $signed(input_fmap_78[7:0]) +
	( 14'sd 5000) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5621) * $signed(input_fmap_80[7:0]) +
	( 16'sd 20592) * $signed(input_fmap_81[7:0]) +
	( 15'sd 14940) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30490) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3660) * $signed(input_fmap_84[7:0]) +
	( 16'sd 32584) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14704) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1830) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22473) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23479) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26497) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27882) * $signed(input_fmap_91[7:0]) +
	( 16'sd 30032) * $signed(input_fmap_92[7:0]) +
	( 15'sd 10678) * $signed(input_fmap_93[7:0]) +
	( 15'sd 11572) * $signed(input_fmap_94[7:0]) +
	( 15'sd 16193) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10525) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19237) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22503) * $signed(input_fmap_98[7:0]) +
	( 9'sd 178) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11011) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15354) * $signed(input_fmap_101[7:0]) +
	( 15'sd 11785) * $signed(input_fmap_102[7:0]) +
	( 16'sd 25653) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17091) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26108) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15595) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4152) * $signed(input_fmap_107[7:0]) +
	( 13'sd 3714) * $signed(input_fmap_108[7:0]) +
	( 15'sd 14029) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9256) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32378) * $signed(input_fmap_111[7:0]) +
	( 16'sd 31293) * $signed(input_fmap_112[7:0]) +
	( 10'sd 492) * $signed(input_fmap_113[7:0]) +
	( 16'sd 22452) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25504) * $signed(input_fmap_115[7:0]) +
	( 16'sd 32304) * $signed(input_fmap_116[7:0]) +
	( 16'sd 18926) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7028) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6137) * $signed(input_fmap_121[7:0]) +
	( 11'sd 860) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25963) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17058) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22746) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4959) * $signed(input_fmap_126[7:0]) +
	( 11'sd 987) * $signed(input_fmap_127[7:0]) +
	( 13'sd 2090) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13452) * $signed(input_fmap_129[7:0]) +
	( 9'sd 157) * $signed(input_fmap_130[7:0]) +
	( 12'sd 1276) * $signed(input_fmap_131[7:0]) +
	( 15'sd 16297) * $signed(input_fmap_132[7:0]) +
	( 16'sd 26022) * $signed(input_fmap_133[7:0]) +
	( 16'sd 28315) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23385) * $signed(input_fmap_135[7:0]) +
	( 15'sd 14837) * $signed(input_fmap_136[7:0]) +
	( 9'sd 215) * $signed(input_fmap_137[7:0]) +
	( 14'sd 6639) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27622) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1319) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24579) * $signed(input_fmap_141[7:0]) +
	( 16'sd 32685) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7245) * $signed(input_fmap_143[7:0]) +
	( 16'sd 24943) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28743) * $signed(input_fmap_145[7:0]) +
	( 15'sd 11054) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14767) * $signed(input_fmap_147[7:0]) +
	( 16'sd 24671) * $signed(input_fmap_148[7:0]) +
	( 16'sd 29536) * $signed(input_fmap_149[7:0]) +
	( 15'sd 14442) * $signed(input_fmap_150[7:0]) +
	( 13'sd 3241) * $signed(input_fmap_151[7:0]) +
	( 16'sd 16397) * $signed(input_fmap_152[7:0]) +
	( 15'sd 9084) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6269) * $signed(input_fmap_154[7:0]) +
	( 16'sd 29875) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10009) * $signed(input_fmap_156[7:0]) +
	( 14'sd 4477) * $signed(input_fmap_157[7:0]) +
	( 16'sd 32321) * $signed(input_fmap_158[7:0]) +
	( 16'sd 25981) * $signed(input_fmap_159[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_160[7:0]) +
	( 15'sd 13859) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14386) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3576) * $signed(input_fmap_163[7:0]) +
	( 16'sd 30319) * $signed(input_fmap_164[7:0]) +
	( 12'sd 1400) * $signed(input_fmap_165[7:0]) +
	( 16'sd 24972) * $signed(input_fmap_166[7:0]) +
	( 16'sd 31548) * $signed(input_fmap_167[7:0]) +
	( 16'sd 21663) * $signed(input_fmap_168[7:0]) +
	( 15'sd 12641) * $signed(input_fmap_169[7:0]) +
	( 16'sd 22910) * $signed(input_fmap_170[7:0]) +
	( 14'sd 5358) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_172[7:0]) +
	( 16'sd 32101) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16795) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1941) * $signed(input_fmap_175[7:0]) +
	( 9'sd 153) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15883) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31999) * $signed(input_fmap_178[7:0]) +
	( 15'sd 10450) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15593) * $signed(input_fmap_180[7:0]) +
	( 16'sd 31177) * $signed(input_fmap_181[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_183[7:0]) +
	( 15'sd 9915) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25989) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_186[7:0]) +
	( 14'sd 7875) * $signed(input_fmap_187[7:0]) +
	( 16'sd 28353) * $signed(input_fmap_188[7:0]) +
	( 15'sd 11013) * $signed(input_fmap_189[7:0]) +
	( 16'sd 16849) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17434) * $signed(input_fmap_191[7:0]) +
	( 16'sd 18697) * $signed(input_fmap_192[7:0]) +
	( 16'sd 24677) * $signed(input_fmap_193[7:0]) +
	( 16'sd 16706) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27629) * $signed(input_fmap_195[7:0]) +
	( 16'sd 30631) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21091) * $signed(input_fmap_197[7:0]) +
	( 13'sd 3197) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24980) * $signed(input_fmap_199[7:0]) +
	( 16'sd 30088) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3410) * $signed(input_fmap_201[7:0]) +
	( 15'sd 15744) * $signed(input_fmap_202[7:0]) +
	( 12'sd 1976) * $signed(input_fmap_203[7:0]) +
	( 15'sd 12978) * $signed(input_fmap_204[7:0]) +
	( 16'sd 27955) * $signed(input_fmap_205[7:0]) +
	( 15'sd 15294) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30911) * $signed(input_fmap_207[7:0]) +
	( 15'sd 8498) * $signed(input_fmap_208[7:0]) +
	( 13'sd 2098) * $signed(input_fmap_209[7:0]) +
	( 14'sd 6710) * $signed(input_fmap_210[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_211[7:0]) +
	( 14'sd 7343) * $signed(input_fmap_212[7:0]) +
	( 12'sd 2039) * $signed(input_fmap_213[7:0]) +
	( 16'sd 18991) * $signed(input_fmap_214[7:0]) +
	( 16'sd 20504) * $signed(input_fmap_215[7:0]) +
	( 15'sd 15463) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9655) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31050) * $signed(input_fmap_218[7:0]) +
	( 16'sd 22996) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1373) * $signed(input_fmap_220[7:0]) +
	( 10'sd 376) * $signed(input_fmap_221[7:0]) +
	( 16'sd 25551) * $signed(input_fmap_222[7:0]) +
	( 16'sd 20801) * $signed(input_fmap_223[7:0]) +
	( 16'sd 32153) * $signed(input_fmap_224[7:0]) +
	( 16'sd 24756) * $signed(input_fmap_225[7:0]) +
	( 16'sd 23348) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20075) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24686) * $signed(input_fmap_228[7:0]) +
	( 15'sd 14741) * $signed(input_fmap_229[7:0]) +
	( 14'sd 6950) * $signed(input_fmap_230[7:0]) +
	( 11'sd 516) * $signed(input_fmap_231[7:0]) +
	( 15'sd 10490) * $signed(input_fmap_232[7:0]) +
	( 16'sd 20065) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18714) * $signed(input_fmap_234[7:0]) +
	( 16'sd 22623) * $signed(input_fmap_235[7:0]) +
	( 16'sd 24424) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2049) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31987) * $signed(input_fmap_239[7:0]) +
	( 15'sd 14489) * $signed(input_fmap_240[7:0]) +
	( 16'sd 20022) * $signed(input_fmap_241[7:0]) +
	( 13'sd 3376) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22592) * $signed(input_fmap_243[7:0]) +
	( 15'sd 15018) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14032) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20672) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15025) * $signed(input_fmap_247[7:0]) +
	( 16'sd 25463) * $signed(input_fmap_248[7:0]) +
	( 15'sd 15388) * $signed(input_fmap_249[7:0]) +
	( 16'sd 17489) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27056) * $signed(input_fmap_251[7:0]) +
	( 16'sd 29575) * $signed(input_fmap_252[7:0]) +
	( 15'sd 9036) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20780) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_223;
assign conv_mac_223 = 
	( 16'sd 20764) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27595) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31485) * $signed(input_fmap_2[7:0]) +
	( 15'sd 14968) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12023) * $signed(input_fmap_4[7:0]) +
	( 16'sd 22910) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21320) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20608) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17340) * $signed(input_fmap_8[7:0]) +
	( 16'sd 21623) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12414) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2641) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21108) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14438) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15289) * $signed(input_fmap_14[7:0]) +
	( 16'sd 20337) * $signed(input_fmap_15[7:0]) +
	( 16'sd 20466) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19303) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5397) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10395) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9664) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20220) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19232) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10254) * $signed(input_fmap_23[7:0]) +
	( 15'sd 12861) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20223) * $signed(input_fmap_25[7:0]) +
	( 15'sd 11703) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26315) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26509) * $signed(input_fmap_28[7:0]) +
	( 16'sd 28770) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5700) * $signed(input_fmap_31[7:0]) +
	( 16'sd 31680) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28548) * $signed(input_fmap_33[7:0]) +
	( 15'sd 8753) * $signed(input_fmap_34[7:0]) +
	( 16'sd 17956) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10555) * $signed(input_fmap_36[7:0]) +
	( 11'sd 793) * $signed(input_fmap_37[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7493) * $signed(input_fmap_39[7:0]) +
	( 16'sd 31477) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5455) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11684) * $signed(input_fmap_42[7:0]) +
	( 14'sd 5389) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17414) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4596) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14167) * $signed(input_fmap_46[7:0]) +
	( 16'sd 19397) * $signed(input_fmap_47[7:0]) +
	( 16'sd 21091) * $signed(input_fmap_48[7:0]) +
	( 15'sd 9633) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12402) * $signed(input_fmap_50[7:0]) +
	( 15'sd 11574) * $signed(input_fmap_51[7:0]) +
	( 6'sd 20) * $signed(input_fmap_52[7:0]) +
	( 10'sd 382) * $signed(input_fmap_53[7:0]) +
	( 13'sd 4036) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19075) * $signed(input_fmap_56[7:0]) +
	( 10'sd 326) * $signed(input_fmap_57[7:0]) +
	( 13'sd 2558) * $signed(input_fmap_58[7:0]) +
	( 16'sd 16643) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9267) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19808) * $signed(input_fmap_61[7:0]) +
	( 12'sd 1213) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29321) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15767) * $signed(input_fmap_64[7:0]) +
	( 15'sd 12323) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30640) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6914) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13098) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29123) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6027) * $signed(input_fmap_70[7:0]) +
	( 11'sd 996) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25941) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14045) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17399) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23132) * $signed(input_fmap_75[7:0]) +
	( 16'sd 27394) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32373) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10344) * $signed(input_fmap_78[7:0]) +
	( 16'sd 18756) * $signed(input_fmap_79[7:0]) +
	( 15'sd 13622) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23779) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9498) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27661) * $signed(input_fmap_83[7:0]) +
	( 15'sd 13246) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12671) * $signed(input_fmap_85[7:0]) +
	( 16'sd 16456) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5304) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6261) * $signed(input_fmap_88[7:0]) +
	( 16'sd 23674) * $signed(input_fmap_89[7:0]) +
	( 16'sd 31228) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8855) * $signed(input_fmap_91[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_92[7:0]) +
	( 14'sd 8021) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25916) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5062) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25341) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1212) * $signed(input_fmap_97[7:0]) +
	( 16'sd 30784) * $signed(input_fmap_98[7:0]) +
	( 16'sd 19217) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23034) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3273) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27312) * $signed(input_fmap_102[7:0]) +
	( 16'sd 30653) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20835) * $signed(input_fmap_104[7:0]) +
	( 12'sd 1468) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3614) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5298) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30452) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24773) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2757) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15200) * $signed(input_fmap_111[7:0]) +
	( 16'sd 18482) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10243) * $signed(input_fmap_113[7:0]) +
	( 16'sd 29450) * $signed(input_fmap_114[7:0]) +
	( 16'sd 30170) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6347) * $signed(input_fmap_116[7:0]) +
	( 15'sd 14319) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13830) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27181) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10563) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17745) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19623) * $signed(input_fmap_122[7:0]) +
	( 14'sd 4428) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22529) * $signed(input_fmap_124[7:0]) +
	( 16'sd 16909) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29510) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10089) * $signed(input_fmap_127[7:0]) +
	( 16'sd 28688) * $signed(input_fmap_128[7:0]) +
	( 15'sd 9796) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22236) * $signed(input_fmap_130[7:0]) +
	( 15'sd 9353) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8814) * $signed(input_fmap_132[7:0]) +
	( 12'sd 1530) * $signed(input_fmap_133[7:0]) +
	( 14'sd 6293) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1850) * $signed(input_fmap_136[7:0]) +
	( 14'sd 8180) * $signed(input_fmap_137[7:0]) +
	( 16'sd 25351) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2085) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28897) * $signed(input_fmap_140[7:0]) +
	( 16'sd 24352) * $signed(input_fmap_141[7:0]) +
	( 15'sd 13420) * $signed(input_fmap_142[7:0]) +
	( 16'sd 27695) * $signed(input_fmap_143[7:0]) +
	( 12'sd 1429) * $signed(input_fmap_144[7:0]) +
	( 15'sd 16026) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7298) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30320) * $signed(input_fmap_147[7:0]) +
	( 16'sd 29225) * $signed(input_fmap_148[7:0]) +
	( 16'sd 27159) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27197) * $signed(input_fmap_150[7:0]) +
	( 15'sd 15096) * $signed(input_fmap_151[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10295) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25981) * $signed(input_fmap_154[7:0]) +
	( 16'sd 28434) * $signed(input_fmap_155[7:0]) +
	( 16'sd 23463) * $signed(input_fmap_156[7:0]) +
	( 16'sd 22055) * $signed(input_fmap_157[7:0]) +
	( 12'sd 1878) * $signed(input_fmap_158[7:0]) +
	( 16'sd 24193) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6188) * $signed(input_fmap_160[7:0]) +
	( 15'sd 11069) * $signed(input_fmap_161[7:0]) +
	( 16'sd 19496) * $signed(input_fmap_162[7:0]) +
	( 11'sd 888) * $signed(input_fmap_163[7:0]) +
	( 15'sd 15731) * $signed(input_fmap_164[7:0]) +
	( 13'sd 4058) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31385) * $signed(input_fmap_166[7:0]) +
	( 14'sd 6097) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9282) * $signed(input_fmap_168[7:0]) +
	( 15'sd 9674) * $signed(input_fmap_169[7:0]) +
	( 16'sd 23991) * $signed(input_fmap_170[7:0]) +
	( 16'sd 25443) * $signed(input_fmap_171[7:0]) +
	( 16'sd 21349) * $signed(input_fmap_172[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_173[7:0]) +
	( 15'sd 13846) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17608) * $signed(input_fmap_175[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_176[7:0]) +
	( 14'sd 8020) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27143) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25656) * $signed(input_fmap_179[7:0]) +
	( 16'sd 18833) * $signed(input_fmap_180[7:0]) +
	( 16'sd 20007) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10089) * $signed(input_fmap_182[7:0]) +
	( 15'sd 11123) * $signed(input_fmap_183[7:0]) +
	( 15'sd 10813) * $signed(input_fmap_184[7:0]) +
	( 16'sd 22219) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18673) * $signed(input_fmap_186[7:0]) +
	( 15'sd 16285) * $signed(input_fmap_187[7:0]) +
	( 14'sd 5518) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3276) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30776) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19176) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20565) * $signed(input_fmap_192[7:0]) +
	( 16'sd 28647) * $signed(input_fmap_193[7:0]) +
	( 16'sd 32674) * $signed(input_fmap_194[7:0]) +
	( 16'sd 32724) * $signed(input_fmap_195[7:0]) +
	( 15'sd 16009) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21297) * $signed(input_fmap_197[7:0]) +
	( 16'sd 32640) * $signed(input_fmap_198[7:0]) +
	( 16'sd 26544) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18150) * $signed(input_fmap_200[7:0]) +
	( 14'sd 7417) * $signed(input_fmap_201[7:0]) +
	( 14'sd 6748) * $signed(input_fmap_202[7:0]) +
	( 11'sd 707) * $signed(input_fmap_203[7:0]) +
	( 16'sd 27127) * $signed(input_fmap_204[7:0]) +
	( 12'sd 1395) * $signed(input_fmap_205[7:0]) +
	( 15'sd 8769) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1551) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15716) * $signed(input_fmap_208[7:0]) +
	( 14'sd 7423) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15214) * $signed(input_fmap_210[7:0]) +
	( 16'sd 16416) * $signed(input_fmap_211[7:0]) +
	( 14'sd 7790) * $signed(input_fmap_212[7:0]) +
	( 9'sd 184) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28653) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10367) * $signed(input_fmap_215[7:0]) +
	( 16'sd 30966) * $signed(input_fmap_216[7:0]) +
	( 16'sd 21887) * $signed(input_fmap_217[7:0]) +
	( 15'sd 11658) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21514) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24238) * $signed(input_fmap_220[7:0]) +
	( 16'sd 26544) * $signed(input_fmap_221[7:0]) +
	( 16'sd 21790) * $signed(input_fmap_222[7:0]) +
	( 15'sd 11970) * $signed(input_fmap_223[7:0]) +
	( 15'sd 13178) * $signed(input_fmap_224[7:0]) +
	( 16'sd 19599) * $signed(input_fmap_225[7:0]) +
	( 14'sd 5654) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5441) * $signed(input_fmap_227[7:0]) +
	( 14'sd 7673) * $signed(input_fmap_228[7:0]) +
	( 14'sd 5387) * $signed(input_fmap_229[7:0]) +
	( 11'sd 1018) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7815) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8193) * $signed(input_fmap_232[7:0]) +
	( 16'sd 32179) * $signed(input_fmap_233[7:0]) +
	( 16'sd 32630) * $signed(input_fmap_234[7:0]) +
	( 16'sd 25793) * $signed(input_fmap_235[7:0]) +
	( 15'sd 16365) * $signed(input_fmap_236[7:0]) +
	( 16'sd 31569) * $signed(input_fmap_237[7:0]) +
	( 15'sd 15344) * $signed(input_fmap_238[7:0]) +
	( 15'sd 10963) * $signed(input_fmap_239[7:0]) +
	( 16'sd 21591) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21444) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11207) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7026) * $signed(input_fmap_243[7:0]) +
	( 15'sd 9233) * $signed(input_fmap_244[7:0]) +
	( 6'sd 20) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19720) * $signed(input_fmap_246[7:0]) +
	( 12'sd 2029) * $signed(input_fmap_247[7:0]) +
	( 14'sd 7679) * $signed(input_fmap_248[7:0]) +
	( 13'sd 3060) * $signed(input_fmap_249[7:0]) +
	( 12'sd 1948) * $signed(input_fmap_250[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_251[7:0]) +
	( 7'sd 45) * $signed(input_fmap_252[7:0]) +
	( 14'sd 7816) * $signed(input_fmap_253[7:0]) +
	( 15'sd 16272) * $signed(input_fmap_254[7:0]) +
	( 16'sd 31182) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_224;
assign conv_mac_224 = 
	( 10'sd 468) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7200) * $signed(input_fmap_1[7:0]) +
	( 16'sd 23176) * $signed(input_fmap_2[7:0]) +
	( 15'sd 10365) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5557) * $signed(input_fmap_4[7:0]) +
	( 13'sd 3366) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17042) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1345) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30579) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29048) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21122) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10230) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7921) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31514) * $signed(input_fmap_13[7:0]) +
	( 16'sd 24515) * $signed(input_fmap_14[7:0]) +
	( 14'sd 6064) * $signed(input_fmap_15[7:0]) +
	( 16'sd 19360) * $signed(input_fmap_16[7:0]) +
	( 16'sd 28828) * $signed(input_fmap_17[7:0]) +
	( 15'sd 9875) * $signed(input_fmap_18[7:0]) +
	( 11'sd 605) * $signed(input_fmap_19[7:0]) +
	( 16'sd 32313) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12203) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7058) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_23[7:0]) +
	( 14'sd 5492) * $signed(input_fmap_24[7:0]) +
	( 10'sd 404) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4545) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22468) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2079) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14335) * $signed(input_fmap_29[7:0]) +
	( 13'sd 3606) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15975) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17181) * $signed(input_fmap_32[7:0]) +
	( 16'sd 22047) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24491) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19870) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7212) * $signed(input_fmap_36[7:0]) +
	( 15'sd 15936) * $signed(input_fmap_37[7:0]) +
	( 16'sd 31868) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25031) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23716) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26799) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31690) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24789) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3561) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9736) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23851) * $signed(input_fmap_46[7:0]) +
	( 16'sd 27307) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24445) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17945) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26820) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12314) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5079) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13223) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13555) * $signed(input_fmap_54[7:0]) +
	( 16'sd 20931) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31924) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28667) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15413) * $signed(input_fmap_58[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26486) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19214) * $signed(input_fmap_61[7:0]) +
	( 14'sd 7598) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1564) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18832) * $signed(input_fmap_64[7:0]) +
	( 16'sd 22582) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25634) * $signed(input_fmap_66[7:0]) +
	( 15'sd 11366) * $signed(input_fmap_67[7:0]) +
	( 15'sd 12556) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8562) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10397) * $signed(input_fmap_70[7:0]) +
	( 13'sd 3750) * $signed(input_fmap_71[7:0]) +
	( 15'sd 11224) * $signed(input_fmap_72[7:0]) +
	( 16'sd 25926) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17858) * $signed(input_fmap_74[7:0]) +
	( 16'sd 18723) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9557) * $signed(input_fmap_76[7:0]) +
	( 16'sd 26785) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12262) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11872) * $signed(input_fmap_79[7:0]) +
	( 15'sd 9980) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25016) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27491) * $signed(input_fmap_82[7:0]) +
	( 14'sd 7356) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11482) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18508) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23549) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18378) * $signed(input_fmap_87[7:0]) +
	( 15'sd 13293) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25750) * $signed(input_fmap_89[7:0]) +
	( 13'sd 3142) * $signed(input_fmap_90[7:0]) +
	( 14'sd 4277) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27754) * $signed(input_fmap_92[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16531) * $signed(input_fmap_94[7:0]) +
	( 16'sd 16855) * $signed(input_fmap_95[7:0]) +
	( 15'sd 12036) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14035) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17048) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5183) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23190) * $signed(input_fmap_100[7:0]) +
	( 12'sd 1757) * $signed(input_fmap_101[7:0]) +
	( 14'sd 5693) * $signed(input_fmap_102[7:0]) +
	( 16'sd 23506) * $signed(input_fmap_103[7:0]) +
	( 15'sd 14944) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9886) * $signed(input_fmap_105[7:0]) +
	( 13'sd 3541) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17805) * $signed(input_fmap_108[7:0]) +
	( 12'sd 1312) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19817) * $signed(input_fmap_110[7:0]) +
	( 13'sd 3795) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22061) * $signed(input_fmap_112[7:0]) +
	( 16'sd 22809) * $signed(input_fmap_113[7:0]) +
	( 16'sd 24312) * $signed(input_fmap_114[7:0]) +
	( 15'sd 9044) * $signed(input_fmap_115[7:0]) +
	( 13'sd 2120) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6345) * $signed(input_fmap_117[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16532) * $signed(input_fmap_119[7:0]) +
	( 16'sd 26979) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30497) * $signed(input_fmap_121[7:0]) +
	( 16'sd 18273) * $signed(input_fmap_122[7:0]) +
	( 13'sd 2797) * $signed(input_fmap_123[7:0]) +
	( 15'sd 14058) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9878) * $signed(input_fmap_125[7:0]) +
	( 16'sd 25756) * $signed(input_fmap_126[7:0]) +
	( 16'sd 27073) * $signed(input_fmap_127[7:0]) +
	( 16'sd 32566) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5889) * $signed(input_fmap_129[7:0]) +
	( 14'sd 7557) * $signed(input_fmap_130[7:0]) +
	( 16'sd 26316) * $signed(input_fmap_131[7:0]) +
	( 11'sd 975) * $signed(input_fmap_132[7:0]) +
	( 15'sd 9822) * $signed(input_fmap_133[7:0]) +
	( 16'sd 16696) * $signed(input_fmap_134[7:0]) +
	( 15'sd 16223) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30182) * $signed(input_fmap_136[7:0]) +
	( 16'sd 25173) * $signed(input_fmap_137[7:0]) +
	( 16'sd 25004) * $signed(input_fmap_138[7:0]) +
	( 16'sd 27928) * $signed(input_fmap_139[7:0]) +
	( 16'sd 16717) * $signed(input_fmap_140[7:0]) +
	( 15'sd 16358) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25452) * $signed(input_fmap_142[7:0]) +
	( 16'sd 29819) * $signed(input_fmap_143[7:0]) +
	( 16'sd 22948) * $signed(input_fmap_144[7:0]) +
	( 12'sd 1795) * $signed(input_fmap_145[7:0]) +
	( 14'sd 7255) * $signed(input_fmap_146[7:0]) +
	( 14'sd 5753) * $signed(input_fmap_147[7:0]) +
	( 16'sd 27268) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12718) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21196) * $signed(input_fmap_150[7:0]) +
	( 16'sd 22687) * $signed(input_fmap_151[7:0]) +
	( 16'sd 25467) * $signed(input_fmap_152[7:0]) +
	( 16'sd 18172) * $signed(input_fmap_153[7:0]) +
	( 15'sd 13854) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19321) * $signed(input_fmap_155[7:0]) +
	( 13'sd 2242) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15065) * $signed(input_fmap_157[7:0]) +
	( 16'sd 24486) * $signed(input_fmap_158[7:0]) +
	( 15'sd 16090) * $signed(input_fmap_159[7:0]) +
	( 10'sd 472) * $signed(input_fmap_160[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21364) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8790) * $signed(input_fmap_163[7:0]) +
	( 16'sd 32419) * $signed(input_fmap_164[7:0]) +
	( 7'sd 45) * $signed(input_fmap_165[7:0]) +
	( 15'sd 14312) * $signed(input_fmap_166[7:0]) +
	( 16'sd 19699) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20692) * $signed(input_fmap_168[7:0]) +
	( 16'sd 19326) * $signed(input_fmap_169[7:0]) +
	( 16'sd 26332) * $signed(input_fmap_170[7:0]) +
	( 16'sd 23427) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12230) * $signed(input_fmap_172[7:0]) +
	( 15'sd 16300) * $signed(input_fmap_173[7:0]) +
	( 15'sd 16128) * $signed(input_fmap_174[7:0]) +
	( 15'sd 8995) * $signed(input_fmap_175[7:0]) +
	( 9'sd 130) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27856) * $signed(input_fmap_177[7:0]) +
	( 11'sd 625) * $signed(input_fmap_178[7:0]) +
	( 15'sd 12232) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24665) * $signed(input_fmap_180[7:0]) +
	( 14'sd 8016) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10618) * $signed(input_fmap_182[7:0]) +
	( 14'sd 4299) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8359) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15145) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26600) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25583) * $signed(input_fmap_187[7:0]) +
	( 16'sd 18732) * $signed(input_fmap_188[7:0]) +
	( 15'sd 8605) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5139) * $signed(input_fmap_190[7:0]) +
	( 16'sd 30425) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15867) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_193[7:0]) +
	( 16'sd 32721) * $signed(input_fmap_194[7:0]) +
	( 15'sd 13197) * $signed(input_fmap_195[7:0]) +
	( 15'sd 13017) * $signed(input_fmap_196[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24065) * $signed(input_fmap_198[7:0]) +
	( 16'sd 17513) * $signed(input_fmap_199[7:0]) +
	( 16'sd 20061) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3558) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2478) * $signed(input_fmap_202[7:0]) +
	( 11'sd 917) * $signed(input_fmap_203[7:0]) +
	( 15'sd 8775) * $signed(input_fmap_204[7:0]) +
	( 16'sd 30605) * $signed(input_fmap_205[7:0]) +
	( 16'sd 17615) * $signed(input_fmap_206[7:0]) +
	( 16'sd 31174) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17588) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13427) * $signed(input_fmap_209[7:0]) +
	( 15'sd 9386) * $signed(input_fmap_210[7:0]) +
	( 16'sd 24846) * $signed(input_fmap_211[7:0]) +
	( 16'sd 28230) * $signed(input_fmap_212[7:0]) +
	( 15'sd 10110) * $signed(input_fmap_213[7:0]) +
	( 16'sd 22532) * $signed(input_fmap_214[7:0]) +
	( 15'sd 13390) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19844) * $signed(input_fmap_216[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_217[7:0]) +
	( 15'sd 13712) * $signed(input_fmap_218[7:0]) +
	( 15'sd 14856) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30499) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13834) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18694) * $signed(input_fmap_222[7:0]) +
	( 12'sd 1511) * $signed(input_fmap_223[7:0]) +
	( 14'sd 7898) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5274) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14158) * $signed(input_fmap_226[7:0]) +
	( 16'sd 28592) * $signed(input_fmap_227[7:0]) +
	( 15'sd 13961) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24111) * $signed(input_fmap_229[7:0]) +
	( 11'sd 885) * $signed(input_fmap_230[7:0]) +
	( 15'sd 15194) * $signed(input_fmap_231[7:0]) +
	( 14'sd 6979) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5758) * $signed(input_fmap_233[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_234[7:0]) +
	( 13'sd 2944) * $signed(input_fmap_235[7:0]) +
	( 11'sd 527) * $signed(input_fmap_236[7:0]) +
	( 16'sd 21293) * $signed(input_fmap_237[7:0]) +
	( 16'sd 32199) * $signed(input_fmap_238[7:0]) +
	( 16'sd 28589) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26206) * $signed(input_fmap_240[7:0]) +
	( 15'sd 12517) * $signed(input_fmap_241[7:0]) +
	( 15'sd 8361) * $signed(input_fmap_242[7:0]) +
	( 16'sd 30513) * $signed(input_fmap_243[7:0]) +
	( 16'sd 27957) * $signed(input_fmap_244[7:0]) +
	( 11'sd 550) * $signed(input_fmap_245[7:0]) +
	( 14'sd 5695) * $signed(input_fmap_246[7:0]) +
	( 14'sd 5524) * $signed(input_fmap_247[7:0]) +
	( 16'sd 17635) * $signed(input_fmap_248[7:0]) +
	( 8'sd 99) * $signed(input_fmap_249[7:0]) +
	( 16'sd 23014) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22563) * $signed(input_fmap_251[7:0]) +
	( 15'sd 9964) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5145) * $signed(input_fmap_253[7:0]) +
	( 14'sd 7775) * $signed(input_fmap_254[7:0]) +
	( 16'sd 21506) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_225;
assign conv_mac_225 = 
	( 16'sd 25828) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10485) * $signed(input_fmap_1[7:0]) +
	( 16'sd 26852) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12501) * $signed(input_fmap_3[7:0]) +
	( 16'sd 23179) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21916) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22508) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18350) * $signed(input_fmap_7[7:0]) +
	( 14'sd 5667) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20468) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10606) * $signed(input_fmap_10[7:0]) +
	( 14'sd 5173) * $signed(input_fmap_11[7:0]) +
	( 16'sd 31815) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15493) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1315) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28040) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25668) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14747) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27135) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23091) * $signed(input_fmap_20[7:0]) +
	( 11'sd 656) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27686) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14688) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28216) * $signed(input_fmap_24[7:0]) +
	( 16'sd 26050) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28439) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23721) * $signed(input_fmap_27[7:0]) +
	( 14'sd 6339) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6587) * $signed(input_fmap_29[7:0]) +
	( 15'sd 16004) * $signed(input_fmap_30[7:0]) +
	( 16'sd 24390) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28086) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4821) * $signed(input_fmap_33[7:0]) +
	( 15'sd 14630) * $signed(input_fmap_34[7:0]) +
	( 16'sd 19514) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20893) * $signed(input_fmap_36[7:0]) +
	( 15'sd 10381) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8437) * $signed(input_fmap_38[7:0]) +
	( 16'sd 32357) * $signed(input_fmap_39[7:0]) +
	( 14'sd 8166) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31095) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12232) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25435) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15078) * $signed(input_fmap_44[7:0]) +
	( 16'sd 20169) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10738) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31927) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8632) * $signed(input_fmap_48[7:0]) +
	( 16'sd 17417) * $signed(input_fmap_49[7:0]) +
	( 16'sd 29702) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29694) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22030) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22091) * $signed(input_fmap_53[7:0]) +
	( 15'sd 10278) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8790) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19140) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4921) * $signed(input_fmap_57[7:0]) +
	( 15'sd 9685) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12680) * $signed(input_fmap_59[7:0]) +
	( 15'sd 8367) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27262) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23797) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25286) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19089) * $signed(input_fmap_64[7:0]) +
	( 16'sd 31795) * $signed(input_fmap_65[7:0]) +
	( 16'sd 22156) * $signed(input_fmap_66[7:0]) +
	( 16'sd 27893) * $signed(input_fmap_67[7:0]) +
	( 16'sd 17088) * $signed(input_fmap_68[7:0]) +
	( 16'sd 18578) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3491) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19693) * $signed(input_fmap_71[7:0]) +
	( 14'sd 5516) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7579) * $signed(input_fmap_73[7:0]) +
	( 16'sd 23282) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15767) * $signed(input_fmap_75[7:0]) +
	( 14'sd 4224) * $signed(input_fmap_76[7:0]) +
	( 16'sd 20706) * $signed(input_fmap_77[7:0]) +
	( 14'sd 7102) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20705) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24136) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25524) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3763) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32194) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2999) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5438) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4577) * $signed(input_fmap_86[7:0]) +
	( 14'sd 7901) * $signed(input_fmap_87[7:0]) +
	( 15'sd 16168) * $signed(input_fmap_88[7:0]) +
	( 16'sd 20353) * $signed(input_fmap_89[7:0]) +
	( 16'sd 18095) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31607) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28529) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32270) * $signed(input_fmap_93[7:0]) +
	( 12'sd 1697) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24350) * $signed(input_fmap_95[7:0]) +
	( 14'sd 5668) * $signed(input_fmap_96[7:0]) +
	( 16'sd 30462) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2101) * $signed(input_fmap_98[7:0]) +
	( 4'sd 7) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13723) * $signed(input_fmap_100[7:0]) +
	( 13'sd 3446) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16251) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11024) * $signed(input_fmap_103[7:0]) +
	( 15'sd 11106) * $signed(input_fmap_104[7:0]) +
	( 13'sd 2274) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1952) * $signed(input_fmap_106[7:0]) +
	( 14'sd 8135) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2783) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2953) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29708) * $signed(input_fmap_110[7:0]) +
	( 14'sd 6153) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17059) * $signed(input_fmap_112[7:0]) +
	( 16'sd 25564) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32326) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1929) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7357) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25048) * $signed(input_fmap_117[7:0]) +
	( 16'sd 30619) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19920) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21129) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16527) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25706) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18072) * $signed(input_fmap_123[7:0]) +
	( 16'sd 29558) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26288) * $signed(input_fmap_125[7:0]) +
	( 16'sd 19171) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15024) * $signed(input_fmap_127[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_128[7:0]) +
	( 15'sd 16164) * $signed(input_fmap_129[7:0]) +
	( 9'sd 140) * $signed(input_fmap_130[7:0]) +
	( 7'sd 51) * $signed(input_fmap_131[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10584) * $signed(input_fmap_133[7:0]) +
	( 15'sd 10778) * $signed(input_fmap_134[7:0]) +
	( 15'sd 15444) * $signed(input_fmap_135[7:0]) +
	( 14'sd 6234) * $signed(input_fmap_136[7:0]) +
	( 15'sd 13379) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29804) * $signed(input_fmap_138[7:0]) +
	( 15'sd 13261) * $signed(input_fmap_139[7:0]) +
	( 14'sd 7090) * $signed(input_fmap_140[7:0]) +
	( 14'sd 4943) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21464) * $signed(input_fmap_142[7:0]) +
	( 13'sd 2297) * $signed(input_fmap_143[7:0]) +
	( 16'sd 16822) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8373) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21093) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8969) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26437) * $signed(input_fmap_148[7:0]) +
	( 15'sd 14032) * $signed(input_fmap_149[7:0]) +
	( 15'sd 11052) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24218) * $signed(input_fmap_151[7:0]) +
	( 16'sd 20583) * $signed(input_fmap_152[7:0]) +
	( 16'sd 32272) * $signed(input_fmap_153[7:0]) +
	( 16'sd 22920) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11458) * $signed(input_fmap_157[7:0]) +
	( 16'sd 30801) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6188) * $signed(input_fmap_159[7:0]) +
	( 15'sd 12147) * $signed(input_fmap_160[7:0]) +
	( 16'sd 20884) * $signed(input_fmap_161[7:0]) +
	( 15'sd 14488) * $signed(input_fmap_162[7:0]) +
	( 16'sd 24570) * $signed(input_fmap_163[7:0]) +
	( 16'sd 20485) * $signed(input_fmap_164[7:0]) +
	( 13'sd 3395) * $signed(input_fmap_165[7:0]) +
	( 16'sd 24099) * $signed(input_fmap_166[7:0]) +
	( 16'sd 20675) * $signed(input_fmap_167[7:0]) +
	( 9'sd 191) * $signed(input_fmap_168[7:0]) +
	( 15'sd 13361) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28527) * $signed(input_fmap_170[7:0]) +
	( 14'sd 8038) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1346) * $signed(input_fmap_172[7:0]) +
	( 14'sd 4894) * $signed(input_fmap_173[7:0]) +
	( 13'sd 3129) * $signed(input_fmap_174[7:0]) +
	( 16'sd 27590) * $signed(input_fmap_175[7:0]) +
	( 15'sd 10195) * $signed(input_fmap_176[7:0]) +
	( 15'sd 15284) * $signed(input_fmap_177[7:0]) +
	( 15'sd 8785) * $signed(input_fmap_178[7:0]) +
	( 16'sd 19803) * $signed(input_fmap_179[7:0]) +
	( 16'sd 28282) * $signed(input_fmap_180[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_181[7:0]) +
	( 16'sd 23836) * $signed(input_fmap_182[7:0]) +
	( 16'sd 16613) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26981) * $signed(input_fmap_184[7:0]) +
	( 16'sd 32338) * $signed(input_fmap_185[7:0]) +
	( 14'sd 5173) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25263) * $signed(input_fmap_187[7:0]) +
	( 16'sd 27025) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_189[7:0]) +
	( 15'sd 13733) * $signed(input_fmap_190[7:0]) +
	( 16'sd 26643) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22835) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9067) * $signed(input_fmap_193[7:0]) +
	( 8'sd 105) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1586) * $signed(input_fmap_195[7:0]) +
	( 12'sd 1827) * $signed(input_fmap_196[7:0]) +
	( 13'sd 4065) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27900) * $signed(input_fmap_198[7:0]) +
	( 16'sd 26298) * $signed(input_fmap_199[7:0]) +
	( 14'sd 5928) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18374) * $signed(input_fmap_201[7:0]) +
	( 10'sd 494) * $signed(input_fmap_202[7:0]) +
	( 12'sd 1704) * $signed(input_fmap_203[7:0]) +
	( 15'sd 9844) * $signed(input_fmap_204[7:0]) +
	( 11'sd 702) * $signed(input_fmap_205[7:0]) +
	( 13'sd 2059) * $signed(input_fmap_206[7:0]) +
	( 14'sd 4629) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18508) * $signed(input_fmap_208[7:0]) +
	( 15'sd 10293) * $signed(input_fmap_209[7:0]) +
	( 16'sd 22206) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23141) * $signed(input_fmap_211[7:0]) +
	( 16'sd 27239) * $signed(input_fmap_212[7:0]) +
	( 15'sd 14804) * $signed(input_fmap_213[7:0]) +
	( 15'sd 11943) * $signed(input_fmap_214[7:0]) +
	( 16'sd 23795) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19129) * $signed(input_fmap_216[7:0]) +
	( 16'sd 18000) * $signed(input_fmap_217[7:0]) +
	( 14'sd 6246) * $signed(input_fmap_218[7:0]) +
	( 13'sd 4033) * $signed(input_fmap_219[7:0]) +
	( 16'sd 22535) * $signed(input_fmap_220[7:0]) +
	( 15'sd 13502) * $signed(input_fmap_221[7:0]) +
	( 15'sd 15899) * $signed(input_fmap_222[7:0]) +
	( 14'sd 4757) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25605) * $signed(input_fmap_224[7:0]) +
	( 16'sd 17668) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11104) * $signed(input_fmap_226[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10479) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23959) * $signed(input_fmap_229[7:0]) +
	( 16'sd 27693) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1801) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29370) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5219) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23697) * $signed(input_fmap_234[7:0]) +
	( 13'sd 2772) * $signed(input_fmap_235[7:0]) +
	( 15'sd 8552) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19147) * $signed(input_fmap_237[7:0]) +
	( 16'sd 32040) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31252) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18139) * $signed(input_fmap_240[7:0]) +
	( 15'sd 9545) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29046) * $signed(input_fmap_242[7:0]) +
	( 15'sd 15193) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_244[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19492) * $signed(input_fmap_246[7:0]) +
	( 12'sd 1970) * $signed(input_fmap_247[7:0]) +
	( 16'sd 24626) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4236) * $signed(input_fmap_249[7:0]) +
	( 13'sd 3754) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4940) * $signed(input_fmap_251[7:0]) +
	( 14'sd 6168) * $signed(input_fmap_252[7:0]) +
	( 16'sd 24290) * $signed(input_fmap_253[7:0]) +
	( 16'sd 29146) * $signed(input_fmap_254[7:0]) +
	( 14'sd 5296) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_226;
assign conv_mac_226 = 
	( 13'sd 4003) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26563) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20742) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24548) * $signed(input_fmap_3[7:0]) +
	( 16'sd 17833) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30673) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10199) * $signed(input_fmap_6[7:0]) +
	( 15'sd 15950) * $signed(input_fmap_7[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_8[7:0]) +
	( 15'sd 11931) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9513) * $signed(input_fmap_10[7:0]) +
	( 16'sd 24147) * $signed(input_fmap_11[7:0]) +
	( 16'sd 21758) * $signed(input_fmap_12[7:0]) +
	( 16'sd 30044) * $signed(input_fmap_13[7:0]) +
	( 15'sd 11731) * $signed(input_fmap_14[7:0]) +
	( 14'sd 5446) * $signed(input_fmap_15[7:0]) +
	( 15'sd 10023) * $signed(input_fmap_16[7:0]) +
	( 15'sd 13413) * $signed(input_fmap_17[7:0]) +
	( 14'sd 5628) * $signed(input_fmap_18[7:0]) +
	( 15'sd 10259) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_20[7:0]) +
	( 14'sd 4431) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4961) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1902) * $signed(input_fmap_24[7:0]) +
	( 16'sd 16770) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14932) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20354) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24706) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13854) * $signed(input_fmap_29[7:0]) +
	( 13'sd 4073) * $signed(input_fmap_30[7:0]) +
	( 16'sd 30794) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10322) * $signed(input_fmap_32[7:0]) +
	( 16'sd 21418) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30679) * $signed(input_fmap_34[7:0]) +
	( 16'sd 32374) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32168) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1853) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13544) * $signed(input_fmap_38[7:0]) +
	( 14'sd 4275) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18457) * $signed(input_fmap_40[7:0]) +
	( 16'sd 31038) * $signed(input_fmap_41[7:0]) +
	( 16'sd 31118) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26226) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23032) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21367) * $signed(input_fmap_45[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_46[7:0]) +
	( 15'sd 14273) * $signed(input_fmap_47[7:0]) +
	( 15'sd 13765) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31404) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6667) * $signed(input_fmap_50[7:0]) +
	( 16'sd 31143) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22551) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16999) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27465) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15342) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16889) * $signed(input_fmap_56[7:0]) +
	( 16'sd 25224) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15400) * $signed(input_fmap_58[7:0]) +
	( 16'sd 24825) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11293) * $signed(input_fmap_61[7:0]) +
	( 13'sd 4051) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21647) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20023) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9488) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14465) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13038) * $signed(input_fmap_67[7:0]) +
	( 15'sd 11124) * $signed(input_fmap_68[7:0]) +
	( 15'sd 15209) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30342) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32166) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26932) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4895) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8383) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3105) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24645) * $signed(input_fmap_76[7:0]) +
	( 15'sd 16105) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29161) * $signed(input_fmap_78[7:0]) +
	( 16'sd 19676) * $signed(input_fmap_79[7:0]) +
	( 16'sd 23354) * $signed(input_fmap_80[7:0]) +
	( 13'sd 3777) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3486) * $signed(input_fmap_82[7:0]) +
	( 16'sd 27394) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15329) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31390) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18605) * $signed(input_fmap_86[7:0]) +
	( 16'sd 24735) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19484) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12944) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6657) * $signed(input_fmap_90[7:0]) +
	( 16'sd 31847) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22105) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20782) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26246) * $signed(input_fmap_94[7:0]) +
	( 16'sd 19582) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15116) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17857) * $signed(input_fmap_97[7:0]) +
	( 15'sd 13743) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29614) * $signed(input_fmap_99[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_100[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_101[7:0]) +
	( 15'sd 14501) * $signed(input_fmap_102[7:0]) +
	( 12'sd 2005) * $signed(input_fmap_103[7:0]) +
	( 14'sd 7655) * $signed(input_fmap_104[7:0]) +
	( 16'sd 29006) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27100) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5766) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5064) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29495) * $signed(input_fmap_109[7:0]) +
	( 12'sd 1177) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15119) * $signed(input_fmap_112[7:0]) +
	( 15'sd 11925) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14878) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_115[7:0]) +
	( 14'sd 4585) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23347) * $signed(input_fmap_117[7:0]) +
	( 16'sd 26503) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27543) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18863) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7020) * $signed(input_fmap_121[7:0]) +
	( 15'sd 9016) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10922) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21586) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28637) * $signed(input_fmap_125[7:0]) +
	( 15'sd 11502) * $signed(input_fmap_126[7:0]) +
	( 16'sd 19954) * $signed(input_fmap_127[7:0]) +
	( 16'sd 22298) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5385) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31458) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14131) * $signed(input_fmap_131[7:0]) +
	( 14'sd 6922) * $signed(input_fmap_132[7:0]) +
	( 14'sd 4467) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2890) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31206) * $signed(input_fmap_135[7:0]) +
	( 15'sd 14385) * $signed(input_fmap_136[7:0]) +
	( 15'sd 9555) * $signed(input_fmap_137[7:0]) +
	( 16'sd 30564) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8470) * $signed(input_fmap_139[7:0]) +
	( 15'sd 12581) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31665) * $signed(input_fmap_141[7:0]) +
	( 16'sd 23809) * $signed(input_fmap_142[7:0]) +
	( 15'sd 13212) * $signed(input_fmap_143[7:0]) +
	( 16'sd 26213) * $signed(input_fmap_144[7:0]) +
	( 15'sd 14061) * $signed(input_fmap_145[7:0]) +
	( 14'sd 4864) * $signed(input_fmap_146[7:0]) +
	( 13'sd 3273) * $signed(input_fmap_147[7:0]) +
	( 14'sd 4249) * $signed(input_fmap_148[7:0]) +
	( 14'sd 5257) * $signed(input_fmap_149[7:0]) +
	( 5'sd 13) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30108) * $signed(input_fmap_151[7:0]) +
	( 10'sd 471) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1220) * $signed(input_fmap_153[7:0]) +
	( 11'sd 593) * $signed(input_fmap_154[7:0]) +
	( 16'sd 24458) * $signed(input_fmap_155[7:0]) +
	( 16'sd 27538) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15800) * $signed(input_fmap_157[7:0]) +
	( 16'sd 26903) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27338) * $signed(input_fmap_159[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_160[7:0]) +
	( 16'sd 24103) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29707) * $signed(input_fmap_162[7:0]) +
	( 16'sd 16796) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3577) * $signed(input_fmap_164[7:0]) +
	( 12'sd 1391) * $signed(input_fmap_165[7:0]) +
	( 16'sd 20186) * $signed(input_fmap_166[7:0]) +
	( 14'sd 6801) * $signed(input_fmap_167[7:0]) +
	( 13'sd 2801) * $signed(input_fmap_168[7:0]) +
	( 15'sd 8422) * $signed(input_fmap_169[7:0]) +
	( 16'sd 32498) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31181) * $signed(input_fmap_171[7:0]) +
	( 16'sd 26588) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19019) * $signed(input_fmap_173[7:0]) +
	( 16'sd 28455) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4987) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21028) * $signed(input_fmap_176[7:0]) +
	( 16'sd 32456) * $signed(input_fmap_177[7:0]) +
	( 15'sd 13541) * $signed(input_fmap_178[7:0]) +
	( 16'sd 30883) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15501) * $signed(input_fmap_180[7:0]) +
	( 16'sd 20134) * $signed(input_fmap_181[7:0]) +
	( 15'sd 11049) * $signed(input_fmap_182[7:0]) +
	( 11'sd 590) * $signed(input_fmap_183[7:0]) +
	( 13'sd 3243) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1765) * $signed(input_fmap_185[7:0]) +
	( 16'sd 26639) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5493) * $signed(input_fmap_187[7:0]) +
	( 16'sd 22402) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17492) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20252) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32144) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_192[7:0]) +
	( 16'sd 17761) * $signed(input_fmap_193[7:0]) +
	( 16'sd 23045) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1034) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22869) * $signed(input_fmap_196[7:0]) +
	( 15'sd 9349) * $signed(input_fmap_197[7:0]) +
	( 15'sd 8363) * $signed(input_fmap_198[7:0]) +
	( 16'sd 24192) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6591) * $signed(input_fmap_200[7:0]) +
	( 16'sd 24058) * $signed(input_fmap_201[7:0]) +
	( 16'sd 20510) * $signed(input_fmap_202[7:0]) +
	( 15'sd 13867) * $signed(input_fmap_203[7:0]) +
	( 15'sd 9553) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31081) * $signed(input_fmap_205[7:0]) +
	( 16'sd 18140) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3657) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30414) * $signed(input_fmap_208[7:0]) +
	( 15'sd 8894) * $signed(input_fmap_209[7:0]) +
	( 16'sd 28183) * $signed(input_fmap_210[7:0]) +
	( 16'sd 16867) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24295) * $signed(input_fmap_212[7:0]) +
	( 16'sd 20589) * $signed(input_fmap_213[7:0]) +
	( 15'sd 13028) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6968) * $signed(input_fmap_215[7:0]) +
	( 11'sd 853) * $signed(input_fmap_216[7:0]) +
	( 14'sd 8109) * $signed(input_fmap_217[7:0]) +
	( 16'sd 20486) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21382) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30991) * $signed(input_fmap_220[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5947) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2796) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_224[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_225[7:0]) +
	( 15'sd 9460) * $signed(input_fmap_226[7:0]) +
	( 15'sd 8335) * $signed(input_fmap_227[7:0]) +
	( 14'sd 5534) * $signed(input_fmap_228[7:0]) +
	( 16'sd 22791) * $signed(input_fmap_229[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_230[7:0]) +
	( 16'sd 21724) * $signed(input_fmap_231[7:0]) +
	( 5'sd 15) * $signed(input_fmap_232[7:0]) +
	( 15'sd 13686) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4931) * $signed(input_fmap_234[7:0]) +
	( 13'sd 2529) * $signed(input_fmap_235[7:0]) +
	( 15'sd 9741) * $signed(input_fmap_236[7:0]) +
	( 16'sd 23070) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28551) * $signed(input_fmap_238[7:0]) +
	( 16'sd 27805) * $signed(input_fmap_239[7:0]) +
	( 15'sd 13345) * $signed(input_fmap_240[7:0]) +
	( 16'sd 28812) * $signed(input_fmap_241[7:0]) +
	( 15'sd 16311) * $signed(input_fmap_242[7:0]) +
	( 16'sd 20018) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6568) * $signed(input_fmap_244[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_245[7:0]) +
	( 16'sd 32252) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27367) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17735) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22521) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6692) * $signed(input_fmap_251[7:0]) +
	( 16'sd 16418) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5858) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23980) * $signed(input_fmap_254[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_227;
assign conv_mac_227 = 
	( 16'sd 22302) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24088) * $signed(input_fmap_1[7:0]) +
	( 16'sd 29856) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13838) * $signed(input_fmap_3[7:0]) +
	( 16'sd 27284) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15632) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17954) * $signed(input_fmap_6[7:0]) +
	( 16'sd 28134) * $signed(input_fmap_7[7:0]) +
	( 16'sd 32083) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22557) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19858) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26939) * $signed(input_fmap_11[7:0]) +
	( 16'sd 28311) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10787) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4504) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22255) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10796) * $signed(input_fmap_17[7:0]) +
	( 15'sd 14562) * $signed(input_fmap_18[7:0]) +
	( 15'sd 9801) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18046) * $signed(input_fmap_20[7:0]) +
	( 16'sd 20981) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24153) * $signed(input_fmap_22[7:0]) +
	( 10'sd 351) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27239) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17679) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8937) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17660) * $signed(input_fmap_27[7:0]) +
	( 16'sd 19788) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7129) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25024) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6824) * $signed(input_fmap_31[7:0]) +
	( 16'sd 19321) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1893) * $signed(input_fmap_33[7:0]) +
	( 14'sd 8158) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_35[7:0]) +
	( 16'sd 23922) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24688) * $signed(input_fmap_37[7:0]) +
	( 10'sd 366) * $signed(input_fmap_38[7:0]) +
	( 11'sd 824) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18267) * $signed(input_fmap_40[7:0]) +
	( 16'sd 22828) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12807) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26198) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22707) * $signed(input_fmap_44[7:0]) +
	( 16'sd 30754) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4656) * $signed(input_fmap_46[7:0]) +
	( 14'sd 4915) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19913) * $signed(input_fmap_48[7:0]) +
	( 11'sd 1009) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25928) * $signed(input_fmap_50[7:0]) +
	( 15'sd 8444) * $signed(input_fmap_51[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11212) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9507) * $signed(input_fmap_54[7:0]) +
	( 16'sd 29786) * $signed(input_fmap_55[7:0]) +
	( 13'sd 3951) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5607) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14383) * $signed(input_fmap_58[7:0]) +
	( 12'sd 1726) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25930) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24749) * $signed(input_fmap_61[7:0]) +
	( 15'sd 12629) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10255) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6934) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32406) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3739) * $signed(input_fmap_66[7:0]) +
	( 14'sd 5041) * $signed(input_fmap_67[7:0]) +
	( 16'sd 19452) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20439) * $signed(input_fmap_69[7:0]) +
	( 12'sd 1841) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27846) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25576) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27727) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28650) * $signed(input_fmap_74[7:0]) +
	( 16'sd 23693) * $signed(input_fmap_75[7:0]) +
	( 13'sd 2298) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32631) * $signed(input_fmap_77[7:0]) +
	( 14'sd 6142) * $signed(input_fmap_78[7:0]) +
	( 16'sd 20507) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20281) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25221) * $signed(input_fmap_81[7:0]) +
	( 16'sd 18985) * $signed(input_fmap_82[7:0]) +
	( 16'sd 20980) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11012) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_85[7:0]) +
	( 15'sd 16321) * $signed(input_fmap_86[7:0]) +
	( 16'sd 28396) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17155) * $signed(input_fmap_88[7:0]) +
	( 15'sd 14835) * $signed(input_fmap_89[7:0]) +
	( 16'sd 16663) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15701) * $signed(input_fmap_91[7:0]) +
	( 16'sd 26065) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25811) * $signed(input_fmap_93[7:0]) +
	( 15'sd 16265) * $signed(input_fmap_94[7:0]) +
	( 15'sd 9987) * $signed(input_fmap_95[7:0]) +
	( 16'sd 22234) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8514) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31767) * $signed(input_fmap_99[7:0]) +
	( 16'sd 19497) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12523) * $signed(input_fmap_101[7:0]) +
	( 12'sd 1367) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19470) * $signed(input_fmap_103[7:0]) +
	( 16'sd 25956) * $signed(input_fmap_104[7:0]) +
	( 14'sd 4967) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17817) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13471) * $signed(input_fmap_107[7:0]) +
	( 16'sd 17774) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4130) * $signed(input_fmap_109[7:0]) +
	( 16'sd 19570) * $signed(input_fmap_110[7:0]) +
	( 16'sd 21801) * $signed(input_fmap_111[7:0]) +
	( 10'sd 325) * $signed(input_fmap_112[7:0]) +
	( 13'sd 2545) * $signed(input_fmap_113[7:0]) +
	( 16'sd 21954) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21535) * $signed(input_fmap_115[7:0]) +
	( 16'sd 24491) * $signed(input_fmap_116[7:0]) +
	( 13'sd 2720) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2914) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12367) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10905) * $signed(input_fmap_120[7:0]) +
	( 16'sd 16873) * $signed(input_fmap_121[7:0]) +
	( 15'sd 13503) * $signed(input_fmap_122[7:0]) +
	( 15'sd 9824) * $signed(input_fmap_123[7:0]) +
	( 16'sd 22333) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30874) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17454) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3448) * $signed(input_fmap_127[7:0]) +
	( 15'sd 10617) * $signed(input_fmap_128[7:0]) +
	( 16'sd 20847) * $signed(input_fmap_129[7:0]) +
	( 16'sd 24662) * $signed(input_fmap_130[7:0]) +
	( 15'sd 12070) * $signed(input_fmap_131[7:0]) +
	( 15'sd 13868) * $signed(input_fmap_132[7:0]) +
	( 15'sd 15187) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2636) * $signed(input_fmap_134[7:0]) +
	( 16'sd 16870) * $signed(input_fmap_135[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_136[7:0]) +
	( 13'sd 2072) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19411) * $signed(input_fmap_138[7:0]) +
	( 13'sd 3696) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30410) * $signed(input_fmap_140[7:0]) +
	( 16'sd 23991) * $signed(input_fmap_141[7:0]) +
	( 16'sd 27666) * $signed(input_fmap_142[7:0]) +
	( 16'sd 18753) * $signed(input_fmap_143[7:0]) +
	( 16'sd 23823) * $signed(input_fmap_144[7:0]) +
	( 14'sd 5011) * $signed(input_fmap_145[7:0]) +
	( 15'sd 10292) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21485) * $signed(input_fmap_147[7:0]) +
	( 13'sd 2852) * $signed(input_fmap_148[7:0]) +
	( 16'sd 31783) * $signed(input_fmap_149[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_150[7:0]) +
	( 16'sd 18834) * $signed(input_fmap_151[7:0]) +
	( 13'sd 3647) * $signed(input_fmap_152[7:0]) +
	( 16'sd 29859) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4417) * $signed(input_fmap_154[7:0]) +
	( 16'sd 16739) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10928) * $signed(input_fmap_156[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_157[7:0]) +
	( 16'sd 29219) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32491) * $signed(input_fmap_159[7:0]) +
	( 15'sd 10930) * $signed(input_fmap_160[7:0]) +
	( 16'sd 17891) * $signed(input_fmap_161[7:0]) +
	( 16'sd 32645) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20253) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3591) * $signed(input_fmap_164[7:0]) +
	( 16'sd 16836) * $signed(input_fmap_165[7:0]) +
	( 12'sd 1976) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9681) * $signed(input_fmap_167[7:0]) +
	( 16'sd 30128) * $signed(input_fmap_168[7:0]) +
	( 12'sd 1572) * $signed(input_fmap_169[7:0]) +
	( 15'sd 14098) * $signed(input_fmap_170[7:0]) +
	( 16'sd 29607) * $signed(input_fmap_171[7:0]) +
	( 15'sd 8934) * $signed(input_fmap_172[7:0]) +
	( 16'sd 24783) * $signed(input_fmap_173[7:0]) +
	( 16'sd 17289) * $signed(input_fmap_174[7:0]) +
	( 14'sd 7397) * $signed(input_fmap_175[7:0]) +
	( 15'sd 11941) * $signed(input_fmap_176[7:0]) +
	( 14'sd 8108) * $signed(input_fmap_177[7:0]) +
	( 16'sd 30820) * $signed(input_fmap_178[7:0]) +
	( 14'sd 4805) * $signed(input_fmap_179[7:0]) +
	( 16'sd 31807) * $signed(input_fmap_180[7:0]) +
	( 16'sd 31868) * $signed(input_fmap_181[7:0]) +
	( 15'sd 11365) * $signed(input_fmap_182[7:0]) +
	( 15'sd 8785) * $signed(input_fmap_183[7:0]) +
	( 16'sd 29715) * $signed(input_fmap_184[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_185[7:0]) +
	( 15'sd 15636) * $signed(input_fmap_186[7:0]) +
	( 13'sd 3116) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4189) * $signed(input_fmap_188[7:0]) +
	( 16'sd 29734) * $signed(input_fmap_189[7:0]) +
	( 14'sd 6092) * $signed(input_fmap_190[7:0]) +
	( 16'sd 21768) * $signed(input_fmap_191[7:0]) +
	( 16'sd 22840) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20584) * $signed(input_fmap_193[7:0]) +
	( 15'sd 13058) * $signed(input_fmap_194[7:0]) +
	( 16'sd 30756) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14195) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14093) * $signed(input_fmap_197[7:0]) +
	( 15'sd 16079) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12370) * $signed(input_fmap_199[7:0]) +
	( 15'sd 16157) * $signed(input_fmap_200[7:0]) +
	( 16'sd 23785) * $signed(input_fmap_201[7:0]) +
	( 16'sd 16527) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30008) * $signed(input_fmap_203[7:0]) +
	( 16'sd 23941) * $signed(input_fmap_204[7:0]) +
	( 16'sd 28551) * $signed(input_fmap_205[7:0]) +
	( 14'sd 8025) * $signed(input_fmap_206[7:0]) +
	( 15'sd 8342) * $signed(input_fmap_207[7:0]) +
	( 15'sd 15651) * $signed(input_fmap_208[7:0]) +
	( 15'sd 14213) * $signed(input_fmap_209[7:0]) +
	( 16'sd 22429) * $signed(input_fmap_210[7:0]) +
	( 16'sd 19953) * $signed(input_fmap_211[7:0]) +
	( 16'sd 24372) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29671) * $signed(input_fmap_213[7:0]) +
	( 16'sd 19344) * $signed(input_fmap_214[7:0]) +
	( 13'sd 3850) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17108) * $signed(input_fmap_216[7:0]) +
	( 16'sd 28036) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22690) * $signed(input_fmap_218[7:0]) +
	( 16'sd 28977) * $signed(input_fmap_219[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_220[7:0]) +
	( 16'sd 17484) * $signed(input_fmap_221[7:0]) +
	( 14'sd 6529) * $signed(input_fmap_222[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1163) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2874) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27557) * $signed(input_fmap_226[7:0]) +
	( 16'sd 23784) * $signed(input_fmap_227[7:0]) +
	( 15'sd 15181) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24179) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18149) * $signed(input_fmap_230[7:0]) +
	( 16'sd 20703) * $signed(input_fmap_231[7:0]) +
	( 16'sd 29011) * $signed(input_fmap_232[7:0]) +
	( 13'sd 2400) * $signed(input_fmap_233[7:0]) +
	( 14'sd 5486) * $signed(input_fmap_234[7:0]) +
	( 15'sd 9996) * $signed(input_fmap_235[7:0]) +
	( 16'sd 23756) * $signed(input_fmap_236[7:0]) +
	( 14'sd 5956) * $signed(input_fmap_237[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_238[7:0]) +
	( 16'sd 21438) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18819) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32189) * $signed(input_fmap_241[7:0]) +
	( 15'sd 9775) * $signed(input_fmap_242[7:0]) +
	( 16'sd 30079) * $signed(input_fmap_243[7:0]) +
	( 16'sd 24254) * $signed(input_fmap_244[7:0]) +
	( 16'sd 22764) * $signed(input_fmap_245[7:0]) +
	( 16'sd 16463) * $signed(input_fmap_246[7:0]) +
	( 16'sd 27833) * $signed(input_fmap_247[7:0]) +
	( 16'sd 17410) * $signed(input_fmap_248[7:0]) +
	( 15'sd 9861) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26400) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26416) * $signed(input_fmap_251[7:0]) +
	( 16'sd 18972) * $signed(input_fmap_252[7:0]) +
	( 12'sd 1096) * $signed(input_fmap_253[7:0]) +
	( 15'sd 8894) * $signed(input_fmap_254[7:0]) +
	( 16'sd 19751) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_228;
assign conv_mac_228 = 
	( 16'sd 23867) * $signed(input_fmap_0[7:0]) +
	( 16'sd 24540) * $signed(input_fmap_1[7:0]) +
	( 16'sd 32395) * $signed(input_fmap_2[7:0]) +
	( 13'sd 3597) * $signed(input_fmap_3[7:0]) +
	( 16'sd 31659) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30322) * $signed(input_fmap_5[7:0]) +
	( 16'sd 17854) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6076) * $signed(input_fmap_7[7:0]) +
	( 14'sd 6393) * $signed(input_fmap_8[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_9[7:0]) +
	( 16'sd 28757) * $signed(input_fmap_10[7:0]) +
	( 16'sd 16866) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25312) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15152) * $signed(input_fmap_13[7:0]) +
	( 16'sd 31817) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4197) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3332) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17451) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26463) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28050) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16823) * $signed(input_fmap_20[7:0]) +
	( 15'sd 9695) * $signed(input_fmap_21[7:0]) +
	( 16'sd 30799) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18623) * $signed(input_fmap_23[7:0]) +
	( 16'sd 30389) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8889) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20344) * $signed(input_fmap_26[7:0]) +
	( 12'sd 1342) * $signed(input_fmap_27[7:0]) +
	( 15'sd 15874) * $signed(input_fmap_28[7:0]) +
	( 15'sd 12899) * $signed(input_fmap_29[7:0]) +
	( 16'sd 31669) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18596) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1046) * $signed(input_fmap_32[7:0]) +
	( 14'sd 5329) * $signed(input_fmap_33[7:0]) +
	( 16'sd 21190) * $signed(input_fmap_34[7:0]) +
	( 16'sd 23661) * $signed(input_fmap_35[7:0]) +
	( 15'sd 12505) * $signed(input_fmap_36[7:0]) +
	( 11'sd 526) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3926) * $signed(input_fmap_38[7:0]) +
	( 14'sd 5616) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3819) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11229) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3405) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15303) * $signed(input_fmap_43[7:0]) +
	( 14'sd 5089) * $signed(input_fmap_44[7:0]) +
	( 16'sd 18257) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9595) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15661) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20229) * $signed(input_fmap_48[7:0]) +
	( 13'sd 3909) * $signed(input_fmap_49[7:0]) +
	( 16'sd 20532) * $signed(input_fmap_50[7:0]) +
	( 16'sd 19310) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2302) * $signed(input_fmap_52[7:0]) +
	( 16'sd 25967) * $signed(input_fmap_53[7:0]) +
	( 9'sd 217) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8798) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19950) * $signed(input_fmap_56[7:0]) +
	( 16'sd 28453) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20358) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15837) * $signed(input_fmap_59[7:0]) +
	( 16'sd 24522) * $signed(input_fmap_60[7:0]) +
	( 14'sd 7193) * $signed(input_fmap_61[7:0]) +
	( 16'sd 24841) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2907) * $signed(input_fmap_63[7:0]) +
	( 7'sd 36) * $signed(input_fmap_64[7:0]) +
	( 13'sd 3158) * $signed(input_fmap_65[7:0]) +
	( 16'sd 21906) * $signed(input_fmap_66[7:0]) +
	( 13'sd 3384) * $signed(input_fmap_67[7:0]) +
	( 15'sd 16110) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30947) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24014) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20057) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12649) * $signed(input_fmap_72[7:0]) +
	( 16'sd 30515) * $signed(input_fmap_73[7:0]) +
	( 14'sd 7544) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29357) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12718) * $signed(input_fmap_76[7:0]) +
	( 14'sd 4735) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24018) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11500) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15349) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30767) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1741) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5385) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28203) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31691) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11693) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22975) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17822) * $signed(input_fmap_88[7:0]) +
	( 16'sd 25541) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32378) * $signed(input_fmap_90[7:0]) +
	( 14'sd 7096) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6087) * $signed(input_fmap_92[7:0]) +
	( 14'sd 4778) * $signed(input_fmap_93[7:0]) +
	( 16'sd 26573) * $signed(input_fmap_94[7:0]) +
	( 14'sd 4885) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32311) * $signed(input_fmap_96[7:0]) +
	( 16'sd 20825) * $signed(input_fmap_97[7:0]) +
	( 15'sd 10367) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11814) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16420) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20526) * $signed(input_fmap_101[7:0]) +
	( 16'sd 24788) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1053) * $signed(input_fmap_103[7:0]) +
	( 14'sd 6151) * $signed(input_fmap_104[7:0]) +
	( 16'sd 25829) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1416) * $signed(input_fmap_106[7:0]) +
	( 16'sd 30029) * $signed(input_fmap_107[7:0]) +
	( 16'sd 32677) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6086) * $signed(input_fmap_109[7:0]) +
	( 16'sd 30399) * $signed(input_fmap_110[7:0]) +
	( 15'sd 8930) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24479) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19166) * $signed(input_fmap_113[7:0]) +
	( 16'sd 30761) * $signed(input_fmap_114[7:0]) +
	( 15'sd 8303) * $signed(input_fmap_115[7:0]) +
	( 14'sd 6193) * $signed(input_fmap_116[7:0]) +
	( 16'sd 16728) * $signed(input_fmap_117[7:0]) +
	( 12'sd 1856) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8308) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20801) * $signed(input_fmap_120[7:0]) +
	( 14'sd 6485) * $signed(input_fmap_121[7:0]) +
	( 13'sd 3652) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27001) * $signed(input_fmap_124[7:0]) +
	( 15'sd 11354) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4338) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18494) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9242) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1204) * $signed(input_fmap_129[7:0]) +
	( 13'sd 2498) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13879) * $signed(input_fmap_131[7:0]) +
	( 15'sd 16306) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29803) * $signed(input_fmap_133[7:0]) +
	( 14'sd 5884) * $signed(input_fmap_134[7:0]) +
	( 12'sd 1507) * $signed(input_fmap_135[7:0]) +
	( 16'sd 20627) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24580) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32315) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11835) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1394) * $signed(input_fmap_140[7:0]) +
	( 16'sd 30254) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30805) * $signed(input_fmap_142[7:0]) +
	( 16'sd 29411) * $signed(input_fmap_143[7:0]) +
	( 16'sd 26671) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23031) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21284) * $signed(input_fmap_146[7:0]) +
	( 15'sd 9762) * $signed(input_fmap_147[7:0]) +
	( 15'sd 10050) * $signed(input_fmap_148[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9306) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4250) * $signed(input_fmap_151[7:0]) +
	( 7'sd 33) * $signed(input_fmap_152[7:0]) +
	( 16'sd 24747) * $signed(input_fmap_153[7:0]) +
	( 16'sd 25138) * $signed(input_fmap_154[7:0]) +
	( 14'sd 6126) * $signed(input_fmap_155[7:0]) +
	( 15'sd 10441) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23007) * $signed(input_fmap_157[7:0]) +
	( 16'sd 22214) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_159[7:0]) +
	( 16'sd 19658) * $signed(input_fmap_160[7:0]) +
	( 16'sd 27648) * $signed(input_fmap_161[7:0]) +
	( 16'sd 17952) * $signed(input_fmap_162[7:0]) +
	( 16'sd 19920) * $signed(input_fmap_163[7:0]) +
	( 16'sd 28341) * $signed(input_fmap_164[7:0]) +
	( 14'sd 6748) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30063) * $signed(input_fmap_166[7:0]) +
	( 13'sd 3834) * $signed(input_fmap_167[7:0]) +
	( 16'sd 28594) * $signed(input_fmap_168[7:0]) +
	( 16'sd 22775) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24872) * $signed(input_fmap_170[7:0]) +
	( 16'sd 25040) * $signed(input_fmap_171[7:0]) +
	( 16'sd 20439) * $signed(input_fmap_172[7:0]) +
	( 14'sd 5857) * $signed(input_fmap_173[7:0]) +
	( 16'sd 25697) * $signed(input_fmap_174[7:0]) +
	( 15'sd 10541) * $signed(input_fmap_175[7:0]) +
	( 12'sd 1861) * $signed(input_fmap_176[7:0]) +
	( 16'sd 23830) * $signed(input_fmap_177[7:0]) +
	( 14'sd 5368) * $signed(input_fmap_178[7:0]) +
	( 9'sd 225) * $signed(input_fmap_179[7:0]) +
	( 14'sd 7966) * $signed(input_fmap_180[7:0]) +
	( 16'sd 18218) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6707) * $signed(input_fmap_182[7:0]) +
	( 15'sd 9728) * $signed(input_fmap_183[7:0]) +
	( 16'sd 26938) * $signed(input_fmap_184[7:0]) +
	( 16'sd 16542) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23627) * $signed(input_fmap_186[7:0]) +
	( 15'sd 10476) * $signed(input_fmap_187[7:0]) +
	( 15'sd 12259) * $signed(input_fmap_188[7:0]) +
	( 14'sd 4132) * $signed(input_fmap_189[7:0]) +
	( 16'sd 20695) * $signed(input_fmap_190[7:0]) +
	( 16'sd 23840) * $signed(input_fmap_191[7:0]) +
	( 16'sd 28364) * $signed(input_fmap_192[7:0]) +
	( 15'sd 12599) * $signed(input_fmap_193[7:0]) +
	( 16'sd 26162) * $signed(input_fmap_194[7:0]) +
	( 16'sd 21962) * $signed(input_fmap_195[7:0]) +
	( 16'sd 17739) * $signed(input_fmap_196[7:0]) +
	( 16'sd 18093) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29813) * $signed(input_fmap_198[7:0]) +
	( 15'sd 15187) * $signed(input_fmap_199[7:0]) +
	( 15'sd 16348) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16809) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5458) * $signed(input_fmap_202[7:0]) +
	( 15'sd 16251) * $signed(input_fmap_203[7:0]) +
	( 16'sd 30400) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2251) * $signed(input_fmap_205[7:0]) +
	( 14'sd 7373) * $signed(input_fmap_206[7:0]) +
	( 16'sd 20507) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28700) * $signed(input_fmap_208[7:0]) +
	( 16'sd 23650) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23808) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30175) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19638) * $signed(input_fmap_212[7:0]) +
	( 16'sd 27854) * $signed(input_fmap_213[7:0]) +
	( 16'sd 21213) * $signed(input_fmap_214[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_215[7:0]) +
	( 15'sd 10838) * $signed(input_fmap_216[7:0]) +
	( 16'sd 28660) * $signed(input_fmap_217[7:0]) +
	( 15'sd 14445) * $signed(input_fmap_218[7:0]) +
	( 14'sd 7516) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31516) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15258) * $signed(input_fmap_221[7:0]) +
	( 15'sd 11975) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28184) * $signed(input_fmap_223[7:0]) +
	( 16'sd 23652) * $signed(input_fmap_224[7:0]) +
	( 16'sd 31092) * $signed(input_fmap_225[7:0]) +
	( 15'sd 15244) * $signed(input_fmap_226[7:0]) +
	( 16'sd 29364) * $signed(input_fmap_227[7:0]) +
	( 16'sd 22857) * $signed(input_fmap_228[7:0]) +
	( 16'sd 22588) * $signed(input_fmap_229[7:0]) +
	( 16'sd 20548) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1122) * $signed(input_fmap_231[7:0]) +
	( 16'sd 25878) * $signed(input_fmap_232[7:0]) +
	( 16'sd 17872) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23978) * $signed(input_fmap_234[7:0]) +
	( 16'sd 17405) * $signed(input_fmap_235[7:0]) +
	( 15'sd 11644) * $signed(input_fmap_236[7:0]) +
	( 16'sd 29759) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13698) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31781) * $signed(input_fmap_239[7:0]) +
	( 16'sd 25148) * $signed(input_fmap_240[7:0]) +
	( 15'sd 12001) * $signed(input_fmap_241[7:0]) +
	( 15'sd 14488) * $signed(input_fmap_242[7:0]) +
	( 15'sd 13126) * $signed(input_fmap_243[7:0]) +
	( 16'sd 25487) * $signed(input_fmap_244[7:0]) +
	( 15'sd 9115) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19638) * $signed(input_fmap_246[7:0]) +
	( 16'sd 25785) * $signed(input_fmap_247[7:0]) +
	( 16'sd 32029) * $signed(input_fmap_248[7:0]) +
	( 16'sd 24040) * $signed(input_fmap_249[7:0]) +
	( 16'sd 20325) * $signed(input_fmap_250[7:0]) +
	( 13'sd 3202) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5017) * $signed(input_fmap_252[7:0]) +
	( 14'sd 6079) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9197) * $signed(input_fmap_254[7:0]) +
	( 16'sd 17529) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_229;
assign conv_mac_229 = 
	( 16'sd 31466) * $signed(input_fmap_0[7:0]) +
	( 16'sd 21771) * $signed(input_fmap_1[7:0]) +
	( 15'sd 14802) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18312) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4304) * $signed(input_fmap_4[7:0]) +
	( 16'sd 23973) * $signed(input_fmap_5[7:0]) +
	( 16'sd 19766) * $signed(input_fmap_6[7:0]) +
	( 16'sd 25001) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28003) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24552) * $signed(input_fmap_9[7:0]) +
	( 16'sd 30172) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6188) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23037) * $signed(input_fmap_12[7:0]) +
	( 16'sd 19745) * $signed(input_fmap_13[7:0]) +
	( 16'sd 17448) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25521) * $signed(input_fmap_15[7:0]) +
	( 15'sd 9725) * $signed(input_fmap_16[7:0]) +
	( 15'sd 12143) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29870) * $signed(input_fmap_18[7:0]) +
	( 16'sd 28886) * $signed(input_fmap_19[7:0]) +
	( 14'sd 8001) * $signed(input_fmap_20[7:0]) +
	( 15'sd 14396) * $signed(input_fmap_21[7:0]) +
	( 16'sd 31641) * $signed(input_fmap_22[7:0]) +
	( 14'sd 6452) * $signed(input_fmap_23[7:0]) +
	( 16'sd 28779) * $signed(input_fmap_24[7:0]) +
	( 14'sd 5094) * $signed(input_fmap_25[7:0]) +
	( 16'sd 26290) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22429) * $signed(input_fmap_27[7:0]) +
	( 13'sd 3541) * $signed(input_fmap_28[7:0]) +
	( 14'sd 5754) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9684) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5491) * $signed(input_fmap_31[7:0]) +
	( 14'sd 5262) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26376) * $signed(input_fmap_33[7:0]) +
	( 14'sd 7931) * $signed(input_fmap_34[7:0]) +
	( 14'sd 6100) * $signed(input_fmap_35[7:0]) +
	( 16'sd 21071) * $signed(input_fmap_36[7:0]) +
	( 13'sd 2184) * $signed(input_fmap_37[7:0]) +
	( 13'sd 3006) * $signed(input_fmap_38[7:0]) +
	( 16'sd 19516) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11555) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20528) * $signed(input_fmap_41[7:0]) +
	( 14'sd 5473) * $signed(input_fmap_42[7:0]) +
	( 13'sd 2713) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13549) * $signed(input_fmap_44[7:0]) +
	( 15'sd 9503) * $signed(input_fmap_45[7:0]) +
	( 16'sd 30110) * $signed(input_fmap_46[7:0]) +
	( 16'sd 26238) * $signed(input_fmap_47[7:0]) +
	( 16'sd 32423) * $signed(input_fmap_48[7:0]) +
	( 16'sd 31402) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27650) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14359) * $signed(input_fmap_51[7:0]) +
	( 15'sd 13742) * $signed(input_fmap_52[7:0]) +
	( 14'sd 4363) * $signed(input_fmap_53[7:0]) +
	( 16'sd 18360) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31703) * $signed(input_fmap_55[7:0]) +
	( 14'sd 7110) * $signed(input_fmap_56[7:0]) +
	( 14'sd 4590) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14863) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19635) * $signed(input_fmap_59[7:0]) +
	( 16'sd 29905) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4876) * $signed(input_fmap_61[7:0]) +
	( 16'sd 21765) * $signed(input_fmap_62[7:0]) +
	( 16'sd 20066) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6543) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2621) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17153) * $signed(input_fmap_66[7:0]) +
	( 14'sd 6818) * $signed(input_fmap_67[7:0]) +
	( 16'sd 21939) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21223) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5641) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20221) * $signed(input_fmap_71[7:0]) +
	( 16'sd 25835) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28447) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26789) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8478) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11979) * $signed(input_fmap_76[7:0]) +
	( 16'sd 24738) * $signed(input_fmap_77[7:0]) +
	( 16'sd 17024) * $signed(input_fmap_78[7:0]) +
	( 14'sd 8055) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31345) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17285) * $signed(input_fmap_81[7:0]) +
	( 16'sd 30674) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25142) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11264) * $signed(input_fmap_84[7:0]) +
	( 10'sd 486) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15197) * $signed(input_fmap_86[7:0]) +
	( 16'sd 19086) * $signed(input_fmap_87[7:0]) +
	( 16'sd 18838) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5086) * $signed(input_fmap_89[7:0]) +
	( 16'sd 20678) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8858) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3128) * $signed(input_fmap_92[7:0]) +
	( 16'sd 26699) * $signed(input_fmap_93[7:0]) +
	( 16'sd 22738) * $signed(input_fmap_94[7:0]) +
	( 15'sd 11756) * $signed(input_fmap_95[7:0]) +
	( 16'sd 18666) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12091) * $signed(input_fmap_97[7:0]) +
	( 16'sd 19102) * $signed(input_fmap_98[7:0]) +
	( 15'sd 13583) * $signed(input_fmap_99[7:0]) +
	( 15'sd 10736) * $signed(input_fmap_100[7:0]) +
	( 16'sd 23068) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21748) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10598) * $signed(input_fmap_103[7:0]) +
	( 11'sd 650) * $signed(input_fmap_104[7:0]) +
	( 15'sd 11368) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21989) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16028) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10854) * $signed(input_fmap_108[7:0]) +
	( 14'sd 5205) * $signed(input_fmap_109[7:0]) +
	( 16'sd 18816) * $signed(input_fmap_110[7:0]) +
	( 15'sd 9881) * $signed(input_fmap_111[7:0]) +
	( 13'sd 3268) * $signed(input_fmap_112[7:0]) +
	( 15'sd 15348) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14310) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_115[7:0]) +
	( 13'sd 3881) * $signed(input_fmap_116[7:0]) +
	( 14'sd 6438) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17841) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32659) * $signed(input_fmap_119[7:0]) +
	( 15'sd 15679) * $signed(input_fmap_120[7:0]) +
	( 11'sd 798) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1146) * $signed(input_fmap_122[7:0]) +
	( 16'sd 21367) * $signed(input_fmap_123[7:0]) +
	( 16'sd 21049) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29885) * $signed(input_fmap_125[7:0]) +
	( 16'sd 31467) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4879) * $signed(input_fmap_128[7:0]) +
	( 16'sd 30016) * $signed(input_fmap_129[7:0]) +
	( 15'sd 15871) * $signed(input_fmap_130[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_131[7:0]) +
	( 16'sd 18469) * $signed(input_fmap_132[7:0]) +
	( 14'sd 5077) * $signed(input_fmap_133[7:0]) +
	( 16'sd 22329) * $signed(input_fmap_134[7:0]) +
	( 14'sd 7941) * $signed(input_fmap_135[7:0]) +
	( 12'sd 1594) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12588) * $signed(input_fmap_137[7:0]) +
	( 16'sd 19653) * $signed(input_fmap_138[7:0]) +
	( 10'sd 341) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26172) * $signed(input_fmap_140[7:0]) +
	( 15'sd 16227) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8303) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17460) * $signed(input_fmap_143[7:0]) +
	( 16'sd 32515) * $signed(input_fmap_144[7:0]) +
	( 16'sd 27185) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15919) * $signed(input_fmap_146[7:0]) +
	( 13'sd 2620) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22073) * $signed(input_fmap_148[7:0]) +
	( 16'sd 28036) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_150[7:0]) +
	( 16'sd 32273) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24451) * $signed(input_fmap_152[7:0]) +
	( 15'sd 13373) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31332) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19344) * $signed(input_fmap_155[7:0]) +
	( 16'sd 22046) * $signed(input_fmap_156[7:0]) +
	( 16'sd 17454) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8989) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3951) * $signed(input_fmap_159[7:0]) +
	( 13'sd 4053) * $signed(input_fmap_160[7:0]) +
	( 7'sd 35) * $signed(input_fmap_161[7:0]) +
	( 15'sd 10747) * $signed(input_fmap_162[7:0]) +
	( 12'sd 1862) * $signed(input_fmap_163[7:0]) +
	( 16'sd 25638) * $signed(input_fmap_164[7:0]) +
	( 16'sd 16664) * $signed(input_fmap_165[7:0]) +
	( 14'sd 7052) * $signed(input_fmap_166[7:0]) +
	( 15'sd 10748) * $signed(input_fmap_167[7:0]) +
	( 16'sd 29848) * $signed(input_fmap_168[7:0]) +
	( 16'sd 18500) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5920) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7182) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12784) * $signed(input_fmap_172[7:0]) +
	( 16'sd 20742) * $signed(input_fmap_173[7:0]) +
	( 14'sd 5490) * $signed(input_fmap_174[7:0]) +
	( 13'sd 3423) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7004) * $signed(input_fmap_176[7:0]) +
	( 11'sd 831) * $signed(input_fmap_177[7:0]) +
	( 15'sd 11821) * $signed(input_fmap_178[7:0]) +
	( 16'sd 24125) * $signed(input_fmap_179[7:0]) +
	( 16'sd 24952) * $signed(input_fmap_180[7:0]) +
	( 16'sd 32126) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12700) * $signed(input_fmap_182[7:0]) +
	( 15'sd 8324) * $signed(input_fmap_183[7:0]) +
	( 16'sd 32725) * $signed(input_fmap_184[7:0]) +
	( 16'sd 17763) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17748) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2168) * $signed(input_fmap_187[7:0]) +
	( 15'sd 9711) * $signed(input_fmap_188[7:0]) +
	( 16'sd 23944) * $signed(input_fmap_189[7:0]) +
	( 15'sd 15904) * $signed(input_fmap_190[7:0]) +
	( 15'sd 10632) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29742) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_193[7:0]) +
	( 16'sd 19573) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22793) * $signed(input_fmap_195[7:0]) +
	( 14'sd 5389) * $signed(input_fmap_196[7:0]) +
	( 13'sd 2902) * $signed(input_fmap_197[7:0]) +
	( 16'sd 29773) * $signed(input_fmap_198[7:0]) +
	( 14'sd 7967) * $signed(input_fmap_199[7:0]) +
	( 15'sd 12815) * $signed(input_fmap_200[7:0]) +
	( 16'sd 32190) * $signed(input_fmap_201[7:0]) +
	( 16'sd 24340) * $signed(input_fmap_202[7:0]) +
	( 16'sd 18881) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32595) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11988) * $signed(input_fmap_205[7:0]) +
	( 16'sd 26358) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5900) * $signed(input_fmap_207[7:0]) +
	( 16'sd 19296) * $signed(input_fmap_208[7:0]) +
	( 15'sd 9399) * $signed(input_fmap_209[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_210[7:0]) +
	( 15'sd 9366) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29476) * $signed(input_fmap_212[7:0]) +
	( 16'sd 31383) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15192) * $signed(input_fmap_214[7:0]) +
	( 15'sd 16234) * $signed(input_fmap_215[7:0]) +
	( 15'sd 11280) * $signed(input_fmap_216[7:0]) +
	( 15'sd 14844) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31177) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10981) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21364) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1150) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5314) * $signed(input_fmap_222[7:0]) +
	( 16'sd 21955) * $signed(input_fmap_223[7:0]) +
	( 16'sd 22439) * $signed(input_fmap_224[7:0]) +
	( 13'sd 3127) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27662) * $signed(input_fmap_226[7:0]) +
	( 15'sd 14989) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1868) * $signed(input_fmap_228[7:0]) +
	( 16'sd 23514) * $signed(input_fmap_229[7:0]) +
	( 16'sd 21678) * $signed(input_fmap_230[7:0]) +
	( 14'sd 7994) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8544) * $signed(input_fmap_232[7:0]) +
	( 15'sd 12611) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19891) * $signed(input_fmap_234[7:0]) +
	( 15'sd 8702) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12306) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19722) * $signed(input_fmap_237[7:0]) +
	( 15'sd 10275) * $signed(input_fmap_238[7:0]) +
	( 16'sd 25518) * $signed(input_fmap_239[7:0]) +
	( 15'sd 14906) * $signed(input_fmap_240[7:0]) +
	( 16'sd 30901) * $signed(input_fmap_241[7:0]) +
	( 15'sd 8988) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2164) * $signed(input_fmap_243[7:0]) +
	( 15'sd 8240) * $signed(input_fmap_244[7:0]) +
	( 16'sd 20269) * $signed(input_fmap_245[7:0]) +
	( 15'sd 12625) * $signed(input_fmap_246[7:0]) +
	( 10'sd 317) * $signed(input_fmap_247[7:0]) +
	( 16'sd 27582) * $signed(input_fmap_248[7:0]) +
	( 16'sd 17543) * $signed(input_fmap_249[7:0]) +
	( 16'sd 16628) * $signed(input_fmap_250[7:0]) +
	( 15'sd 8679) * $signed(input_fmap_251[7:0]) +
	( 15'sd 11494) * $signed(input_fmap_252[7:0]) +
	( 15'sd 14645) * $signed(input_fmap_253[7:0]) +
	( 15'sd 13355) * $signed(input_fmap_254[7:0]) +
	( 16'sd 19981) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_230;
assign conv_mac_230 = 
	( 16'sd 23603) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10065) * $signed(input_fmap_1[7:0]) +
	( 15'sd 13720) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25366) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_4[7:0]) +
	( 11'sd 766) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1939) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31477) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9149) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15077) * $signed(input_fmap_9[7:0]) +
	( 16'sd 23121) * $signed(input_fmap_10[7:0]) +
	( 5'sd 11) * $signed(input_fmap_11[7:0]) +
	( 16'sd 27188) * $signed(input_fmap_12[7:0]) +
	( 16'sd 31015) * $signed(input_fmap_13[7:0]) +
	( 16'sd 19725) * $signed(input_fmap_14[7:0]) +
	( 16'sd 17858) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28918) * $signed(input_fmap_16[7:0]) +
	( 15'sd 10119) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29385) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23844) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2827) * $signed(input_fmap_20[7:0]) +
	( 11'sd 595) * $signed(input_fmap_21[7:0]) +
	( 15'sd 16260) * $signed(input_fmap_22[7:0]) +
	( 14'sd 7455) * $signed(input_fmap_23[7:0]) +
	( 15'sd 8800) * $signed(input_fmap_24[7:0]) +
	( 16'sd 31207) * $signed(input_fmap_25[7:0]) +
	( 16'sd 24325) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20190) * $signed(input_fmap_27[7:0]) +
	( 16'sd 31647) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19017) * $signed(input_fmap_29[7:0]) +
	( 16'sd 17975) * $signed(input_fmap_30[7:0]) +
	( 16'sd 32662) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28459) * $signed(input_fmap_32[7:0]) +
	( 16'sd 27259) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10713) * $signed(input_fmap_34[7:0]) +
	( 13'sd 3319) * $signed(input_fmap_35[7:0]) +
	( 15'sd 9637) * $signed(input_fmap_36[7:0]) +
	( 16'sd 20367) * $signed(input_fmap_37[7:0]) +
	( 15'sd 10454) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6149) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23121) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26980) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23362) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_43[7:0]) +
	( 16'sd 25492) * $signed(input_fmap_44[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_45[7:0]) +
	( 15'sd 9054) * $signed(input_fmap_46[7:0]) +
	( 16'sd 21391) * $signed(input_fmap_47[7:0]) +
	( 16'sd 29952) * $signed(input_fmap_48[7:0]) +
	( 15'sd 12225) * $signed(input_fmap_49[7:0]) +
	( 16'sd 21833) * $signed(input_fmap_50[7:0]) +
	( 16'sd 17028) * $signed(input_fmap_51[7:0]) +
	( 16'sd 19018) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32641) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6340) * $signed(input_fmap_54[7:0]) +
	( 7'sd 47) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4231) * $signed(input_fmap_56[7:0]) +
	( 14'sd 7178) * $signed(input_fmap_57[7:0]) +
	( 15'sd 15275) * $signed(input_fmap_58[7:0]) +
	( 15'sd 9375) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11614) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25394) * $signed(input_fmap_61[7:0]) +
	( 16'sd 28094) * $signed(input_fmap_62[7:0]) +
	( 14'sd 5158) * $signed(input_fmap_63[7:0]) +
	( 16'sd 17517) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32071) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30409) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24486) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6863) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7297) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4361) * $signed(input_fmap_70[7:0]) +
	( 16'sd 32399) * $signed(input_fmap_71[7:0]) +
	( 14'sd 4196) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32377) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16677) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29570) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20498) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21674) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4548) * $signed(input_fmap_78[7:0]) +
	( 16'sd 30574) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26886) * $signed(input_fmap_80[7:0]) +
	( 16'sd 16438) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22543) * $signed(input_fmap_82[7:0]) +
	( 16'sd 22342) * $signed(input_fmap_83[7:0]) +
	( 13'sd 2453) * $signed(input_fmap_84[7:0]) +
	( 14'sd 4096) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21281) * $signed(input_fmap_87[7:0]) +
	( 13'sd 2616) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19688) * $signed(input_fmap_89[7:0]) +
	( 15'sd 15596) * $signed(input_fmap_90[7:0]) +
	( 14'sd 6482) * $signed(input_fmap_91[7:0]) +
	( 15'sd 11243) * $signed(input_fmap_92[7:0]) +
	( 16'sd 19072) * $signed(input_fmap_93[7:0]) +
	( 16'sd 23020) * $signed(input_fmap_94[7:0]) +
	( 16'sd 31487) * $signed(input_fmap_95[7:0]) +
	( 15'sd 16102) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27214) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4265) * $signed(input_fmap_98[7:0]) +
	( 16'sd 28155) * $signed(input_fmap_99[7:0]) +
	( 14'sd 5888) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8364) * $signed(input_fmap_101[7:0]) +
	( 16'sd 26128) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19807) * $signed(input_fmap_103[7:0]) +
	( 9'sd 185) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15907) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17719) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23791) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16850) * $signed(input_fmap_108[7:0]) +
	( 16'sd 31353) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12748) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29774) * $signed(input_fmap_111[7:0]) +
	( 15'sd 15214) * $signed(input_fmap_112[7:0]) +
	( 16'sd 29503) * $signed(input_fmap_113[7:0]) +
	( 16'sd 28195) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12145) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22851) * $signed(input_fmap_116[7:0]) +
	( 11'sd 685) * $signed(input_fmap_117[7:0]) +
	( 16'sd 22490) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12986) * $signed(input_fmap_119[7:0]) +
	( 16'sd 29543) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1417) * $signed(input_fmap_121[7:0]) +
	( 13'sd 4084) * $signed(input_fmap_122[7:0]) +
	( 15'sd 8636) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12335) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13167) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_126[7:0]) +
	( 16'sd 16391) * $signed(input_fmap_127[7:0]) +
	( 16'sd 31591) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28531) * $signed(input_fmap_129[7:0]) +
	( 15'sd 9218) * $signed(input_fmap_130[7:0]) +
	( 16'sd 27295) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8525) * $signed(input_fmap_132[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_133[7:0]) +
	( 16'sd 22301) * $signed(input_fmap_134[7:0]) +
	( 15'sd 8437) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2205) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24473) * $signed(input_fmap_137[7:0]) +
	( 16'sd 30608) * $signed(input_fmap_138[7:0]) +
	( 15'sd 10327) * $signed(input_fmap_139[7:0]) +
	( 16'sd 22125) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5433) * $signed(input_fmap_141[7:0]) +
	( 16'sd 31752) * $signed(input_fmap_142[7:0]) +
	( 16'sd 29360) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5370) * $signed(input_fmap_144[7:0]) +
	( 15'sd 9479) * $signed(input_fmap_145[7:0]) +
	( 16'sd 24515) * $signed(input_fmap_146[7:0]) +
	( 16'sd 20995) * $signed(input_fmap_147[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_148[7:0]) +
	( 16'sd 20043) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23502) * $signed(input_fmap_150[7:0]) +
	( 15'sd 16275) * $signed(input_fmap_151[7:0]) +
	( 10'sd 444) * $signed(input_fmap_152[7:0]) +
	( 16'sd 23743) * $signed(input_fmap_153[7:0]) +
	( 14'sd 4935) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22887) * $signed(input_fmap_155[7:0]) +
	( 15'sd 15148) * $signed(input_fmap_156[7:0]) +
	( 16'sd 17556) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4297) * $signed(input_fmap_158[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6853) * $signed(input_fmap_160[7:0]) +
	( 16'sd 24824) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21125) * $signed(input_fmap_162[7:0]) +
	( 15'sd 14035) * $signed(input_fmap_163[7:0]) +
	( 16'sd 21892) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2671) * $signed(input_fmap_165[7:0]) +
	( 14'sd 5957) * $signed(input_fmap_166[7:0]) +
	( 15'sd 14233) * $signed(input_fmap_167[7:0]) +
	( 16'sd 23421) * $signed(input_fmap_168[7:0]) +
	( 16'sd 16566) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28805) * $signed(input_fmap_170[7:0]) +
	( 14'sd 6152) * $signed(input_fmap_171[7:0]) +
	( 13'sd 3530) * $signed(input_fmap_172[7:0]) +
	( 16'sd 30816) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7847) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4436) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21899) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30791) * $signed(input_fmap_177[7:0]) +
	( 13'sd 2799) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25418) * $signed(input_fmap_179[7:0]) +
	( 16'sd 22589) * $signed(input_fmap_180[7:0]) +
	( 16'sd 22880) * $signed(input_fmap_181[7:0]) +
	( 15'sd 8615) * $signed(input_fmap_182[7:0]) +
	( 16'sd 21905) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22122) * $signed(input_fmap_184[7:0]) +
	( 15'sd 15736) * $signed(input_fmap_185[7:0]) +
	( 16'sd 20544) * $signed(input_fmap_186[7:0]) +
	( 15'sd 16244) * $signed(input_fmap_187[7:0]) +
	( 13'sd 2538) * $signed(input_fmap_188[7:0]) +
	( 16'sd 18579) * $signed(input_fmap_189[7:0]) +
	( 16'sd 19805) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29389) * $signed(input_fmap_191[7:0]) +
	( 13'sd 2151) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11242) * $signed(input_fmap_193[7:0]) +
	( 16'sd 24272) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17514) * $signed(input_fmap_195[7:0]) +
	( 16'sd 27991) * $signed(input_fmap_196[7:0]) +
	( 15'sd 8810) * $signed(input_fmap_197[7:0]) +
	( 16'sd 32638) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6906) * $signed(input_fmap_199[7:0]) +
	( 15'sd 11990) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16929) * $signed(input_fmap_201[7:0]) +
	( 15'sd 11285) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21096) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14299) * $signed(input_fmap_204[7:0]) +
	( 15'sd 9699) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9916) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7913) * $signed(input_fmap_207[7:0]) +
	( 16'sd 19110) * $signed(input_fmap_208[7:0]) +
	( 11'sd 828) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3899) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28048) * $signed(input_fmap_211[7:0]) +
	( 16'sd 23611) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29863) * $signed(input_fmap_213[7:0]) +
	( 14'sd 5064) * $signed(input_fmap_214[7:0]) +
	( 15'sd 14533) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18135) * $signed(input_fmap_216[7:0]) +
	( 14'sd 7037) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30128) * $signed(input_fmap_218[7:0]) +
	( 16'sd 16659) * $signed(input_fmap_219[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_220[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14422) * $signed(input_fmap_222[7:0]) +
	( 13'sd 3059) * $signed(input_fmap_223[7:0]) +
	( 13'sd 2138) * $signed(input_fmap_224[7:0]) +
	( 14'sd 7063) * $signed(input_fmap_225[7:0]) +
	( 15'sd 8676) * $signed(input_fmap_226[7:0]) +
	( 14'sd 4520) * $signed(input_fmap_227[7:0]) +
	( 13'sd 3568) * $signed(input_fmap_228[7:0]) +
	( 13'sd 2072) * $signed(input_fmap_229[7:0]) +
	( 11'sd 1001) * $signed(input_fmap_230[7:0]) +
	( 15'sd 8604) * $signed(input_fmap_231[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_232[7:0]) +
	( 16'sd 31239) * $signed(input_fmap_233[7:0]) +
	( 11'sd 628) * $signed(input_fmap_234[7:0]) +
	( 16'sd 23489) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27339) * $signed(input_fmap_236[7:0]) +
	( 12'sd 1323) * $signed(input_fmap_237[7:0]) +
	( 15'sd 14350) * $signed(input_fmap_238[7:0]) +
	( 15'sd 11200) * $signed(input_fmap_239[7:0]) +
	( 14'sd 8116) * $signed(input_fmap_240[7:0]) +
	( 15'sd 9927) * $signed(input_fmap_241[7:0]) +
	( 16'sd 19824) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22814) * $signed(input_fmap_243[7:0]) +
	( 12'sd 1640) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28468) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19671) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11852) * $signed(input_fmap_247[7:0]) +
	( 13'sd 2552) * $signed(input_fmap_248[7:0]) +
	( 15'sd 14679) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6546) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26829) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27175) * $signed(input_fmap_253[7:0]) +
	( 16'sd 18239) * $signed(input_fmap_254[7:0]) +
	( 15'sd 11862) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_231;
assign conv_mac_231 = 
	( 15'sd 9053) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13207) * $signed(input_fmap_1[7:0]) +
	( 15'sd 8310) * $signed(input_fmap_2[7:0]) +
	( 16'sd 24406) * $signed(input_fmap_3[7:0]) +
	( 15'sd 14710) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11127) * $signed(input_fmap_5[7:0]) +
	( 16'sd 29337) * $signed(input_fmap_6[7:0]) +
	( 16'sd 24704) * $signed(input_fmap_7[7:0]) +
	( 13'sd 3157) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25629) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7393) * $signed(input_fmap_10[7:0]) +
	( 14'sd 8161) * $signed(input_fmap_11[7:0]) +
	( 14'sd 7241) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20619) * $signed(input_fmap_13[7:0]) +
	( 16'sd 32131) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21798) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31449) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1436) * $signed(input_fmap_17[7:0]) +
	( 15'sd 10687) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17705) * $signed(input_fmap_19[7:0]) +
	( 15'sd 8943) * $signed(input_fmap_20[7:0]) +
	( 16'sd 24845) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14206) * $signed(input_fmap_22[7:0]) +
	( 16'sd 26779) * $signed(input_fmap_23[7:0]) +
	( 16'sd 21213) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27812) * $signed(input_fmap_25[7:0]) +
	( 16'sd 23104) * $signed(input_fmap_26[7:0]) +
	( 16'sd 23660) * $signed(input_fmap_27[7:0]) +
	( 11'sd 669) * $signed(input_fmap_28[7:0]) +
	( 15'sd 13813) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25201) * $signed(input_fmap_30[7:0]) +
	( 14'sd 6143) * $signed(input_fmap_31[7:0]) +
	( 16'sd 17548) * $signed(input_fmap_32[7:0]) +
	( 16'sd 25642) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19897) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12367) * $signed(input_fmap_35[7:0]) +
	( 16'sd 32170) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25040) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7034) * $signed(input_fmap_38[7:0]) +
	( 15'sd 12423) * $signed(input_fmap_39[7:0]) +
	( 11'sd 557) * $signed(input_fmap_40[7:0]) +
	( 15'sd 13321) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8202) * $signed(input_fmap_42[7:0]) +
	( 16'sd 21073) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11491) * $signed(input_fmap_44[7:0]) +
	( 16'sd 28241) * $signed(input_fmap_45[7:0]) +
	( 12'sd 1098) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13054) * $signed(input_fmap_47[7:0]) +
	( 16'sd 26046) * $signed(input_fmap_48[7:0]) +
	( 16'sd 21272) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26548) * $signed(input_fmap_50[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22576) * $signed(input_fmap_52[7:0]) +
	( 9'sd 136) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1029) * $signed(input_fmap_54[7:0]) +
	( 16'sd 23202) * $signed(input_fmap_55[7:0]) +
	( 16'sd 16644) * $signed(input_fmap_56[7:0]) +
	( 16'sd 30540) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3964) * $signed(input_fmap_58[7:0]) +
	( 15'sd 15160) * $signed(input_fmap_59[7:0]) +
	( 14'sd 4645) * $signed(input_fmap_60[7:0]) +
	( 16'sd 16880) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8519) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21042) * $signed(input_fmap_63[7:0]) +
	( 16'sd 29767) * $signed(input_fmap_64[7:0]) +
	( 11'sd 977) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11704) * $signed(input_fmap_66[7:0]) +
	( 15'sd 15797) * $signed(input_fmap_67[7:0]) +
	( 14'sd 6217) * $signed(input_fmap_68[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_69[7:0]) +
	( 13'sd 3794) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25468) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17342) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7417) * $signed(input_fmap_73[7:0]) +
	( 15'sd 13992) * $signed(input_fmap_74[7:0]) +
	( 15'sd 14565) * $signed(input_fmap_75[7:0]) +
	( 16'sd 24675) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9898) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10826) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7184) * $signed(input_fmap_79[7:0]) +
	( 14'sd 5534) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14705) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28847) * $signed(input_fmap_82[7:0]) +
	( 16'sd 30759) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3737) * $signed(input_fmap_84[7:0]) +
	( 14'sd 5099) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28935) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29301) * $signed(input_fmap_87[7:0]) +
	( 16'sd 28073) * $signed(input_fmap_88[7:0]) +
	( 15'sd 10539) * $signed(input_fmap_89[7:0]) +
	( 15'sd 9474) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19204) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3591) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25761) * $signed(input_fmap_93[7:0]) +
	( 16'sd 18403) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30458) * $signed(input_fmap_95[7:0]) +
	( 16'sd 20757) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19159) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2241) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7236) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23383) * $signed(input_fmap_100[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_101[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_102[7:0]) +
	( 16'sd 21911) * $signed(input_fmap_103[7:0]) +
	( 15'sd 8377) * $signed(input_fmap_104[7:0]) +
	( 15'sd 9386) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27718) * $signed(input_fmap_106[7:0]) +
	( 14'sd 5315) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4109) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29232) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29394) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23453) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22553) * $signed(input_fmap_112[7:0]) +
	( 16'sd 24993) * $signed(input_fmap_113[7:0]) +
	( 14'sd 8008) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31994) * $signed(input_fmap_115[7:0]) +
	( 11'sd 815) * $signed(input_fmap_116[7:0]) +
	( 16'sd 29252) * $signed(input_fmap_117[7:0]) +
	( 16'sd 29118) * $signed(input_fmap_118[7:0]) +
	( 16'sd 16548) * $signed(input_fmap_119[7:0]) +
	( 16'sd 18273) * $signed(input_fmap_120[7:0]) +
	( 14'sd 5390) * $signed(input_fmap_121[7:0]) +
	( 16'sd 29495) * $signed(input_fmap_122[7:0]) +
	( 8'sd 108) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24772) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27861) * $signed(input_fmap_125[7:0]) +
	( 16'sd 24054) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26447) * $signed(input_fmap_127[7:0]) +
	( 15'sd 8453) * $signed(input_fmap_128[7:0]) +
	( 14'sd 6623) * $signed(input_fmap_129[7:0]) +
	( 16'sd 24654) * $signed(input_fmap_130[7:0]) +
	( 15'sd 10277) * $signed(input_fmap_131[7:0]) +
	( 16'sd 30164) * $signed(input_fmap_132[7:0]) +
	( 15'sd 10495) * $signed(input_fmap_133[7:0]) +
	( 15'sd 9593) * $signed(input_fmap_134[7:0]) +
	( 15'sd 10897) * $signed(input_fmap_135[7:0]) +
	( 14'sd 6478) * $signed(input_fmap_136[7:0]) +
	( 16'sd 23815) * $signed(input_fmap_137[7:0]) +
	( 16'sd 30800) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31852) * $signed(input_fmap_139[7:0]) +
	( 16'sd 30885) * $signed(input_fmap_140[7:0]) +
	( 16'sd 21078) * $signed(input_fmap_141[7:0]) +
	( 13'sd 3069) * $signed(input_fmap_142[7:0]) +
	( 16'sd 26279) * $signed(input_fmap_143[7:0]) +
	( 16'sd 26694) * $signed(input_fmap_144[7:0]) +
	( 15'sd 10681) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1346) * $signed(input_fmap_146[7:0]) +
	( 16'sd 16593) * $signed(input_fmap_147[7:0]) +
	( 14'sd 6668) * $signed(input_fmap_148[7:0]) +
	( 15'sd 10759) * $signed(input_fmap_149[7:0]) +
	( 16'sd 30576) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19923) * $signed(input_fmap_151[7:0]) +
	( 15'sd 15189) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4373) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11836) * $signed(input_fmap_154[7:0]) +
	( 16'sd 27929) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25321) * $signed(input_fmap_156[7:0]) +
	( 16'sd 28606) * $signed(input_fmap_157[7:0]) +
	( 15'sd 10203) * $signed(input_fmap_158[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_159[7:0]) +
	( 16'sd 19616) * $signed(input_fmap_160[7:0]) +
	( 16'sd 32159) * $signed(input_fmap_161[7:0]) +
	( 16'sd 20931) * $signed(input_fmap_162[7:0]) +
	( 16'sd 18699) * $signed(input_fmap_163[7:0]) +
	( 15'sd 12847) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22004) * $signed(input_fmap_165[7:0]) +
	( 9'sd 201) * $signed(input_fmap_166[7:0]) +
	( 16'sd 18024) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1473) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26383) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11663) * $signed(input_fmap_170[7:0]) +
	( 16'sd 28356) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19586) * $signed(input_fmap_172[7:0]) +
	( 16'sd 18539) * $signed(input_fmap_173[7:0]) +
	( 16'sd 23809) * $signed(input_fmap_174[7:0]) +
	( 15'sd 13429) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18948) * $signed(input_fmap_176[7:0]) +
	( 16'sd 22021) * $signed(input_fmap_177[7:0]) +
	( 15'sd 15927) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6151) * $signed(input_fmap_179[7:0]) +
	( 14'sd 6927) * $signed(input_fmap_180[7:0]) +
	( 16'sd 26123) * $signed(input_fmap_181[7:0]) +
	( 15'sd 15592) * $signed(input_fmap_182[7:0]) +
	( 16'sd 26676) * $signed(input_fmap_183[7:0]) +
	( 16'sd 23488) * $signed(input_fmap_184[7:0]) +
	( 16'sd 23487) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_186[7:0]) +
	( 16'sd 30596) * $signed(input_fmap_187[7:0]) +
	( 15'sd 16359) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7455) * $signed(input_fmap_189[7:0]) +
	( 15'sd 10332) * $signed(input_fmap_190[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_191[7:0]) +
	( 16'sd 16706) * $signed(input_fmap_192[7:0]) +
	( 15'sd 9174) * $signed(input_fmap_193[7:0]) +
	( 15'sd 8940) * $signed(input_fmap_194[7:0]) +
	( 16'sd 18461) * $signed(input_fmap_195[7:0]) +
	( 16'sd 22342) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21303) * $signed(input_fmap_197[7:0]) +
	( 15'sd 9791) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12959) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13419) * $signed(input_fmap_200[7:0]) +
	( 14'sd 7343) * $signed(input_fmap_201[7:0]) +
	( 14'sd 4241) * $signed(input_fmap_202[7:0]) +
	( 16'sd 28574) * $signed(input_fmap_203[7:0]) +
	( 14'sd 7760) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6040) * $signed(input_fmap_205[7:0]) +
	( 16'sd 20733) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12026) * $signed(input_fmap_207[7:0]) +
	( 16'sd 21954) * $signed(input_fmap_208[7:0]) +
	( 15'sd 15085) * $signed(input_fmap_209[7:0]) +
	( 16'sd 26462) * $signed(input_fmap_210[7:0]) +
	( 15'sd 12491) * $signed(input_fmap_211[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_212[7:0]) +
	( 16'sd 18646) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15536) * $signed(input_fmap_214[7:0]) +
	( 14'sd 8095) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24842) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9894) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28393) * $signed(input_fmap_218[7:0]) +
	( 13'sd 3075) * $signed(input_fmap_219[7:0]) +
	( 11'sd 993) * $signed(input_fmap_220[7:0]) +
	( 14'sd 7064) * $signed(input_fmap_221[7:0]) +
	( 16'sd 30908) * $signed(input_fmap_222[7:0]) +
	( 16'sd 28744) * $signed(input_fmap_223[7:0]) +
	( 11'sd 551) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13015) * $signed(input_fmap_225[7:0]) +
	( 16'sd 16892) * $signed(input_fmap_226[7:0]) +
	( 15'sd 15885) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10956) * $signed(input_fmap_228[7:0]) +
	( 16'sd 22162) * $signed(input_fmap_229[7:0]) +
	( 14'sd 4429) * $signed(input_fmap_230[7:0]) +
	( 16'sd 27659) * $signed(input_fmap_231[7:0]) +
	( 15'sd 9774) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5509) * $signed(input_fmap_233[7:0]) +
	( 13'sd 2175) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29542) * $signed(input_fmap_235[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_236[7:0]) +
	( 16'sd 16431) * $signed(input_fmap_237[7:0]) +
	( 15'sd 11332) * $signed(input_fmap_238[7:0]) +
	( 15'sd 11400) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19500) * $signed(input_fmap_240[7:0]) +
	( 16'sd 26125) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27135) * $signed(input_fmap_242[7:0]) +
	( 15'sd 8593) * $signed(input_fmap_243[7:0]) +
	( 15'sd 10267) * $signed(input_fmap_244[7:0]) +
	( 16'sd 17415) * $signed(input_fmap_245[7:0]) +
	( 16'sd 26533) * $signed(input_fmap_246[7:0]) +
	( 16'sd 19684) * $signed(input_fmap_247[7:0]) +
	( 16'sd 19735) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30176) * $signed(input_fmap_249[7:0]) +
	( 16'sd 19788) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12424) * $signed(input_fmap_251[7:0]) +
	( 16'sd 21072) * $signed(input_fmap_252[7:0]) +
	( 15'sd 8290) * $signed(input_fmap_253[7:0]) +
	( 15'sd 14365) * $signed(input_fmap_254[7:0]) +
	( 15'sd 14897) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_232;
assign conv_mac_232 = 
	( 16'sd 26552) * $signed(input_fmap_0[7:0]) +
	( 16'sd 28386) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18466) * $signed(input_fmap_2[7:0]) +
	( 16'sd 26718) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7651) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11805) * $signed(input_fmap_5[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_6[7:0]) +
	( 15'sd 14950) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15048) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24769) * $signed(input_fmap_9[7:0]) +
	( 15'sd 9394) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2338) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12843) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10027) * $signed(input_fmap_13[7:0]) +
	( 16'sd 20124) * $signed(input_fmap_14[7:0]) +
	( 5'sd 11) * $signed(input_fmap_15[7:0]) +
	( 16'sd 21500) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14019) * $signed(input_fmap_17[7:0]) +
	( 16'sd 29753) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26179) * $signed(input_fmap_19[7:0]) +
	( 12'sd 1282) * $signed(input_fmap_20[7:0]) +
	( 15'sd 15845) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18768) * $signed(input_fmap_22[7:0]) +
	( 15'sd 8395) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14188) * $signed(input_fmap_24[7:0]) +
	( 14'sd 4520) * $signed(input_fmap_25[7:0]) +
	( 15'sd 14837) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3140) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10359) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26767) * $signed(input_fmap_29[7:0]) +
	( 16'sd 16453) * $signed(input_fmap_30[7:0]) +
	( 14'sd 7703) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28321) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3086) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5585) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26645) * $signed(input_fmap_35[7:0]) +
	( 10'sd 363) * $signed(input_fmap_36[7:0]) +
	( 16'sd 19836) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7158) * $signed(input_fmap_38[7:0]) +
	( 15'sd 14676) * $signed(input_fmap_39[7:0]) +
	( 16'sd 19733) * $signed(input_fmap_40[7:0]) +
	( 16'sd 27546) * $signed(input_fmap_41[7:0]) +
	( 16'sd 28931) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26105) * $signed(input_fmap_43[7:0]) +
	( 12'sd 1388) * $signed(input_fmap_44[7:0]) +
	( 13'sd 2985) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21529) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12443) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28050) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5108) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32082) * $signed(input_fmap_50[7:0]) +
	( 14'sd 8111) * $signed(input_fmap_51[7:0]) +
	( 13'sd 3886) * $signed(input_fmap_52[7:0]) +
	( 15'sd 11837) * $signed(input_fmap_53[7:0]) +
	( 14'sd 8163) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24360) * $signed(input_fmap_55[7:0]) +
	( 14'sd 4295) * $signed(input_fmap_56[7:0]) +
	( 16'sd 17216) * $signed(input_fmap_57[7:0]) +
	( 16'sd 21749) * $signed(input_fmap_58[7:0]) +
	( 15'sd 14859) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26208) * $signed(input_fmap_60[7:0]) +
	( 15'sd 10140) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17545) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32737) * $signed(input_fmap_63[7:0]) +
	( 15'sd 12416) * $signed(input_fmap_64[7:0]) +
	( 6'sd 21) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17514) * $signed(input_fmap_66[7:0]) +
	( 16'sd 28848) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24920) * $signed(input_fmap_68[7:0]) +
	( 8'sd 106) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27462) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1557) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26477) * $signed(input_fmap_72[7:0]) +
	( 13'sd 2815) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5220) * $signed(input_fmap_74[7:0]) +
	( 16'sd 27136) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19255) * $signed(input_fmap_76[7:0]) +
	( 16'sd 18631) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18596) * $signed(input_fmap_78[7:0]) +
	( 15'sd 13574) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27666) * $signed(input_fmap_80[7:0]) +
	( 16'sd 25435) * $signed(input_fmap_81[7:0]) +
	( 15'sd 8698) * $signed(input_fmap_82[7:0]) +
	( 13'sd 3304) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9071) * $signed(input_fmap_84[7:0]) +
	( 16'sd 18833) * $signed(input_fmap_85[7:0]) +
	( 16'sd 19877) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22634) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1280) * $signed(input_fmap_88[7:0]) +
	( 14'sd 8005) * $signed(input_fmap_89[7:0]) +
	( 11'sd 831) * $signed(input_fmap_90[7:0]) +
	( 15'sd 8383) * $signed(input_fmap_91[7:0]) +
	( 16'sd 27428) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11496) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2393) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14606) * $signed(input_fmap_95[7:0]) +
	( 16'sd 17985) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11382) * $signed(input_fmap_97[7:0]) +
	( 14'sd 4747) * $signed(input_fmap_98[7:0]) +
	( 14'sd 5864) * $signed(input_fmap_99[7:0]) +
	( 16'sd 23541) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_101[7:0]) +
	( 15'sd 12354) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13363) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12003) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9189) * $signed(input_fmap_106[7:0]) +
	( 16'sd 29575) * $signed(input_fmap_107[7:0]) +
	( 16'sd 16421) * $signed(input_fmap_108[7:0]) +
	( 13'sd 2548) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5823) * $signed(input_fmap_110[7:0]) +
	( 15'sd 12388) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22378) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30679) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15741) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20838) * $signed(input_fmap_115[7:0]) +
	( 15'sd 11214) * $signed(input_fmap_116[7:0]) +
	( 16'sd 31224) * $signed(input_fmap_117[7:0]) +
	( 15'sd 9509) * $signed(input_fmap_118[7:0]) +
	( 16'sd 24870) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10456) * $signed(input_fmap_120[7:0]) +
	( 16'sd 23885) * $signed(input_fmap_121[7:0]) +
	( 16'sd 31798) * $signed(input_fmap_122[7:0]) +
	( 16'sd 30994) * $signed(input_fmap_123[7:0]) +
	( 15'sd 9792) * $signed(input_fmap_124[7:0]) +
	( 16'sd 24929) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12762) * $signed(input_fmap_126[7:0]) +
	( 13'sd 3933) * $signed(input_fmap_127[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_128[7:0]) +
	( 13'sd 3550) * $signed(input_fmap_129[7:0]) +
	( 16'sd 22567) * $signed(input_fmap_130[7:0]) +
	( 16'sd 17750) * $signed(input_fmap_131[7:0]) +
	( 16'sd 22591) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_133[7:0]) +
	( 16'sd 29234) * $signed(input_fmap_134[7:0]) +
	( 14'sd 4867) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15405) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26720) * $signed(input_fmap_137[7:0]) +
	( 13'sd 2132) * $signed(input_fmap_138[7:0]) +
	( 16'sd 23768) * $signed(input_fmap_139[7:0]) +
	( 16'sd 28208) * $signed(input_fmap_140[7:0]) +
	( 14'sd 6310) * $signed(input_fmap_141[7:0]) +
	( 13'sd 2130) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12626) * $signed(input_fmap_143[7:0]) +
	( 15'sd 14115) * $signed(input_fmap_144[7:0]) +
	( 13'sd 3952) * $signed(input_fmap_145[7:0]) +
	( 16'sd 30001) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21910) * $signed(input_fmap_147[7:0]) +
	( 16'sd 29288) * $signed(input_fmap_148[7:0]) +
	( 15'sd 12942) * $signed(input_fmap_149[7:0]) +
	( 14'sd 4644) * $signed(input_fmap_150[7:0]) +
	( 16'sd 22360) * $signed(input_fmap_151[7:0]) +
	( 14'sd 4254) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10368) * $signed(input_fmap_153[7:0]) +
	( 15'sd 8592) * $signed(input_fmap_154[7:0]) +
	( 15'sd 13898) * $signed(input_fmap_155[7:0]) +
	( 16'sd 25749) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15138) * $signed(input_fmap_157[7:0]) +
	( 11'sd 558) * $signed(input_fmap_158[7:0]) +
	( 11'sd 730) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26549) * $signed(input_fmap_160[7:0]) +
	( 16'sd 32428) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2826) * $signed(input_fmap_162[7:0]) +
	( 15'sd 14264) * $signed(input_fmap_163[7:0]) +
	( 16'sd 30732) * $signed(input_fmap_164[7:0]) +
	( 16'sd 26398) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3348) * $signed(input_fmap_166[7:0]) +
	( 15'sd 11406) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9020) * $signed(input_fmap_168[7:0]) +
	( 16'sd 24884) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24249) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7559) * $signed(input_fmap_171[7:0]) +
	( 15'sd 10674) * $signed(input_fmap_172[7:0]) +
	( 14'sd 6434) * $signed(input_fmap_173[7:0]) +
	( 15'sd 15590) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28641) * $signed(input_fmap_175[7:0]) +
	( 16'sd 20542) * $signed(input_fmap_176[7:0]) +
	( 14'sd 7600) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14001) * $signed(input_fmap_178[7:0]) +
	( 16'sd 18478) * $signed(input_fmap_179[7:0]) +
	( 16'sd 29101) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11118) * $signed(input_fmap_181[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17768) * $signed(input_fmap_183[7:0]) +
	( 15'sd 12661) * $signed(input_fmap_184[7:0]) +
	( 16'sd 31842) * $signed(input_fmap_185[7:0]) +
	( 15'sd 13910) * $signed(input_fmap_186[7:0]) +
	( 15'sd 10446) * $signed(input_fmap_187[7:0]) +
	( 12'sd 1375) * $signed(input_fmap_188[7:0]) +
	( 16'sd 21025) * $signed(input_fmap_189[7:0]) +
	( 16'sd 32109) * $signed(input_fmap_190[7:0]) +
	( 13'sd 2884) * $signed(input_fmap_191[7:0]) +
	( 16'sd 30359) * $signed(input_fmap_192[7:0]) +
	( 13'sd 3581) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3459) * $signed(input_fmap_194[7:0]) +
	( 16'sd 17352) * $signed(input_fmap_195[7:0]) +
	( 15'sd 8276) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10500) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10419) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6566) * $signed(input_fmap_199[7:0]) +
	( 16'sd 17204) * $signed(input_fmap_200[7:0]) +
	( 15'sd 8451) * $signed(input_fmap_201[7:0]) +
	( 16'sd 22016) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21853) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4227) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5159) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31451) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3779) * $signed(input_fmap_207[7:0]) +
	( 11'sd 552) * $signed(input_fmap_208[7:0]) +
	( 16'sd 16884) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18543) * $signed(input_fmap_210[7:0]) +
	( 13'sd 3751) * $signed(input_fmap_211[7:0]) +
	( 14'sd 6702) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29714) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31373) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5227) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1263) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30927) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22558) * $signed(input_fmap_218[7:0]) +
	( 16'sd 30165) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30065) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27947) * $signed(input_fmap_221[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_222[7:0]) +
	( 16'sd 17080) * $signed(input_fmap_223[7:0]) +
	( 15'sd 10089) * $signed(input_fmap_224[7:0]) +
	( 14'sd 6787) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10208) * $signed(input_fmap_226[7:0]) +
	( 15'sd 10613) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10587) * $signed(input_fmap_228[7:0]) +
	( 15'sd 9146) * $signed(input_fmap_229[7:0]) +
	( 16'sd 17512) * $signed(input_fmap_230[7:0]) +
	( 16'sd 30169) * $signed(input_fmap_231[7:0]) +
	( 16'sd 21715) * $signed(input_fmap_232[7:0]) +
	( 16'sd 28087) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23354) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12849) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12361) * $signed(input_fmap_236[7:0]) +
	( 14'sd 4548) * $signed(input_fmap_237[7:0]) +
	( 16'sd 26306) * $signed(input_fmap_238[7:0]) +
	( 14'sd 6100) * $signed(input_fmap_239[7:0]) +
	( 13'sd 4079) * $signed(input_fmap_240[7:0]) +
	( 15'sd 14207) * $signed(input_fmap_241[7:0]) +
	( 15'sd 8193) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22667) * $signed(input_fmap_243[7:0]) +
	( 14'sd 4144) * $signed(input_fmap_244[7:0]) +
	( 15'sd 13814) * $signed(input_fmap_245[7:0]) +
	( 12'sd 1760) * $signed(input_fmap_246[7:0]) +
	( 15'sd 13371) * $signed(input_fmap_247[7:0]) +
	( 16'sd 19030) * $signed(input_fmap_248[7:0]) +
	( 14'sd 5661) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12120) * $signed(input_fmap_250[7:0]) +
	( 16'sd 19007) * $signed(input_fmap_251[7:0]) +
	( 16'sd 22569) * $signed(input_fmap_252[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_253[7:0]) +
	( 11'sd 990) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24549) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_233;
assign conv_mac_233 = 
	( 16'sd 26617) * $signed(input_fmap_0[7:0]) +
	( 14'sd 5498) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17984) * $signed(input_fmap_2[7:0]) +
	( 15'sd 13772) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6018) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30414) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3535) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8748) * $signed(input_fmap_7[7:0]) +
	( 15'sd 15713) * $signed(input_fmap_8[7:0]) +
	( 11'sd 929) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20451) * $signed(input_fmap_10[7:0]) +
	( 16'sd 21206) * $signed(input_fmap_11[7:0]) +
	( 11'sd 805) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20205) * $signed(input_fmap_13[7:0]) +
	( 16'sd 26358) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24190) * $signed(input_fmap_15[7:0]) +
	( 12'sd 1530) * $signed(input_fmap_16[7:0]) +
	( 14'sd 7330) * $signed(input_fmap_17[7:0]) +
	( 16'sd 16926) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26815) * $signed(input_fmap_19[7:0]) +
	( 16'sd 17030) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12122) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21150) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2149) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10834) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32741) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16046) * $signed(input_fmap_26[7:0]) +
	( 14'sd 8137) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24199) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22401) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5632) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28682) * $signed(input_fmap_31[7:0]) +
	( 15'sd 10280) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4863) * $signed(input_fmap_33[7:0]) +
	( 16'sd 25024) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22596) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18476) * $signed(input_fmap_36[7:0]) +
	( 15'sd 14872) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7582) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13060) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13716) * $signed(input_fmap_40[7:0]) +
	( 8'sd 113) * $signed(input_fmap_41[7:0]) +
	( 16'sd 25033) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1553) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6947) * $signed(input_fmap_44[7:0]) +
	( 16'sd 25384) * $signed(input_fmap_45[7:0]) +
	( 16'sd 16982) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13399) * $signed(input_fmap_47[7:0]) +
	( 12'sd 1517) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6750) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15271) * $signed(input_fmap_50[7:0]) +
	( 15'sd 13163) * $signed(input_fmap_51[7:0]) +
	( 16'sd 18928) * $signed(input_fmap_52[7:0]) +
	( 16'sd 32169) * $signed(input_fmap_53[7:0]) +
	( 16'sd 17037) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17551) * $signed(input_fmap_55[7:0]) +
	( 16'sd 23965) * $signed(input_fmap_56[7:0]) +
	( 15'sd 12544) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4561) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12153) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6296) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25735) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6377) * $signed(input_fmap_62[7:0]) +
	( 16'sd 26486) * $signed(input_fmap_63[7:0]) +
	( 15'sd 16197) * $signed(input_fmap_64[7:0]) +
	( 16'sd 28739) * $signed(input_fmap_65[7:0]) +
	( 14'sd 8155) * $signed(input_fmap_66[7:0]) +
	( 15'sd 9558) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3785) * $signed(input_fmap_68[7:0]) +
	( 16'sd 21680) * $signed(input_fmap_69[7:0]) +
	( 16'sd 23510) * $signed(input_fmap_70[7:0]) +
	( 15'sd 9259) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2474) * $signed(input_fmap_72[7:0]) +
	( 15'sd 8487) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9080) * $signed(input_fmap_74[7:0]) +
	( 15'sd 15308) * $signed(input_fmap_75[7:0]) +
	( 16'sd 20249) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25434) * $signed(input_fmap_77[7:0]) +
	( 15'sd 10265) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3981) * $signed(input_fmap_79[7:0]) +
	( 16'sd 26245) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2595) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23637) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28854) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11872) * $signed(input_fmap_84[7:0]) +
	( 16'sd 23682) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4209) * $signed(input_fmap_86[7:0]) +
	( 16'sd 22752) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17702) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2396) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6082) * $signed(input_fmap_90[7:0]) +
	( 16'sd 25734) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6086) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21818) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25275) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29583) * $signed(input_fmap_95[7:0]) +
	( 11'sd 882) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28132) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23830) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31128) * $signed(input_fmap_99[7:0]) +
	( 16'sd 18385) * $signed(input_fmap_100[7:0]) +
	( 16'sd 32590) * $signed(input_fmap_101[7:0]) +
	( 16'sd 21413) * $signed(input_fmap_102[7:0]) +
	( 15'sd 9888) * $signed(input_fmap_103[7:0]) +
	( 16'sd 24967) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17264) * $signed(input_fmap_105[7:0]) +
	( 16'sd 19815) * $signed(input_fmap_106[7:0]) +
	( 13'sd 2590) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27533) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21493) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13552) * $signed(input_fmap_110[7:0]) +
	( 13'sd 4036) * $signed(input_fmap_111[7:0]) +
	( 15'sd 11217) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30233) * $signed(input_fmap_113[7:0]) +
	( 16'sd 19979) * $signed(input_fmap_114[7:0]) +
	( 15'sd 13727) * $signed(input_fmap_115[7:0]) +
	( 14'sd 7540) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24043) * $signed(input_fmap_117[7:0]) +
	( 13'sd 2852) * $signed(input_fmap_118[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_119[7:0]) +
	( 16'sd 20199) * $signed(input_fmap_120[7:0]) +
	( 16'sd 27802) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24121) * $signed(input_fmap_122[7:0]) +
	( 16'sd 25958) * $signed(input_fmap_123[7:0]) +
	( 16'sd 16470) * $signed(input_fmap_124[7:0]) +
	( 16'sd 29665) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14814) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7202) * $signed(input_fmap_127[7:0]) +
	( 15'sd 16068) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5145) * $signed(input_fmap_129[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_130[7:0]) +
	( 16'sd 23996) * $signed(input_fmap_131[7:0]) +
	( 15'sd 10525) * $signed(input_fmap_132[7:0]) +
	( 14'sd 6090) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1301) * $signed(input_fmap_134[7:0]) +
	( 15'sd 12904) * $signed(input_fmap_135[7:0]) +
	( 16'sd 18642) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27405) * $signed(input_fmap_137[7:0]) +
	( 16'sd 32680) * $signed(input_fmap_138[7:0]) +
	( 15'sd 16195) * $signed(input_fmap_139[7:0]) +
	( 14'sd 5577) * $signed(input_fmap_140[7:0]) +
	( 16'sd 30573) * $signed(input_fmap_141[7:0]) +
	( 16'sd 30803) * $signed(input_fmap_142[7:0]) +
	( 12'sd 1756) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2718) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_145[7:0]) +
	( 16'sd 27936) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11051) * $signed(input_fmap_147[7:0]) +
	( 15'sd 16016) * $signed(input_fmap_148[7:0]) +
	( 15'sd 15654) * $signed(input_fmap_149[7:0]) +
	( 16'sd 17233) * $signed(input_fmap_150[7:0]) +
	( 12'sd 1789) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_152[7:0]) +
	( 14'sd 6344) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6246) * $signed(input_fmap_154[7:0]) +
	( 15'sd 11274) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20915) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30441) * $signed(input_fmap_157[7:0]) +
	( 16'sd 25267) * $signed(input_fmap_158[7:0]) +
	( 16'sd 31720) * $signed(input_fmap_159[7:0]) +
	( 15'sd 9582) * $signed(input_fmap_160[7:0]) +
	( 16'sd 24944) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2824) * $signed(input_fmap_162[7:0]) +
	( 16'sd 21833) * $signed(input_fmap_163[7:0]) +
	( 9'sd 201) * $signed(input_fmap_164[7:0]) +
	( 16'sd 16777) * $signed(input_fmap_165[7:0]) +
	( 11'sd 787) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7007) * $signed(input_fmap_167[7:0]) +
	( 15'sd 16363) * $signed(input_fmap_168[7:0]) +
	( 16'sd 23696) * $signed(input_fmap_169[7:0]) +
	( 16'sd 21470) * $signed(input_fmap_170[7:0]) +
	( 15'sd 10720) * $signed(input_fmap_171[7:0]) +
	( 14'sd 6389) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23189) * $signed(input_fmap_173[7:0]) +
	( 16'sd 30647) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5000) * $signed(input_fmap_175[7:0]) +
	( 16'sd 26152) * $signed(input_fmap_176[7:0]) +
	( 14'sd 6552) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14934) * $signed(input_fmap_178[7:0]) +
	( 15'sd 10668) * $signed(input_fmap_179[7:0]) +
	( 15'sd 11587) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15144) * $signed(input_fmap_181[7:0]) +
	( 15'sd 14689) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17697) * $signed(input_fmap_183[7:0]) +
	( 16'sd 19680) * $signed(input_fmap_184[7:0]) +
	( 15'sd 10050) * $signed(input_fmap_185[7:0]) +
	( 15'sd 9190) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5871) * $signed(input_fmap_187[7:0]) +
	( 16'sd 24897) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17143) * $signed(input_fmap_189[7:0]) +
	( 16'sd 25587) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3634) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19635) * $signed(input_fmap_192[7:0]) +
	( 13'sd 3662) * $signed(input_fmap_193[7:0]) +
	( 12'sd 2047) * $signed(input_fmap_194[7:0]) +
	( 14'sd 6791) * $signed(input_fmap_195[7:0]) +
	( 13'sd 3254) * $signed(input_fmap_196[7:0]) +
	( 15'sd 12159) * $signed(input_fmap_197[7:0]) +
	( 16'sd 24277) * $signed(input_fmap_198[7:0]) +
	( 16'sd 27231) * $signed(input_fmap_199[7:0]) +
	( 6'sd 31) * $signed(input_fmap_200[7:0]) +
	( 15'sd 13725) * $signed(input_fmap_201[7:0]) +
	( 16'sd 31297) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19941) * $signed(input_fmap_203[7:0]) +
	( 12'sd 1376) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15490) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29178) * $signed(input_fmap_206[7:0]) +
	( 14'sd 5638) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17563) * $signed(input_fmap_208[7:0]) +
	( 16'sd 28797) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18506) * $signed(input_fmap_210[7:0]) +
	( 14'sd 4615) * $signed(input_fmap_211[7:0]) +
	( 9'sd 143) * $signed(input_fmap_212[7:0]) +
	( 16'sd 27388) * $signed(input_fmap_213[7:0]) +
	( 16'sd 19236) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2949) * $signed(input_fmap_215[7:0]) +
	( 16'sd 29488) * $signed(input_fmap_216[7:0]) +
	( 16'sd 30837) * $signed(input_fmap_217[7:0]) +
	( 16'sd 16513) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15726) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30777) * $signed(input_fmap_220[7:0]) +
	( 16'sd 30559) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28325) * $signed(input_fmap_222[7:0]) +
	( 16'sd 31971) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17722) * $signed(input_fmap_224[7:0]) +
	( 16'sd 22670) * $signed(input_fmap_225[7:0]) +
	( 16'sd 24500) * $signed(input_fmap_226[7:0]) +
	( 16'sd 28594) * $signed(input_fmap_227[7:0]) +
	( 16'sd 18343) * $signed(input_fmap_228[7:0]) +
	( 16'sd 31254) * $signed(input_fmap_229[7:0]) +
	( 13'sd 3916) * $signed(input_fmap_230[7:0]) +
	( 13'sd 3311) * $signed(input_fmap_231[7:0]) +
	( 16'sd 16647) * $signed(input_fmap_232[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_233[7:0]) +
	( 14'sd 7504) * $signed(input_fmap_234[7:0]) +
	( 15'sd 14304) * $signed(input_fmap_235[7:0]) +
	( 16'sd 26486) * $signed(input_fmap_236[7:0]) +
	( 11'sd 893) * $signed(input_fmap_237[7:0]) +
	( 13'sd 2885) * $signed(input_fmap_238[7:0]) +
	( 15'sd 9869) * $signed(input_fmap_239[7:0]) +
	( 7'sd 61) * $signed(input_fmap_240[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_241[7:0]) +
	( 16'sd 25826) * $signed(input_fmap_242[7:0]) +
	( 16'sd 27180) * $signed(input_fmap_243[7:0]) +
	( 14'sd 5864) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_245[7:0]) +
	( 15'sd 13092) * $signed(input_fmap_246[7:0]) +
	( 16'sd 22891) * $signed(input_fmap_247[7:0]) +
	( 16'sd 30090) * $signed(input_fmap_248[7:0]) +
	( 16'sd 26089) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7197) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14422) * $signed(input_fmap_251[7:0]) +
	( 16'sd 18211) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27054) * $signed(input_fmap_253[7:0]) +
	( 15'sd 8676) * $signed(input_fmap_254[7:0]) +
	( 16'sd 23929) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_234;
assign conv_mac_234 = 
	( 15'sd 14886) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18161) * $signed(input_fmap_1[7:0]) +
	( 12'sd 1322) * $signed(input_fmap_2[7:0]) +
	( 16'sd 18245) * $signed(input_fmap_3[7:0]) +
	( 16'sd 25694) * $signed(input_fmap_4[7:0]) +
	( 13'sd 2187) * $signed(input_fmap_5[7:0]) +
	( 14'sd 7055) * $signed(input_fmap_6[7:0]) +
	( 16'sd 18961) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12120) * $signed(input_fmap_8[7:0]) +
	( 15'sd 12008) * $signed(input_fmap_9[7:0]) +
	( 11'sd 1015) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17488) * $signed(input_fmap_11[7:0]) +
	( 11'sd 858) * $signed(input_fmap_12[7:0]) +
	( 16'sd 18547) * $signed(input_fmap_13[7:0]) +
	( 16'sd 16655) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1764) * $signed(input_fmap_15[7:0]) +
	( 16'sd 22704) * $signed(input_fmap_16[7:0]) +
	( 12'sd 1984) * $signed(input_fmap_17[7:0]) +
	( 11'sd 991) * $signed(input_fmap_18[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_19[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23677) * $signed(input_fmap_21[7:0]) +
	( 14'sd 5437) * $signed(input_fmap_22[7:0]) +
	( 10'sd 400) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1313) * $signed(input_fmap_24[7:0]) +
	( 16'sd 27436) * $signed(input_fmap_25[7:0]) +
	( 16'sd 16541) * $signed(input_fmap_26[7:0]) +
	( 16'sd 22734) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23081) * $signed(input_fmap_28[7:0]) +
	( 15'sd 14906) * $signed(input_fmap_29[7:0]) +
	( 11'sd 971) * $signed(input_fmap_30[7:0]) +
	( 16'sd 25745) * $signed(input_fmap_31[7:0]) +
	( 14'sd 6173) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8529) * $signed(input_fmap_33[7:0]) +
	( 16'sd 28765) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13770) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31692) * $signed(input_fmap_36[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6518) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23021) * $signed(input_fmap_39[7:0]) +
	( 16'sd 26017) * $signed(input_fmap_40[7:0]) +
	( 14'sd 5167) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1081) * $signed(input_fmap_42[7:0]) +
	( 16'sd 22212) * $signed(input_fmap_43[7:0]) +
	( 16'sd 23854) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21488) * $signed(input_fmap_45[7:0]) +
	( 14'sd 4836) * $signed(input_fmap_46[7:0]) +
	( 15'sd 13496) * $signed(input_fmap_47[7:0]) +
	( 16'sd 20828) * $signed(input_fmap_48[7:0]) +
	( 16'sd 28958) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15646) * $signed(input_fmap_50[7:0]) +
	( 14'sd 5566) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8892) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16011) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23254) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22436) * $signed(input_fmap_55[7:0]) +
	( 15'sd 15473) * $signed(input_fmap_56[7:0]) +
	( 14'sd 6211) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6050) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21745) * $signed(input_fmap_59[7:0]) +
	( 16'sd 31827) * $signed(input_fmap_60[7:0]) +
	( 16'sd 32208) * $signed(input_fmap_61[7:0]) +
	( 16'sd 18257) * $signed(input_fmap_62[7:0]) +
	( 16'sd 27979) * $signed(input_fmap_63[7:0]) +
	( 13'sd 2567) * $signed(input_fmap_64[7:0]) +
	( 15'sd 16246) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14533) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32301) * $signed(input_fmap_67[7:0]) +
	( 16'sd 28753) * $signed(input_fmap_68[7:0]) +
	( 15'sd 10340) * $signed(input_fmap_69[7:0]) +
	( 16'sd 30885) * $signed(input_fmap_70[7:0]) +
	( 16'sd 16964) * $signed(input_fmap_71[7:0]) +
	( 14'sd 6880) * $signed(input_fmap_72[7:0]) +
	( 16'sd 26067) * $signed(input_fmap_73[7:0]) +
	( 16'sd 32570) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7484) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15460) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11410) * $signed(input_fmap_77[7:0]) +
	( 13'sd 2549) * $signed(input_fmap_78[7:0]) +
	( 14'sd 7292) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10421) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32220) * $signed(input_fmap_82[7:0]) +
	( 14'sd 4499) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_84[7:0]) +
	( 12'sd 1085) * $signed(input_fmap_85[7:0]) +
	( 16'sd 23978) * $signed(input_fmap_86[7:0]) +
	( 12'sd 1993) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17333) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2911) * $signed(input_fmap_89[7:0]) +
	( 16'sd 24117) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10656) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6495) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25509) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5487) * $signed(input_fmap_94[7:0]) +
	( 15'sd 10398) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21526) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1634) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28481) * $signed(input_fmap_98[7:0]) +
	( 13'sd 2724) * $signed(input_fmap_99[7:0]) +
	( 16'sd 21757) * $signed(input_fmap_100[7:0]) +
	( 16'sd 27567) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6474) * $signed(input_fmap_102[7:0]) +
	( 16'sd 31006) * $signed(input_fmap_103[7:0]) +
	( 16'sd 31686) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13533) * $signed(input_fmap_105[7:0]) +
	( 16'sd 31341) * $signed(input_fmap_106[7:0]) +
	( 16'sd 16950) * $signed(input_fmap_107[7:0]) +
	( 16'sd 20657) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16600) * $signed(input_fmap_109[7:0]) +
	( 14'sd 5410) * $signed(input_fmap_110[7:0]) +
	( 16'sd 32207) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5151) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19723) * $signed(input_fmap_113[7:0]) +
	( 15'sd 14592) * $signed(input_fmap_114[7:0]) +
	( 16'sd 17539) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12183) * $signed(input_fmap_116[7:0]) +
	( 16'sd 28719) * $signed(input_fmap_117[7:0]) +
	( 15'sd 13402) * $signed(input_fmap_118[7:0]) +
	( 16'sd 21174) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10631) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1516) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5503) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24630) * $signed(input_fmap_123[7:0]) +
	( 12'sd 1798) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9595) * $signed(input_fmap_125[7:0]) +
	( 16'sd 26558) * $signed(input_fmap_126[7:0]) +
	( 16'sd 24745) * $signed(input_fmap_127[7:0]) +
	( 16'sd 27056) * $signed(input_fmap_128[7:0]) +
	( 12'sd 1884) * $signed(input_fmap_129[7:0]) +
	( 16'sd 23808) * $signed(input_fmap_130[7:0]) +
	( 14'sd 4703) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25978) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31501) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3178) * $signed(input_fmap_134[7:0]) +
	( 11'sd 958) * $signed(input_fmap_135[7:0]) +
	( 16'sd 31114) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24289) * $signed(input_fmap_137[7:0]) +
	( 16'sd 20025) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2428) * $signed(input_fmap_139[7:0]) +
	( 15'sd 8631) * $signed(input_fmap_140[7:0]) +
	( 14'sd 6278) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14390) * $signed(input_fmap_142[7:0]) +
	( 15'sd 11088) * $signed(input_fmap_143[7:0]) +
	( 12'sd 1241) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23374) * $signed(input_fmap_145[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_146[7:0]) +
	( 16'sd 28589) * $signed(input_fmap_147[7:0]) +
	( 16'sd 30413) * $signed(input_fmap_148[7:0]) +
	( 16'sd 17060) * $signed(input_fmap_149[7:0]) +
	( 16'sd 31131) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19371) * $signed(input_fmap_151[7:0]) +
	( 16'sd 32378) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17056) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10032) * $signed(input_fmap_154[7:0]) +
	( 16'sd 18894) * $signed(input_fmap_155[7:0]) +
	( 16'sd 26535) * $signed(input_fmap_156[7:0]) +
	( 16'sd 26161) * $signed(input_fmap_157[7:0]) +
	( 14'sd 6243) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27859) * $signed(input_fmap_159[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_160[7:0]) +
	( 15'sd 15220) * $signed(input_fmap_161[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_162[7:0]) +
	( 16'sd 23244) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6743) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19830) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31959) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24206) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1406) * $signed(input_fmap_168[7:0]) +
	( 15'sd 10043) * $signed(input_fmap_169[7:0]) +
	( 15'sd 11347) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31828) * $signed(input_fmap_171[7:0]) +
	( 16'sd 23337) * $signed(input_fmap_172[7:0]) +
	( 12'sd 1324) * $signed(input_fmap_173[7:0]) +
	( 16'sd 23331) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4912) * $signed(input_fmap_175[7:0]) +
	( 16'sd 21356) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18820) * $signed(input_fmap_177[7:0]) +
	( 16'sd 24112) * $signed(input_fmap_178[7:0]) +
	( 16'sd 27587) * $signed(input_fmap_179[7:0]) +
	( 16'sd 25238) * $signed(input_fmap_180[7:0]) +
	( 16'sd 32552) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16750) * $signed(input_fmap_182[7:0]) +
	( 16'sd 31119) * $signed(input_fmap_183[7:0]) +
	( 12'sd 1115) * $signed(input_fmap_184[7:0]) +
	( 15'sd 12513) * $signed(input_fmap_185[7:0]) +
	( 15'sd 15189) * $signed(input_fmap_186[7:0]) +
	( 13'sd 2559) * $signed(input_fmap_187[7:0]) +
	( 16'sd 29446) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7935) * $signed(input_fmap_189[7:0]) +
	( 15'sd 10850) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3992) * $signed(input_fmap_191[7:0]) +
	( 15'sd 14193) * $signed(input_fmap_192[7:0]) +
	( 16'sd 26649) * $signed(input_fmap_193[7:0]) +
	( 16'sd 19466) * $signed(input_fmap_194[7:0]) +
	( 15'sd 15496) * $signed(input_fmap_195[7:0]) +
	( 16'sd 30969) * $signed(input_fmap_196[7:0]) +
	( 15'sd 12387) * $signed(input_fmap_197[7:0]) +
	( 11'sd 963) * $signed(input_fmap_198[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_199[7:0]) +
	( 16'sd 17251) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18873) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2730) * $signed(input_fmap_202[7:0]) +
	( 16'sd 31197) * $signed(input_fmap_203[7:0]) +
	( 10'sd 415) * $signed(input_fmap_204[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12788) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7781) * $signed(input_fmap_207[7:0]) +
	( 16'sd 21522) * $signed(input_fmap_208[7:0]) +
	( 15'sd 8385) * $signed(input_fmap_209[7:0]) +
	( 16'sd 19808) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26870) * $signed(input_fmap_211[7:0]) +
	( 16'sd 25535) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1442) * $signed(input_fmap_213[7:0]) +
	( 13'sd 3551) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6556) * $signed(input_fmap_215[7:0]) +
	( 16'sd 25255) * $signed(input_fmap_216[7:0]) +
	( 16'sd 17530) * $signed(input_fmap_217[7:0]) +
	( 14'sd 6688) * $signed(input_fmap_218[7:0]) +
	( 16'sd 16457) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19623) * $signed(input_fmap_220[7:0]) +
	( 16'sd 26131) * $signed(input_fmap_221[7:0]) +
	( 14'sd 6663) * $signed(input_fmap_222[7:0]) +
	( 16'sd 16452) * $signed(input_fmap_223[7:0]) +
	( 16'sd 26381) * $signed(input_fmap_224[7:0]) +
	( 16'sd 31984) * $signed(input_fmap_225[7:0]) +
	( 16'sd 21419) * $signed(input_fmap_226[7:0]) +
	( 16'sd 32683) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31152) * $signed(input_fmap_228[7:0]) +
	( 16'sd 30120) * $signed(input_fmap_229[7:0]) +
	( 8'sd 123) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14833) * $signed(input_fmap_231[7:0]) +
	( 16'sd 22713) * $signed(input_fmap_232[7:0]) +
	( 13'sd 2788) * $signed(input_fmap_233[7:0]) +
	( 16'sd 18555) * $signed(input_fmap_234[7:0]) +
	( 15'sd 15622) * $signed(input_fmap_235[7:0]) +
	( 16'sd 22555) * $signed(input_fmap_236[7:0]) +
	( 15'sd 8707) * $signed(input_fmap_237[7:0]) +
	( 13'sd 3498) * $signed(input_fmap_238[7:0]) +
	( 16'sd 25178) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1292) * $signed(input_fmap_240[7:0]) +
	( 16'sd 27576) * $signed(input_fmap_241[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_242[7:0]) +
	( 11'sd 788) * $signed(input_fmap_243[7:0]) +
	( 14'sd 6815) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10851) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19161) * $signed(input_fmap_246[7:0]) +
	( 15'sd 14602) * $signed(input_fmap_247[7:0]) +
	( 14'sd 6553) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12265) * $signed(input_fmap_249[7:0]) +
	( 14'sd 4748) * $signed(input_fmap_250[7:0]) +
	( 16'sd 18736) * $signed(input_fmap_251[7:0]) +
	( 12'sd 1881) * $signed(input_fmap_252[7:0]) +
	( 14'sd 4848) * $signed(input_fmap_253[7:0]) +
	( 15'sd 9137) * $signed(input_fmap_254[7:0]) +
	( 16'sd 27109) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_235;
assign conv_mac_235 = 
	( 16'sd 26308) * $signed(input_fmap_0[7:0]) +
	( 14'sd 4677) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15431) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30924) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24805) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26306) * $signed(input_fmap_5[7:0]) +
	( 12'sd 1713) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20670) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12399) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22736) * $signed(input_fmap_9[7:0]) +
	( 16'sd 21211) * $signed(input_fmap_10[7:0]) +
	( 11'sd 952) * $signed(input_fmap_11[7:0]) +
	( 16'sd 20921) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11794) * $signed(input_fmap_13[7:0]) +
	( 13'sd 2572) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3715) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14323) * $signed(input_fmap_16[7:0]) +
	( 15'sd 14982) * $signed(input_fmap_17[7:0]) +
	( 16'sd 23800) * $signed(input_fmap_18[7:0]) +
	( 16'sd 29648) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4825) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16274) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27641) * $signed(input_fmap_22[7:0]) +
	( 15'sd 12115) * $signed(input_fmap_23[7:0]) +
	( 16'sd 22624) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14846) * $signed(input_fmap_25[7:0]) +
	( 16'sd 29572) * $signed(input_fmap_26[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17877) * $signed(input_fmap_28[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_29[7:0]) +
	( 16'sd 25179) * $signed(input_fmap_30[7:0]) +
	( 15'sd 15752) * $signed(input_fmap_31[7:0]) +
	( 16'sd 23498) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8839) * $signed(input_fmap_33[7:0]) +
	( 15'sd 16068) * $signed(input_fmap_34[7:0]) +
	( 16'sd 25006) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19258) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13799) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8588) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29723) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6263) * $signed(input_fmap_40[7:0]) +
	( 16'sd 32622) * $signed(input_fmap_41[7:0]) +
	( 15'sd 16300) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15902) * $signed(input_fmap_43[7:0]) +
	( 15'sd 9416) * $signed(input_fmap_44[7:0]) +
	( 14'sd 7188) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5199) * $signed(input_fmap_46[7:0]) +
	( 15'sd 15462) * $signed(input_fmap_47[7:0]) +
	( 16'sd 27386) * $signed(input_fmap_48[7:0]) +
	( 16'sd 32604) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5543) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15157) * $signed(input_fmap_51[7:0]) +
	( 16'sd 25567) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22556) * $signed(input_fmap_53[7:0]) +
	( 12'sd 1679) * $signed(input_fmap_54[7:0]) +
	( 16'sd 26457) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17317) * $signed(input_fmap_56[7:0]) +
	( 15'sd 9573) * $signed(input_fmap_57[7:0]) +
	( 16'sd 24030) * $signed(input_fmap_58[7:0]) +
	( 16'sd 32427) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25651) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24294) * $signed(input_fmap_61[7:0]) +
	( 11'sd 741) * $signed(input_fmap_62[7:0]) +
	( 16'sd 30616) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28370) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4990) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3325) * $signed(input_fmap_66[7:0]) +
	( 9'sd 221) * $signed(input_fmap_67[7:0]) +
	( 16'sd 27817) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30943) * $signed(input_fmap_69[7:0]) +
	( 16'sd 17477) * $signed(input_fmap_70[7:0]) +
	( 16'sd 28520) * $signed(input_fmap_71[7:0]) +
	( 14'sd 7652) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10925) * $signed(input_fmap_73[7:0]) +
	( 13'sd 3280) * $signed(input_fmap_74[7:0]) +
	( 15'sd 10261) * $signed(input_fmap_75[7:0]) +
	( 11'sd 617) * $signed(input_fmap_76[7:0]) +
	( 16'sd 32196) * $signed(input_fmap_77[7:0]) +
	( 16'sd 26561) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22957) * $signed(input_fmap_79[7:0]) +
	( 11'sd 703) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18221) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2653) * $signed(input_fmap_82[7:0]) +
	( 16'sd 24377) * $signed(input_fmap_83[7:0]) +
	( 16'sd 30741) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22846) * $signed(input_fmap_85[7:0]) +
	( 16'sd 18678) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5863) * $signed(input_fmap_87[7:0]) +
	( 13'sd 4005) * $signed(input_fmap_88[7:0]) +
	( 16'sd 29757) * $signed(input_fmap_89[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_90[7:0]) +
	( 16'sd 30038) * $signed(input_fmap_91[7:0]) +
	( 16'sd 17814) * $signed(input_fmap_92[7:0]) +
	( 16'sd 17991) * $signed(input_fmap_93[7:0]) +
	( 16'sd 29782) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29551) * $signed(input_fmap_95[7:0]) +
	( 15'sd 9395) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27190) * $signed(input_fmap_97[7:0]) +
	( 15'sd 11770) * $signed(input_fmap_98[7:0]) +
	( 16'sd 31915) * $signed(input_fmap_99[7:0]) +
	( 15'sd 14867) * $signed(input_fmap_100[7:0]) +
	( 15'sd 9182) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18451) * $signed(input_fmap_102[7:0]) +
	( 15'sd 8483) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30886) * $signed(input_fmap_105[7:0]) +
	( 16'sd 26222) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13651) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23454) * $signed(input_fmap_108[7:0]) +
	( 14'sd 4351) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9806) * $signed(input_fmap_110[7:0]) +
	( 15'sd 13059) * $signed(input_fmap_111[7:0]) +
	( 16'sd 17262) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26371) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6511) * $signed(input_fmap_114[7:0]) +
	( 15'sd 12696) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9575) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24130) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24843) * $signed(input_fmap_118[7:0]) +
	( 16'sd 18146) * $signed(input_fmap_119[7:0]) +
	( 15'sd 10992) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17711) * $signed(input_fmap_121[7:0]) +
	( 16'sd 24092) * $signed(input_fmap_122[7:0]) +
	( 13'sd 3249) * $signed(input_fmap_123[7:0]) +
	( 16'sd 20980) * $signed(input_fmap_124[7:0]) +
	( 15'sd 10524) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29382) * $signed(input_fmap_126[7:0]) +
	( 15'sd 15022) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17104) * $signed(input_fmap_128[7:0]) +
	( 13'sd 3419) * $signed(input_fmap_129[7:0]) +
	( 16'sd 28315) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24087) * $signed(input_fmap_131[7:0]) +
	( 16'sd 31210) * $signed(input_fmap_132[7:0]) +
	( 14'sd 8041) * $signed(input_fmap_133[7:0]) +
	( 15'sd 13353) * $signed(input_fmap_134[7:0]) +
	( 15'sd 11388) * $signed(input_fmap_135[7:0]) +
	( 15'sd 10060) * $signed(input_fmap_136[7:0]) +
	( 16'sd 17609) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11599) * $signed(input_fmap_138[7:0]) +
	( 15'sd 9754) * $signed(input_fmap_139[7:0]) +
	( 14'sd 7079) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5145) * $signed(input_fmap_141[7:0]) +
	( 15'sd 11801) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23849) * $signed(input_fmap_143[7:0]) +
	( 15'sd 11850) * $signed(input_fmap_144[7:0]) +
	( 15'sd 11848) * $signed(input_fmap_145[7:0]) +
	( 10'sd 359) * $signed(input_fmap_146[7:0]) +
	( 14'sd 5792) * $signed(input_fmap_147[7:0]) +
	( 16'sd 23633) * $signed(input_fmap_148[7:0]) +
	( 16'sd 22451) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21483) * $signed(input_fmap_150[7:0]) +
	( 16'sd 21174) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30648) * $signed(input_fmap_152[7:0]) +
	( 16'sd 25852) * $signed(input_fmap_153[7:0]) +
	( 16'sd 18890) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12900) * $signed(input_fmap_155[7:0]) +
	( 16'sd 21059) * $signed(input_fmap_156[7:0]) +
	( 16'sd 29315) * $signed(input_fmap_157[7:0]) +
	( 16'sd 17850) * $signed(input_fmap_158[7:0]) +
	( 16'sd 26865) * $signed(input_fmap_159[7:0]) +
	( 16'sd 29842) * $signed(input_fmap_160[7:0]) +
	( 12'sd 1890) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24588) * $signed(input_fmap_162[7:0]) +
	( 15'sd 15115) * $signed(input_fmap_163[7:0]) +
	( 16'sd 19205) * $signed(input_fmap_164[7:0]) +
	( 16'sd 29697) * $signed(input_fmap_165[7:0]) +
	( 12'sd 1531) * $signed(input_fmap_166[7:0]) +
	( 15'sd 12451) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6365) * $signed(input_fmap_168[7:0]) +
	( 16'sd 19754) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18986) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7633) * $signed(input_fmap_171[7:0]) +
	( 15'sd 9749) * $signed(input_fmap_172[7:0]) +
	( 15'sd 14192) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32752) * $signed(input_fmap_174[7:0]) +
	( 16'sd 17767) * $signed(input_fmap_175[7:0]) +
	( 16'sd 32111) * $signed(input_fmap_176[7:0]) +
	( 15'sd 11711) * $signed(input_fmap_177[7:0]) +
	( 15'sd 14413) * $signed(input_fmap_178[7:0]) +
	( 16'sd 19126) * $signed(input_fmap_179[7:0]) +
	( 16'sd 31421) * $signed(input_fmap_180[7:0]) +
	( 13'sd 3821) * $signed(input_fmap_181[7:0]) +
	( 13'sd 3295) * $signed(input_fmap_182[7:0]) +
	( 16'sd 22998) * $signed(input_fmap_183[7:0]) +
	( 14'sd 6773) * $signed(input_fmap_184[7:0]) +
	( 12'sd 1041) * $signed(input_fmap_185[7:0]) +
	( 14'sd 7723) * $signed(input_fmap_186[7:0]) +
	( 15'sd 12308) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32503) * $signed(input_fmap_188[7:0]) +
	( 16'sd 30587) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17454) * $signed(input_fmap_190[7:0]) +
	( 16'sd 17577) * $signed(input_fmap_191[7:0]) +
	( 16'sd 27423) * $signed(input_fmap_192[7:0]) +
	( 16'sd 21750) * $signed(input_fmap_193[7:0]) +
	( 16'sd 25305) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5622) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12703) * $signed(input_fmap_196[7:0]) +
	( 16'sd 27028) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2865) * $signed(input_fmap_198[7:0]) +
	( 14'sd 6354) * $signed(input_fmap_199[7:0]) +
	( 15'sd 11953) * $signed(input_fmap_200[7:0]) +
	( 15'sd 9917) * $signed(input_fmap_201[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_202[7:0]) +
	( 15'sd 9762) * $signed(input_fmap_203[7:0]) +
	( 16'sd 25447) * $signed(input_fmap_204[7:0]) +
	( 11'sd 750) * $signed(input_fmap_205[7:0]) +
	( 15'sd 12679) * $signed(input_fmap_206[7:0]) +
	( 16'sd 27236) * $signed(input_fmap_207[7:0]) +
	( 16'sd 28152) * $signed(input_fmap_208[7:0]) +
	( 16'sd 32503) * $signed(input_fmap_209[7:0]) +
	( 16'sd 24690) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6721) * $signed(input_fmap_211[7:0]) +
	( 13'sd 2946) * $signed(input_fmap_212[7:0]) +
	( 16'sd 23568) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7569) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9435) * $signed(input_fmap_215[7:0]) +
	( 15'sd 9414) * $signed(input_fmap_216[7:0]) +
	( 16'sd 22510) * $signed(input_fmap_217[7:0]) +
	( 16'sd 30722) * $signed(input_fmap_218[7:0]) +
	( 16'sd 18362) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31861) * $signed(input_fmap_220[7:0]) +
	( 16'sd 26321) * $signed(input_fmap_221[7:0]) +
	( 16'sd 28282) * $signed(input_fmap_222[7:0]) +
	( 16'sd 25604) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30847) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18502) * $signed(input_fmap_225[7:0]) +
	( 16'sd 17358) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2429) * $signed(input_fmap_227[7:0]) +
	( 15'sd 14028) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8695) * $signed(input_fmap_229[7:0]) +
	( 12'sd 1207) * $signed(input_fmap_230[7:0]) +
	( 9'sd 184) * $signed(input_fmap_231[7:0]) +
	( 16'sd 16560) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18796) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14443) * $signed(input_fmap_234[7:0]) +
	( 16'sd 27615) * $signed(input_fmap_235[7:0]) +
	( 15'sd 15904) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19442) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13971) * $signed(input_fmap_238[7:0]) +
	( 16'sd 25422) * $signed(input_fmap_239[7:0]) +
	( 14'sd 8176) * $signed(input_fmap_240[7:0]) +
	( 16'sd 21983) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15977) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28753) * $signed(input_fmap_243[7:0]) +
	( 16'sd 25090) * $signed(input_fmap_244[7:0]) +
	( 15'sd 13745) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9436) * $signed(input_fmap_246[7:0]) +
	( 16'sd 16739) * $signed(input_fmap_247[7:0]) +
	( 16'sd 29986) * $signed(input_fmap_248[7:0]) +
	( 16'sd 25900) * $signed(input_fmap_249[7:0]) +
	( 16'sd 30719) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27993) * $signed(input_fmap_251[7:0]) +
	( 16'sd 16946) * $signed(input_fmap_252[7:0]) +
	( 16'sd 17073) * $signed(input_fmap_253[7:0]) +
	( 16'sd 17264) * $signed(input_fmap_254[7:0]) +
	( 16'sd 22383) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_236;
assign conv_mac_236 = 
	( 14'sd 6339) * $signed(input_fmap_0[7:0]) +
	( 16'sd 27258) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28343) * $signed(input_fmap_2[7:0]) +
	( 16'sd 30888) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21574) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7374) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8532) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19784) * $signed(input_fmap_7[7:0]) +
	( 14'sd 8054) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7150) * $signed(input_fmap_9[7:0]) +
	( 16'sd 27083) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31138) * $signed(input_fmap_11[7:0]) +
	( 13'sd 2882) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10489) * $signed(input_fmap_13[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2197) * $signed(input_fmap_15[7:0]) +
	( 15'sd 14729) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18017) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6644) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2853) * $signed(input_fmap_19[7:0]) +
	( 13'sd 2362) * $signed(input_fmap_20[7:0]) +
	( 16'sd 23541) * $signed(input_fmap_21[7:0]) +
	( 16'sd 27129) * $signed(input_fmap_22[7:0]) +
	( 15'sd 11443) * $signed(input_fmap_23[7:0]) +
	( 13'sd 3411) * $signed(input_fmap_24[7:0]) +
	( 16'sd 22373) * $signed(input_fmap_25[7:0]) +
	( 11'sd 600) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6494) * $signed(input_fmap_27[7:0]) +
	( 14'sd 4962) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1528) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2077) * $signed(input_fmap_30[7:0]) +
	( 16'sd 28738) * $signed(input_fmap_31[7:0]) +
	( 16'sd 24235) * $signed(input_fmap_32[7:0]) +
	( 16'sd 20399) * $signed(input_fmap_33[7:0]) +
	( 14'sd 8066) * $signed(input_fmap_34[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29247) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25526) * $signed(input_fmap_37[7:0]) +
	( 14'sd 6400) * $signed(input_fmap_38[7:0]) +
	( 13'sd 3317) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18583) * $signed(input_fmap_40[7:0]) +
	( 16'sd 18991) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15417) * $signed(input_fmap_42[7:0]) +
	( 15'sd 16216) * $signed(input_fmap_43[7:0]) +
	( 13'sd 2557) * $signed(input_fmap_44[7:0]) +
	( 16'sd 26555) * $signed(input_fmap_45[7:0]) +
	( 15'sd 10208) * $signed(input_fmap_46[7:0]) +
	( 11'sd 1023) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22266) * $signed(input_fmap_48[7:0]) +
	( 16'sd 16446) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10087) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23749) * $signed(input_fmap_51[7:0]) +
	( 16'sd 22484) * $signed(input_fmap_52[7:0]) +
	( 15'sd 8864) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21451) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19623) * $signed(input_fmap_55[7:0]) +
	( 15'sd 8553) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23895) * $signed(input_fmap_57[7:0]) +
	( 7'sd 39) * $signed(input_fmap_58[7:0]) +
	( 16'sd 25699) * $signed(input_fmap_59[7:0]) +
	( 16'sd 25590) * $signed(input_fmap_60[7:0]) +
	( 16'sd 31701) * $signed(input_fmap_61[7:0]) +
	( 16'sd 20479) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18270) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5227) * $signed(input_fmap_64[7:0]) +
	( 16'sd 17776) * $signed(input_fmap_65[7:0]) +
	( 16'sd 16623) * $signed(input_fmap_66[7:0]) +
	( 15'sd 8348) * $signed(input_fmap_67[7:0]) +
	( 16'sd 31681) * $signed(input_fmap_68[7:0]) +
	( 16'sd 27537) * $signed(input_fmap_69[7:0]) +
	( 10'sd 333) * $signed(input_fmap_70[7:0]) +
	( 14'sd 7868) * $signed(input_fmap_71[7:0]) +
	( 15'sd 15377) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6003) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11160) * $signed(input_fmap_74[7:0]) +
	( 15'sd 9779) * $signed(input_fmap_75[7:0]) +
	( 16'sd 19723) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1094) * $signed(input_fmap_77[7:0]) +
	( 15'sd 12673) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3566) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16407) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1061) * $signed(input_fmap_81[7:0]) +
	( 16'sd 23892) * $signed(input_fmap_82[7:0]) +
	( 16'sd 25955) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6167) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31215) * $signed(input_fmap_85[7:0]) +
	( 16'sd 31436) * $signed(input_fmap_86[7:0]) +
	( 10'sd 385) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6826) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27975) * $signed(input_fmap_89[7:0]) +
	( 16'sd 32154) * $signed(input_fmap_90[7:0]) +
	( 16'sd 19660) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20220) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30743) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20202) * $signed(input_fmap_94[7:0]) +
	( 16'sd 23527) * $signed(input_fmap_95[7:0]) +
	( 15'sd 11902) * $signed(input_fmap_96[7:0]) +
	( 15'sd 8250) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17329) * $signed(input_fmap_98[7:0]) +
	( 15'sd 9335) * $signed(input_fmap_99[7:0]) +
	( 16'sd 28643) * $signed(input_fmap_100[7:0]) +
	( 14'sd 4816) * $signed(input_fmap_101[7:0]) +
	( 16'sd 16397) * $signed(input_fmap_102[7:0]) +
	( 12'sd 1526) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16042) * $signed(input_fmap_104[7:0]) +
	( 15'sd 8914) * $signed(input_fmap_105[7:0]) +
	( 16'sd 23398) * $signed(input_fmap_106[7:0]) +
	( 15'sd 13357) * $signed(input_fmap_107[7:0]) +
	( 16'sd 26994) * $signed(input_fmap_108[7:0]) +
	( 16'sd 18617) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9227) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17097) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22630) * $signed(input_fmap_112[7:0]) +
	( 16'sd 32108) * $signed(input_fmap_113[7:0]) +
	( 16'sd 23036) * $signed(input_fmap_114[7:0]) +
	( 16'sd 25917) * $signed(input_fmap_115[7:0]) +
	( 15'sd 10819) * $signed(input_fmap_116[7:0]) +
	( 15'sd 8450) * $signed(input_fmap_117[7:0]) +
	( 11'sd 689) * $signed(input_fmap_118[7:0]) +
	( 14'sd 4235) * $signed(input_fmap_119[7:0]) +
	( 16'sd 23243) * $signed(input_fmap_120[7:0]) +
	( 16'sd 20311) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4245) * $signed(input_fmap_122[7:0]) +
	( 16'sd 18702) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10570) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25051) * $signed(input_fmap_125[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_126[7:0]) +
	( 3'sd 2) * $signed(input_fmap_127[7:0]) +
	( 16'sd 24484) * $signed(input_fmap_128[7:0]) +
	( 15'sd 13526) * $signed(input_fmap_129[7:0]) +
	( 16'sd 24648) * $signed(input_fmap_130[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_131[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_132[7:0]) +
	( 14'sd 6708) * $signed(input_fmap_133[7:0]) +
	( 16'sd 28342) * $signed(input_fmap_134[7:0]) +
	( 16'sd 19001) * $signed(input_fmap_135[7:0]) +
	( 15'sd 13053) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6170) * $signed(input_fmap_137[7:0]) +
	( 16'sd 30734) * $signed(input_fmap_138[7:0]) +
	( 15'sd 8322) * $signed(input_fmap_139[7:0]) +
	( 16'sd 18839) * $signed(input_fmap_140[7:0]) +
	( 13'sd 2734) * $signed(input_fmap_141[7:0]) +
	( 10'sd 325) * $signed(input_fmap_142[7:0]) +
	( 14'sd 5017) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5178) * $signed(input_fmap_144[7:0]) +
	( 16'sd 26516) * $signed(input_fmap_145[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_146[7:0]) +
	( 15'sd 14800) * $signed(input_fmap_147[7:0]) +
	( 16'sd 32722) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18314) * $signed(input_fmap_149[7:0]) +
	( 16'sd 20609) * $signed(input_fmap_150[7:0]) +
	( 15'sd 14012) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30457) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4406) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31447) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20436) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18045) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6195) * $signed(input_fmap_157[7:0]) +
	( 16'sd 21252) * $signed(input_fmap_158[7:0]) +
	( 15'sd 11222) * $signed(input_fmap_159[7:0]) +
	( 16'sd 18909) * $signed(input_fmap_160[7:0]) +
	( 16'sd 16951) * $signed(input_fmap_161[7:0]) +
	( 14'sd 4360) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2374) * $signed(input_fmap_163[7:0]) +
	( 14'sd 5322) * $signed(input_fmap_164[7:0]) +
	( 16'sd 32253) * $signed(input_fmap_165[7:0]) +
	( 15'sd 9756) * $signed(input_fmap_166[7:0]) +
	( 14'sd 7455) * $signed(input_fmap_167[7:0]) +
	( 13'sd 2223) * $signed(input_fmap_168[7:0]) +
	( 15'sd 8425) * $signed(input_fmap_169[7:0]) +
	( 16'sd 17648) * $signed(input_fmap_170[7:0]) +
	( 13'sd 2749) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31980) * $signed(input_fmap_172[7:0]) +
	( 16'sd 28469) * $signed(input_fmap_173[7:0]) +
	( 15'sd 15252) * $signed(input_fmap_174[7:0]) +
	( 15'sd 13974) * $signed(input_fmap_175[7:0]) +
	( 16'sd 26020) * $signed(input_fmap_176[7:0]) +
	( 16'sd 29358) * $signed(input_fmap_177[7:0]) +
	( 16'sd 22261) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25586) * $signed(input_fmap_179[7:0]) +
	( 16'sd 21083) * $signed(input_fmap_180[7:0]) +
	( 16'sd 19154) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26318) * $signed(input_fmap_182[7:0]) +
	( 10'sd 441) * $signed(input_fmap_183[7:0]) +
	( 15'sd 16042) * $signed(input_fmap_184[7:0]) +
	( 14'sd 6153) * $signed(input_fmap_185[7:0]) +
	( 14'sd 5428) * $signed(input_fmap_186[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_187[7:0]) +
	( 15'sd 15836) * $signed(input_fmap_188[7:0]) +
	( 16'sd 24797) * $signed(input_fmap_189[7:0]) +
	( 16'sd 27675) * $signed(input_fmap_190[7:0]) +
	( 14'sd 6921) * $signed(input_fmap_191[7:0]) +
	( 16'sd 25041) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22738) * $signed(input_fmap_193[7:0]) +
	( 16'sd 28352) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25701) * $signed(input_fmap_195[7:0]) +
	( 15'sd 15725) * $signed(input_fmap_196[7:0]) +
	( 16'sd 18564) * $signed(input_fmap_197[7:0]) +
	( 16'sd 23575) * $signed(input_fmap_198[7:0]) +
	( 12'sd 1520) * $signed(input_fmap_199[7:0]) +
	( 16'sd 19131) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18497) * $signed(input_fmap_201[7:0]) +
	( 14'sd 4555) * $signed(input_fmap_202[7:0]) +
	( 15'sd 9880) * $signed(input_fmap_203[7:0]) +
	( 11'sd 823) * $signed(input_fmap_204[7:0]) +
	( 15'sd 10952) * $signed(input_fmap_205[7:0]) +
	( 16'sd 27022) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12011) * $signed(input_fmap_207[7:0]) +
	( 15'sd 9101) * $signed(input_fmap_208[7:0]) +
	( 16'sd 27192) * $signed(input_fmap_209[7:0]) +
	( 16'sd 31795) * $signed(input_fmap_210[7:0]) +
	( 16'sd 16930) * $signed(input_fmap_211[7:0]) +
	( 15'sd 13333) * $signed(input_fmap_212[7:0]) +
	( 14'sd 5038) * $signed(input_fmap_213[7:0]) +
	( 15'sd 10679) * $signed(input_fmap_214[7:0]) +
	( 15'sd 15338) * $signed(input_fmap_215[7:0]) +
	( 16'sd 18215) * $signed(input_fmap_216[7:0]) +
	( 13'sd 2463) * $signed(input_fmap_217[7:0]) +
	( 16'sd 24303) * $signed(input_fmap_218[7:0]) +
	( 14'sd 8162) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31328) * $signed(input_fmap_220[7:0]) +
	( 16'sd 30534) * $signed(input_fmap_221[7:0]) +
	( 15'sd 13438) * $signed(input_fmap_222[7:0]) +
	( 14'sd 5692) * $signed(input_fmap_223[7:0]) +
	( 16'sd 16385) * $signed(input_fmap_224[7:0]) +
	( 16'sd 18200) * $signed(input_fmap_225[7:0]) +
	( 15'sd 14041) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27552) * $signed(input_fmap_227[7:0]) +
	( 16'sd 31112) * $signed(input_fmap_228[7:0]) +
	( 15'sd 14264) * $signed(input_fmap_229[7:0]) +
	( 15'sd 15598) * $signed(input_fmap_230[7:0]) +
	( 10'sd 344) * $signed(input_fmap_231[7:0]) +
	( 13'sd 2342) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3817) * $signed(input_fmap_233[7:0]) +
	( 10'sd 285) * $signed(input_fmap_234[7:0]) +
	( 16'sd 20792) * $signed(input_fmap_235[7:0]) +
	( 15'sd 8588) * $signed(input_fmap_236[7:0]) +
	( 16'sd 27309) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12399) * $signed(input_fmap_238[7:0]) +
	( 16'sd 24610) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9649) * $signed(input_fmap_240[7:0]) +
	( 16'sd 24522) * $signed(input_fmap_241[7:0]) +
	( 15'sd 10323) * $signed(input_fmap_242[7:0]) +
	( 15'sd 12328) * $signed(input_fmap_243[7:0]) +
	( 15'sd 8951) * $signed(input_fmap_244[7:0]) +
	( 16'sd 28555) * $signed(input_fmap_245[7:0]) +
	( 16'sd 29553) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12328) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21234) * $signed(input_fmap_248[7:0]) +
	( 11'sd 547) * $signed(input_fmap_249[7:0]) +
	( 15'sd 16085) * $signed(input_fmap_250[7:0]) +
	( 16'sd 32353) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4174) * $signed(input_fmap_252[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_253[7:0]) +
	( 15'sd 12758) * $signed(input_fmap_254[7:0]) +
	( 13'sd 2633) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_237;
assign conv_mac_237 = 
	( 14'sd 4298) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32518) * $signed(input_fmap_1[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_2[7:0]) +
	( 15'sd 15808) * $signed(input_fmap_3[7:0]) +
	( 8'sd 106) * $signed(input_fmap_4[7:0]) +
	( 16'sd 21909) * $signed(input_fmap_5[7:0]) +
	( 15'sd 15721) * $signed(input_fmap_6[7:0]) +
	( 16'sd 31665) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17422) * $signed(input_fmap_8[7:0]) +
	( 16'sd 22728) * $signed(input_fmap_9[7:0]) +
	( 16'sd 20752) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10187) * $signed(input_fmap_11[7:0]) +
	( 14'sd 6722) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3434) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7525) * $signed(input_fmap_14[7:0]) +
	( 14'sd 4273) * $signed(input_fmap_15[7:0]) +
	( 15'sd 11337) * $signed(input_fmap_16[7:0]) +
	( 16'sd 30497) * $signed(input_fmap_17[7:0]) +
	( 16'sd 26335) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13484) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23896) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21286) * $signed(input_fmap_21[7:0]) +
	( 14'sd 6156) * $signed(input_fmap_22[7:0]) +
	( 15'sd 16354) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1897) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12619) * $signed(input_fmap_25[7:0]) +
	( 14'sd 4432) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26225) * $signed(input_fmap_27[7:0]) +
	( 16'sd 24595) * $signed(input_fmap_28[7:0]) +
	( 14'sd 6544) * $signed(input_fmap_29[7:0]) +
	( 14'sd 4463) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1512) * $signed(input_fmap_31[7:0]) +
	( 14'sd 4744) * $signed(input_fmap_32[7:0]) +
	( 15'sd 10414) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24415) * $signed(input_fmap_34[7:0]) +
	( 16'sd 22611) * $signed(input_fmap_35[7:0]) +
	( 14'sd 5347) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3474) * $signed(input_fmap_37[7:0]) +
	( 15'sd 14829) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29160) * $signed(input_fmap_39[7:0]) +
	( 16'sd 23505) * $signed(input_fmap_40[7:0]) +
	( 15'sd 8287) * $signed(input_fmap_41[7:0]) +
	( 15'sd 8728) * $signed(input_fmap_42[7:0]) +
	( 15'sd 10177) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3068) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15539) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24269) * $signed(input_fmap_46[7:0]) +
	( 16'sd 32079) * $signed(input_fmap_47[7:0]) +
	( 16'sd 30445) * $signed(input_fmap_48[7:0]) +
	( 15'sd 16265) * $signed(input_fmap_49[7:0]) +
	( 16'sd 25432) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30942) * $signed(input_fmap_51[7:0]) +
	( 13'sd 2329) * $signed(input_fmap_52[7:0]) +
	( 15'sd 14358) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27606) * $signed(input_fmap_54[7:0]) +
	( 16'sd 25839) * $signed(input_fmap_55[7:0]) +
	( 15'sd 10393) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24684) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29645) * $signed(input_fmap_58[7:0]) +
	( 14'sd 4741) * $signed(input_fmap_59[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_60[7:0]) +
	( 8'sd 124) * $signed(input_fmap_61[7:0]) +
	( 14'sd 6069) * $signed(input_fmap_62[7:0]) +
	( 12'sd 1665) * $signed(input_fmap_63[7:0]) +
	( 13'sd 3303) * $signed(input_fmap_64[7:0]) +
	( 15'sd 9835) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26637) * $signed(input_fmap_66[7:0]) +
	( 16'sd 24116) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9845) * $signed(input_fmap_68[7:0]) +
	( 15'sd 13284) * $signed(input_fmap_69[7:0]) +
	( 15'sd 10914) * $signed(input_fmap_70[7:0]) +
	( 16'sd 23320) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17414) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11128) * $signed(input_fmap_73[7:0]) +
	( 15'sd 11943) * $signed(input_fmap_74[7:0]) +
	( 16'sd 17206) * $signed(input_fmap_75[7:0]) +
	( 16'sd 21498) * $signed(input_fmap_76[7:0]) +
	( 16'sd 23651) * $signed(input_fmap_77[7:0]) +
	( 14'sd 5865) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27018) * $signed(input_fmap_79[7:0]) +
	( 11'sd 659) * $signed(input_fmap_80[7:0]) +
	( 16'sd 30510) * $signed(input_fmap_81[7:0]) +
	( 16'sd 20591) * $signed(input_fmap_82[7:0]) +
	( 16'sd 31889) * $signed(input_fmap_83[7:0]) +
	( 16'sd 31930) * $signed(input_fmap_84[7:0]) +
	( 16'sd 27345) * $signed(input_fmap_85[7:0]) +
	( 12'sd 1893) * $signed(input_fmap_86[7:0]) +
	( 15'sd 8987) * $signed(input_fmap_87[7:0]) +
	( 15'sd 11324) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28344) * $signed(input_fmap_89[7:0]) +
	( 15'sd 12774) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11211) * $signed(input_fmap_91[7:0]) +
	( 16'sd 23882) * $signed(input_fmap_92[7:0]) +
	( 12'sd 2022) * $signed(input_fmap_93[7:0]) +
	( 16'sd 25838) * $signed(input_fmap_94[7:0]) +
	( 16'sd 28601) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4414) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27145) * $signed(input_fmap_97[7:0]) +
	( 15'sd 12134) * $signed(input_fmap_98[7:0]) +
	( 16'sd 24917) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7340) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28454) * $signed(input_fmap_101[7:0]) +
	( 16'sd 22804) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19485) * $signed(input_fmap_103[7:0]) +
	( 15'sd 16185) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21621) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24988) * $signed(input_fmap_106[7:0]) +
	( 16'sd 24280) * $signed(input_fmap_107[7:0]) +
	( 15'sd 10110) * $signed(input_fmap_108[7:0]) +
	( 15'sd 13102) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11596) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5438) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27125) * $signed(input_fmap_112[7:0]) +
	( 9'sd 201) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27841) * $signed(input_fmap_114[7:0]) +
	( 14'sd 4942) * $signed(input_fmap_115[7:0]) +
	( 15'sd 9831) * $signed(input_fmap_116[7:0]) +
	( 14'sd 4764) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18911) * $signed(input_fmap_118[7:0]) +
	( 7'sd 43) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8424) * $signed(input_fmap_120[7:0]) +
	( 15'sd 12524) * $signed(input_fmap_121[7:0]) +
	( 16'sd 17464) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22241) * $signed(input_fmap_123[7:0]) +
	( 13'sd 2772) * $signed(input_fmap_124[7:0]) +
	( 16'sd 23504) * $signed(input_fmap_125[7:0]) +
	( 16'sd 21475) * $signed(input_fmap_126[7:0]) +
	( 15'sd 11678) * $signed(input_fmap_127[7:0]) +
	( 16'sd 19127) * $signed(input_fmap_128[7:0]) +
	( 11'sd 531) * $signed(input_fmap_129[7:0]) +
	( 15'sd 9624) * $signed(input_fmap_130[7:0]) +
	( 15'sd 13908) * $signed(input_fmap_131[7:0]) +
	( 16'sd 32656) * $signed(input_fmap_132[7:0]) +
	( 11'sd 609) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1143) * $signed(input_fmap_134[7:0]) +
	( 15'sd 15776) * $signed(input_fmap_135[7:0]) +
	( 15'sd 15073) * $signed(input_fmap_136[7:0]) +
	( 14'sd 8051) * $signed(input_fmap_137[7:0]) +
	( 15'sd 10185) * $signed(input_fmap_138[7:0]) +
	( 14'sd 7736) * $signed(input_fmap_139[7:0]) +
	( 14'sd 4600) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19558) * $signed(input_fmap_141[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7692) * $signed(input_fmap_143[7:0]) +
	( 16'sd 30594) * $signed(input_fmap_144[7:0]) +
	( 14'sd 6803) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1890) * $signed(input_fmap_146[7:0]) +
	( 16'sd 17964) * $signed(input_fmap_147[7:0]) +
	( 13'sd 2201) * $signed(input_fmap_148[7:0]) +
	( 16'sd 23666) * $signed(input_fmap_149[7:0]) +
	( 11'sd 910) * $signed(input_fmap_150[7:0]) +
	( 14'sd 7228) * $signed(input_fmap_151[7:0]) +
	( 16'sd 28323) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11710) * $signed(input_fmap_153[7:0]) +
	( 16'sd 24642) * $signed(input_fmap_154[7:0]) +
	( 14'sd 7479) * $signed(input_fmap_155[7:0]) +
	( 10'sd 491) * $signed(input_fmap_156[7:0]) +
	( 14'sd 6145) * $signed(input_fmap_157[7:0]) +
	( 16'sd 23484) * $signed(input_fmap_158[7:0]) +
	( 14'sd 5063) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_160[7:0]) +
	( 16'sd 31431) * $signed(input_fmap_161[7:0]) +
	( 16'sd 25423) * $signed(input_fmap_162[7:0]) +
	( 16'sd 30153) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_164[7:0]) +
	( 13'sd 2122) * $signed(input_fmap_165[7:0]) +
	( 14'sd 6983) * $signed(input_fmap_166[7:0]) +
	( 16'sd 29003) * $signed(input_fmap_167[7:0]) +
	( 14'sd 7820) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11042) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18580) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16861) * $signed(input_fmap_171[7:0]) +
	( 16'sd 28427) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29363) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7174) * $signed(input_fmap_174[7:0]) +
	( 16'sd 30528) * $signed(input_fmap_175[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2836) * $signed(input_fmap_177[7:0]) +
	( 15'sd 12725) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22811) * $signed(input_fmap_179[7:0]) +
	( 13'sd 2394) * $signed(input_fmap_180[7:0]) +
	( 15'sd 16291) * $signed(input_fmap_181[7:0]) +
	( 15'sd 15097) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17105) * $signed(input_fmap_183[7:0]) +
	( 16'sd 28680) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11038) * $signed(input_fmap_185[7:0]) +
	( 15'sd 10567) * $signed(input_fmap_186[7:0]) +
	( 16'sd 28664) * $signed(input_fmap_187[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_188[7:0]) +
	( 16'sd 22856) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4889) * $signed(input_fmap_190[7:0]) +
	( 16'sd 25121) * $signed(input_fmap_191[7:0]) +
	( 16'sd 23142) * $signed(input_fmap_192[7:0]) +
	( 14'sd 4262) * $signed(input_fmap_193[7:0]) +
	( 14'sd 7846) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22554) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19353) * $signed(input_fmap_196[7:0]) +
	( 16'sd 31666) * $signed(input_fmap_197[7:0]) +
	( 16'sd 20737) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5887) * $signed(input_fmap_199[7:0]) +
	( 16'sd 32088) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22216) * $signed(input_fmap_201[7:0]) +
	( 16'sd 22498) * $signed(input_fmap_202[7:0]) +
	( 16'sd 25592) * $signed(input_fmap_203[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_204[7:0]) +
	( 15'sd 11314) * $signed(input_fmap_205[7:0]) +
	( 15'sd 14742) * $signed(input_fmap_206[7:0]) +
	( 15'sd 12571) * $signed(input_fmap_207[7:0]) +
	( 16'sd 30511) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20516) * $signed(input_fmap_209[7:0]) +
	( 13'sd 3382) * $signed(input_fmap_210[7:0]) +
	( 16'sd 23884) * $signed(input_fmap_211[7:0]) +
	( 16'sd 28037) * $signed(input_fmap_212[7:0]) +
	( 16'sd 32286) * $signed(input_fmap_213[7:0]) +
	( 14'sd 8120) * $signed(input_fmap_214[7:0]) +
	( 14'sd 5020) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4287) * $signed(input_fmap_216[7:0]) +
	( 16'sd 26490) * $signed(input_fmap_217[7:0]) +
	( 16'sd 28998) * $signed(input_fmap_218[7:0]) +
	( 15'sd 10290) * $signed(input_fmap_219[7:0]) +
	( 16'sd 21902) * $signed(input_fmap_220[7:0]) +
	( 15'sd 11772) * $signed(input_fmap_221[7:0]) +
	( 16'sd 30414) * $signed(input_fmap_222[7:0]) +
	( 16'sd 18762) * $signed(input_fmap_223[7:0]) +
	( 16'sd 16726) * $signed(input_fmap_224[7:0]) +
	( 16'sd 26404) * $signed(input_fmap_225[7:0]) +
	( 15'sd 15487) * $signed(input_fmap_226[7:0]) +
	( 16'sd 19328) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26743) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24311) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30314) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24007) * $signed(input_fmap_231[7:0]) +
	( 15'sd 11577) * $signed(input_fmap_232[7:0]) +
	( 14'sd 6120) * $signed(input_fmap_233[7:0]) +
	( 15'sd 10961) * $signed(input_fmap_234[7:0]) +
	( 15'sd 10058) * $signed(input_fmap_235[7:0]) +
	( 15'sd 14119) * $signed(input_fmap_236[7:0]) +
	( 14'sd 7717) * $signed(input_fmap_237[7:0]) +
	( 15'sd 10804) * $signed(input_fmap_238[7:0]) +
	( 16'sd 26784) * $signed(input_fmap_239[7:0]) +
	( 16'sd 19786) * $signed(input_fmap_240[7:0]) +
	( 15'sd 13220) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5246) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6969) * $signed(input_fmap_243[7:0]) +
	( 16'sd 32038) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30718) * $signed(input_fmap_245[7:0]) +
	( 16'sd 25542) * $signed(input_fmap_246[7:0]) +
	( 14'sd 6867) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18295) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2061) * $signed(input_fmap_249[7:0]) +
	( 16'sd 26354) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22947) * $signed(input_fmap_251[7:0]) +
	( 16'sd 29314) * $signed(input_fmap_252[7:0]) +
	( 15'sd 8636) * $signed(input_fmap_253[7:0]) +
	( 16'sd 16734) * $signed(input_fmap_254[7:0]) +
	( 15'sd 9572) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_238;
assign conv_mac_238 = 
	( 15'sd 9505) * $signed(input_fmap_0[7:0]) +
	( 16'sd 31686) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20734) * $signed(input_fmap_2[7:0]) +
	( 16'sd 19640) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24485) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7564) * $signed(input_fmap_5[7:0]) +
	( 16'sd 28785) * $signed(input_fmap_6[7:0]) +
	( 14'sd 6716) * $signed(input_fmap_7[7:0]) +
	( 16'sd 23655) * $signed(input_fmap_8[7:0]) +
	( 16'sd 24007) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32576) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12939) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8666) * $signed(input_fmap_12[7:0]) +
	( 15'sd 8559) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9525) * $signed(input_fmap_14[7:0]) +
	( 16'sd 25125) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12603) * $signed(input_fmap_16[7:0]) +
	( 16'sd 18482) * $signed(input_fmap_17[7:0]) +
	( 16'sd 30697) * $signed(input_fmap_18[7:0]) +
	( 16'sd 26696) * $signed(input_fmap_19[7:0]) +
	( 16'sd 23558) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1262) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9983) * $signed(input_fmap_22[7:0]) +
	( 16'sd 32696) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1426) * $signed(input_fmap_24[7:0]) +
	( 15'sd 8456) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16026) * $signed(input_fmap_26[7:0]) +
	( 16'sd 26505) * $signed(input_fmap_27[7:0]) +
	( 10'sd 458) * $signed(input_fmap_28[7:0]) +
	( 15'sd 9628) * $signed(input_fmap_29[7:0]) +
	( 16'sd 29786) * $signed(input_fmap_30[7:0]) +
	( 16'sd 22020) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28118) * $signed(input_fmap_32[7:0]) +
	( 14'sd 8172) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10202) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15883) * $signed(input_fmap_35[7:0]) +
	( 11'sd 972) * $signed(input_fmap_36[7:0]) +
	( 12'sd 1775) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30232) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17112) * $signed(input_fmap_39[7:0]) +
	( 16'sd 27401) * $signed(input_fmap_40[7:0]) +
	( 16'sd 20291) * $signed(input_fmap_41[7:0]) +
	( 15'sd 11667) * $signed(input_fmap_42[7:0]) +
	( 16'sd 32267) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17342) * $signed(input_fmap_44[7:0]) +
	( 15'sd 13381) * $signed(input_fmap_45[7:0]) +
	( 15'sd 15671) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8165) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14221) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23192) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32297) * $signed(input_fmap_50[7:0]) +
	( 12'sd 1171) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9530) * $signed(input_fmap_52[7:0]) +
	( 16'sd 18862) * $signed(input_fmap_53[7:0]) +
	( 16'sd 22757) * $signed(input_fmap_54[7:0]) +
	( 16'sd 22569) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18878) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10916) * $signed(input_fmap_57[7:0]) +
	( 14'sd 7677) * $signed(input_fmap_58[7:0]) +
	( 16'sd 18477) * $signed(input_fmap_59[7:0]) +
	( 16'sd 22568) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11892) * $signed(input_fmap_61[7:0]) +
	( 14'sd 4944) * $signed(input_fmap_62[7:0]) +
	( 13'sd 2086) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21209) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30430) * $signed(input_fmap_65[7:0]) +
	( 14'sd 6473) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10775) * $signed(input_fmap_67[7:0]) +
	( 13'sd 2122) * $signed(input_fmap_68[7:0]) +
	( 16'sd 25370) * $signed(input_fmap_69[7:0]) +
	( 14'sd 4099) * $signed(input_fmap_70[7:0]) +
	( 13'sd 4054) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23120) * $signed(input_fmap_72[7:0]) +
	( 16'sd 28522) * $signed(input_fmap_73[7:0]) +
	( 16'sd 29645) * $signed(input_fmap_74[7:0]) +
	( 13'sd 3582) * $signed(input_fmap_75[7:0]) +
	( 15'sd 11156) * $signed(input_fmap_76[7:0]) +
	( 16'sd 19102) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24847) * $signed(input_fmap_78[7:0]) +
	( 9'sd 133) * $signed(input_fmap_79[7:0]) +
	( 12'sd 1174) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22543) * $signed(input_fmap_81[7:0]) +
	( 13'sd 3412) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19793) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3716) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_85[7:0]) +
	( 14'sd 4314) * $signed(input_fmap_86[7:0]) +
	( 13'sd 3069) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25255) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19429) * $signed(input_fmap_89[7:0]) +
	( 15'sd 8435) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24706) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9989) * $signed(input_fmap_92[7:0]) +
	( 16'sd 25986) * $signed(input_fmap_93[7:0]) +
	( 16'sd 20800) * $signed(input_fmap_94[7:0]) +
	( 14'sd 8121) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6190) * $signed(input_fmap_96[7:0]) +
	( 16'sd 18443) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2335) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27810) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13088) * $signed(input_fmap_100[7:0]) +
	( 16'sd 21683) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4481) * $signed(input_fmap_102[7:0]) +
	( 16'sd 20898) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12620) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30842) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17268) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7443) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30221) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28894) * $signed(input_fmap_109[7:0]) +
	( 13'sd 3240) * $signed(input_fmap_110[7:0]) +
	( 16'sd 20593) * $signed(input_fmap_111[7:0]) +
	( 16'sd 21859) * $signed(input_fmap_112[7:0]) +
	( 16'sd 30828) * $signed(input_fmap_113[7:0]) +
	( 15'sd 15346) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1061) * $signed(input_fmap_115[7:0]) +
	( 16'sd 31382) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17255) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7157) * $signed(input_fmap_118[7:0]) +
	( 16'sd 30733) * $signed(input_fmap_119[7:0]) +
	( 16'sd 17909) * $signed(input_fmap_120[7:0]) +
	( 12'sd 1136) * $signed(input_fmap_121[7:0]) +
	( 16'sd 21519) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22939) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28410) * $signed(input_fmap_124[7:0]) +
	( 16'sd 32664) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1742) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2200) * $signed(input_fmap_127[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_128[7:0]) +
	( 16'sd 19297) * $signed(input_fmap_129[7:0]) +
	( 14'sd 7997) * $signed(input_fmap_130[7:0]) +
	( 16'sd 30424) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_132[7:0]) +
	( 16'sd 18667) * $signed(input_fmap_133[7:0]) +
	( 11'sd 515) * $signed(input_fmap_134[7:0]) +
	( 16'sd 31095) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30136) * $signed(input_fmap_136[7:0]) +
	( 15'sd 14582) * $signed(input_fmap_137[7:0]) +
	( 16'sd 30689) * $signed(input_fmap_138[7:0]) +
	( 15'sd 15834) * $signed(input_fmap_139[7:0]) +
	( 16'sd 25812) * $signed(input_fmap_140[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_141[7:0]) +
	( 16'sd 21558) * $signed(input_fmap_142[7:0]) +
	( 16'sd 18802) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18348) * $signed(input_fmap_144[7:0]) +
	( 16'sd 32538) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21199) * $signed(input_fmap_146[7:0]) +
	( 16'sd 23256) * $signed(input_fmap_147[7:0]) +
	( 14'sd 7681) * $signed(input_fmap_148[7:0]) +
	( 16'sd 26386) * $signed(input_fmap_149[7:0]) +
	( 14'sd 6308) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19850) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24438) * $signed(input_fmap_152[7:0]) +
	( 16'sd 22001) * $signed(input_fmap_153[7:0]) +
	( 16'sd 21826) * $signed(input_fmap_154[7:0]) +
	( 16'sd 19484) * $signed(input_fmap_155[7:0]) +
	( 15'sd 8342) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30821) * $signed(input_fmap_157[7:0]) +
	( 14'sd 5545) * $signed(input_fmap_158[7:0]) +
	( 15'sd 11985) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27900) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23416) * $signed(input_fmap_161[7:0]) +
	( 15'sd 9818) * $signed(input_fmap_162[7:0]) +
	( 16'sd 18661) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6030) * $signed(input_fmap_164[7:0]) +
	( 13'sd 3667) * $signed(input_fmap_165[7:0]) +
	( 16'sd 17218) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13762) * $signed(input_fmap_167[7:0]) +
	( 16'sd 20051) * $signed(input_fmap_168[7:0]) +
	( 16'sd 27055) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5082) * $signed(input_fmap_170[7:0]) +
	( 16'sd 32057) * $signed(input_fmap_171[7:0]) +
	( 15'sd 13897) * $signed(input_fmap_172[7:0]) +
	( 15'sd 12565) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7812) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4436) * $signed(input_fmap_175[7:0]) +
	( 15'sd 9755) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2985) * $signed(input_fmap_177[7:0]) +
	( 15'sd 12577) * $signed(input_fmap_178[7:0]) +
	( 15'sd 16177) * $signed(input_fmap_179[7:0]) +
	( 12'sd 1980) * $signed(input_fmap_180[7:0]) +
	( 14'sd 6221) * $signed(input_fmap_181[7:0]) +
	( 16'sd 16468) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2602) * $signed(input_fmap_183[7:0]) +
	( 13'sd 3088) * $signed(input_fmap_184[7:0]) +
	( 16'sd 21061) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6137) * $signed(input_fmap_186[7:0]) +
	( 11'sd 768) * $signed(input_fmap_187[7:0]) +
	( 15'sd 15258) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7034) * $signed(input_fmap_189[7:0]) +
	( 16'sd 30493) * $signed(input_fmap_190[7:0]) +
	( 16'sd 24333) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31660) * $signed(input_fmap_192[7:0]) +
	( 16'sd 17588) * $signed(input_fmap_193[7:0]) +
	( 16'sd 18301) * $signed(input_fmap_194[7:0]) +
	( 11'sd 755) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7621) * $signed(input_fmap_196[7:0]) +
	( 14'sd 5555) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27422) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12667) * $signed(input_fmap_199[7:0]) +
	( 12'sd 1157) * $signed(input_fmap_200[7:0]) +
	( 15'sd 12605) * $signed(input_fmap_201[7:0]) +
	( 16'sd 26779) * $signed(input_fmap_202[7:0]) +
	( 15'sd 15454) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32222) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5067) * $signed(input_fmap_205[7:0]) +
	( 11'sd 556) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28745) * $signed(input_fmap_207[7:0]) +
	( 15'sd 10746) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11815) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18376) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6378) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12033) * $signed(input_fmap_212[7:0]) +
	( 16'sd 24476) * $signed(input_fmap_213[7:0]) +
	( 16'sd 25697) * $signed(input_fmap_214[7:0]) +
	( 16'sd 20368) * $signed(input_fmap_215[7:0]) +
	( 16'sd 28933) * $signed(input_fmap_216[7:0]) +
	( 15'sd 13004) * $signed(input_fmap_217[7:0]) +
	( 14'sd 5420) * $signed(input_fmap_218[7:0]) +
	( 16'sd 30700) * $signed(input_fmap_219[7:0]) +
	( 16'sd 31758) * $signed(input_fmap_220[7:0]) +
	( 15'sd 15928) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5752) * $signed(input_fmap_222[7:0]) +
	( 16'sd 24585) * $signed(input_fmap_223[7:0]) +
	( 16'sd 17454) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20344) * $signed(input_fmap_225[7:0]) +
	( 12'sd 1487) * $signed(input_fmap_226[7:0]) +
	( 15'sd 12861) * $signed(input_fmap_227[7:0]) +
	( 16'sd 27252) * $signed(input_fmap_228[7:0]) +
	( 16'sd 17946) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29950) * $signed(input_fmap_230[7:0]) +
	( 14'sd 6809) * $signed(input_fmap_231[7:0]) +
	( 15'sd 11196) * $signed(input_fmap_232[7:0]) +
	( 16'sd 32468) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14279) * $signed(input_fmap_234[7:0]) +
	( 16'sd 28975) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30333) * $signed(input_fmap_236[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_237[7:0]) +
	( 16'sd 28055) * $signed(input_fmap_238[7:0]) +
	( 15'sd 10800) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9345) * $signed(input_fmap_240[7:0]) +
	( 16'sd 32386) * $signed(input_fmap_241[7:0]) +
	( 16'sd 25455) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7480) * $signed(input_fmap_243[7:0]) +
	( 15'sd 11698) * $signed(input_fmap_244[7:0]) +
	( 15'sd 15211) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22474) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30129) * $signed(input_fmap_247[7:0]) +
	( 16'sd 20067) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21710) * $signed(input_fmap_249[7:0]) +
	( 15'sd 15815) * $signed(input_fmap_250[7:0]) +
	( 16'sd 26602) * $signed(input_fmap_251[7:0]) +
	( 15'sd 10983) * $signed(input_fmap_252[7:0]) +
	( 15'sd 12193) * $signed(input_fmap_253[7:0]) +
	( 15'sd 12946) * $signed(input_fmap_254[7:0]) +
	( 16'sd 21674) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_239;
assign conv_mac_239 = 
	( 15'sd 15307) * $signed(input_fmap_0[7:0]) +
	( 14'sd 7019) * $signed(input_fmap_1[7:0]) +
	( 16'sd 17740) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9969) * $signed(input_fmap_3[7:0]) +
	( 16'sd 28984) * $signed(input_fmap_4[7:0]) +
	( 14'sd 4733) * $signed(input_fmap_5[7:0]) +
	( 16'sd 21732) * $signed(input_fmap_6[7:0]) +
	( 15'sd 9051) * $signed(input_fmap_7[7:0]) +
	( 14'sd 4337) * $signed(input_fmap_8[7:0]) +
	( 15'sd 9476) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26647) * $signed(input_fmap_10[7:0]) +
	( 15'sd 9309) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25627) * $signed(input_fmap_12[7:0]) +
	( 15'sd 14569) * $signed(input_fmap_13[7:0]) +
	( 15'sd 14987) * $signed(input_fmap_14[7:0]) +
	( 15'sd 15818) * $signed(input_fmap_15[7:0]) +
	( 16'sd 32469) * $signed(input_fmap_16[7:0]) +
	( 16'sd 17985) * $signed(input_fmap_17[7:0]) +
	( 12'sd 1668) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18320) * $signed(input_fmap_19[7:0]) +
	( 16'sd 29014) * $signed(input_fmap_20[7:0]) +
	( 16'sd 21013) * $signed(input_fmap_21[7:0]) +
	( 16'sd 29814) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18626) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20418) * $signed(input_fmap_24[7:0]) +
	( 13'sd 3286) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28938) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20791) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16630) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15863) * $signed(input_fmap_29[7:0]) +
	( 16'sd 18071) * $signed(input_fmap_30[7:0]) +
	( 16'sd 17257) * $signed(input_fmap_31[7:0]) +
	( 11'sd 807) * $signed(input_fmap_32[7:0]) +
	( 13'sd 3819) * $signed(input_fmap_33[7:0]) +
	( 15'sd 10283) * $signed(input_fmap_34[7:0]) +
	( 15'sd 10048) * $signed(input_fmap_35[7:0]) +
	( 14'sd 6607) * $signed(input_fmap_36[7:0]) +
	( 15'sd 8819) * $signed(input_fmap_37[7:0]) +
	( 15'sd 9301) * $signed(input_fmap_38[7:0]) +
	( 16'sd 29863) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20630) * $signed(input_fmap_40[7:0]) +
	( 8'sd 123) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6119) * $signed(input_fmap_42[7:0]) +
	( 12'sd 1891) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26298) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27638) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14068) * $signed(input_fmap_46[7:0]) +
	( 16'sd 20904) * $signed(input_fmap_47[7:0]) +
	( 14'sd 6844) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8399) * $signed(input_fmap_49[7:0]) +
	( 16'sd 23774) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27169) * $signed(input_fmap_51[7:0]) +
	( 14'sd 7353) * $signed(input_fmap_52[7:0]) +
	( 13'sd 3674) * $signed(input_fmap_53[7:0]) +
	( 16'sd 30518) * $signed(input_fmap_54[7:0]) +
	( 15'sd 8229) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26798) * $signed(input_fmap_56[7:0]) +
	( 14'sd 5767) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3123) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19482) * $signed(input_fmap_59[7:0]) +
	( 16'sd 26313) * $signed(input_fmap_60[7:0]) +
	( 16'sd 23005) * $signed(input_fmap_61[7:0]) +
	( 15'sd 14541) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13332) * $signed(input_fmap_63[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_64[7:0]) +
	( 15'sd 15190) * $signed(input_fmap_65[7:0]) +
	( 16'sd 20897) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13311) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14347) * $signed(input_fmap_68[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20376) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27336) * $signed(input_fmap_71[7:0]) +
	( 9'sd 233) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29235) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21799) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6909) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30819) * $signed(input_fmap_76[7:0]) +
	( 16'sd 21162) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24442) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3774) * $signed(input_fmap_79[7:0]) +
	( 16'sd 24035) * $signed(input_fmap_80[7:0]) +
	( 15'sd 14714) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9909) * $signed(input_fmap_82[7:0]) +
	( 13'sd 2796) * $signed(input_fmap_83[7:0]) +
	( 15'sd 9796) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19476) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8967) * $signed(input_fmap_86[7:0]) +
	( 16'sd 21375) * $signed(input_fmap_87[7:0]) +
	( 16'sd 25989) * $signed(input_fmap_88[7:0]) +
	( 10'sd 345) * $signed(input_fmap_89[7:0]) +
	( 14'sd 4796) * $signed(input_fmap_90[7:0]) +
	( 16'sd 20495) * $signed(input_fmap_91[7:0]) +
	( 16'sd 19547) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22290) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13578) * $signed(input_fmap_94[7:0]) +
	( 12'sd 1275) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8393) * $signed(input_fmap_96[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22542) * $signed(input_fmap_98[7:0]) +
	( 15'sd 8520) * $signed(input_fmap_99[7:0]) +
	( 11'sd 996) * $signed(input_fmap_100[7:0]) +
	( 15'sd 16188) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28701) * $signed(input_fmap_102[7:0]) +
	( 16'sd 17999) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30463) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28272) * $signed(input_fmap_105[7:0]) +
	( 15'sd 8411) * $signed(input_fmap_106[7:0]) +
	( 14'sd 6246) * $signed(input_fmap_107[7:0]) +
	( 16'sd 25178) * $signed(input_fmap_108[7:0]) +
	( 16'sd 16762) * $signed(input_fmap_109[7:0]) +
	( 16'sd 24501) * $signed(input_fmap_110[7:0]) +
	( 14'sd 5480) * $signed(input_fmap_111[7:0]) +
	( 15'sd 16298) * $signed(input_fmap_112[7:0]) +
	( 16'sd 26701) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32451) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5955) * $signed(input_fmap_115[7:0]) +
	( 16'sd 30763) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27597) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4428) * $signed(input_fmap_118[7:0]) +
	( 15'sd 13795) * $signed(input_fmap_119[7:0]) +
	( 13'sd 2913) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7216) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1540) * $signed(input_fmap_122[7:0]) +
	( 14'sd 5623) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23145) * $signed(input_fmap_124[7:0]) +
	( 11'sd 941) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29240) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26276) * $signed(input_fmap_127[7:0]) +
	( 15'sd 11733) * $signed(input_fmap_128[7:0]) +
	( 15'sd 14205) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25167) * $signed(input_fmap_130[7:0]) +
	( 16'sd 24059) * $signed(input_fmap_131[7:0]) +
	( 16'sd 17796) * $signed(input_fmap_132[7:0]) +
	( 16'sd 19809) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32024) * $signed(input_fmap_134[7:0]) +
	( 15'sd 14217) * $signed(input_fmap_135[7:0]) +
	( 14'sd 8146) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27355) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11784) * $signed(input_fmap_138[7:0]) +
	( 16'sd 26110) * $signed(input_fmap_139[7:0]) +
	( 15'sd 13120) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10912) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6881) * $signed(input_fmap_142[7:0]) +
	( 15'sd 15930) * $signed(input_fmap_143[7:0]) +
	( 16'sd 32533) * $signed(input_fmap_144[7:0]) +
	( 16'sd 29103) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21996) * $signed(input_fmap_146[7:0]) +
	( 16'sd 32674) * $signed(input_fmap_147[7:0]) +
	( 16'sd 17651) * $signed(input_fmap_148[7:0]) +
	( 16'sd 22691) * $signed(input_fmap_149[7:0]) +
	( 16'sd 21095) * $signed(input_fmap_150[7:0]) +
	( 16'sd 21376) * $signed(input_fmap_151[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_152[7:0]) +
	( 16'sd 29291) * $signed(input_fmap_153[7:0]) +
	( 9'sd 183) * $signed(input_fmap_154[7:0]) +
	( 16'sd 21031) * $signed(input_fmap_155[7:0]) +
	( 15'sd 13665) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13840) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4495) * $signed(input_fmap_158[7:0]) +
	( 15'sd 9538) * $signed(input_fmap_159[7:0]) +
	( 16'sd 31724) * $signed(input_fmap_160[7:0]) +
	( 9'sd 168) * $signed(input_fmap_161[7:0]) +
	( 13'sd 3129) * $signed(input_fmap_162[7:0]) +
	( 16'sd 20210) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24010) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10911) * $signed(input_fmap_165[7:0]) +
	( 15'sd 14585) * $signed(input_fmap_166[7:0]) +
	( 16'sd 27380) * $signed(input_fmap_167[7:0]) +
	( 13'sd 2711) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11192) * $signed(input_fmap_169[7:0]) +
	( 15'sd 12876) * $signed(input_fmap_170[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_171[7:0]) +
	( 16'sd 31122) * $signed(input_fmap_172[7:0]) +
	( 14'sd 4575) * $signed(input_fmap_173[7:0]) +
	( 10'sd 409) * $signed(input_fmap_174[7:0]) +
	( 14'sd 5359) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7941) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30904) * $signed(input_fmap_177[7:0]) +
	( 16'sd 31778) * $signed(input_fmap_178[7:0]) +
	( 13'sd 2803) * $signed(input_fmap_179[7:0]) +
	( 14'sd 8047) * $signed(input_fmap_180[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12193) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2516) * $signed(input_fmap_183[7:0]) +
	( 16'sd 22595) * $signed(input_fmap_184[7:0]) +
	( 16'sd 32741) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12475) * $signed(input_fmap_186[7:0]) +
	( 15'sd 15964) * $signed(input_fmap_187[7:0]) +
	( 14'sd 7457) * $signed(input_fmap_188[7:0]) +
	( 16'sd 26483) * $signed(input_fmap_189[7:0]) +
	( 16'sd 26188) * $signed(input_fmap_190[7:0]) +
	( 15'sd 14954) * $signed(input_fmap_191[7:0]) +
	( 14'sd 5518) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22810) * $signed(input_fmap_193[7:0]) +
	( 16'sd 24575) * $signed(input_fmap_194[7:0]) +
	( 16'sd 28582) * $signed(input_fmap_195[7:0]) +
	( 14'sd 4588) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_197[7:0]) +
	( 16'sd 21891) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10139) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13414) * $signed(input_fmap_200[7:0]) +
	( 16'sd 17501) * $signed(input_fmap_201[7:0]) +
	( 14'sd 6823) * $signed(input_fmap_202[7:0]) +
	( 14'sd 5678) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6086) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15514) * $signed(input_fmap_205[7:0]) +
	( 15'sd 14078) * $signed(input_fmap_206[7:0]) +
	( 16'sd 20405) * $signed(input_fmap_207[7:0]) +
	( 14'sd 6104) * $signed(input_fmap_208[7:0]) +
	( 16'sd 16768) * $signed(input_fmap_209[7:0]) +
	( 15'sd 14945) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17202) * $signed(input_fmap_211[7:0]) +
	( 16'sd 29984) * $signed(input_fmap_212[7:0]) +
	( 12'sd 1344) * $signed(input_fmap_213[7:0]) +
	( 15'sd 10676) * $signed(input_fmap_214[7:0]) +
	( 13'sd 2372) * $signed(input_fmap_215[7:0]) +
	( 14'sd 5113) * $signed(input_fmap_216[7:0]) +
	( 16'sd 18364) * $signed(input_fmap_217[7:0]) +
	( 15'sd 15540) * $signed(input_fmap_218[7:0]) +
	( 16'sd 26061) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24336) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28315) * $signed(input_fmap_221[7:0]) +
	( 15'sd 12292) * $signed(input_fmap_222[7:0]) +
	( 16'sd 31228) * $signed(input_fmap_223[7:0]) +
	( 14'sd 6094) * $signed(input_fmap_224[7:0]) +
	( 15'sd 11848) * $signed(input_fmap_225[7:0]) +
	( 15'sd 15287) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2925) * $signed(input_fmap_227[7:0]) +
	( 14'sd 7487) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3916) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28583) * $signed(input_fmap_230[7:0]) +
	( 16'sd 18106) * $signed(input_fmap_231[7:0]) +
	( 16'sd 26348) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14735) * $signed(input_fmap_233[7:0]) +
	( 15'sd 8302) * $signed(input_fmap_234[7:0]) +
	( 16'sd 20006) * $signed(input_fmap_235[7:0]) +
	( 16'sd 31517) * $signed(input_fmap_236[7:0]) +
	( 16'sd 27423) * $signed(input_fmap_237[7:0]) +
	( 14'sd 5312) * $signed(input_fmap_238[7:0]) +
	( 15'sd 13123) * $signed(input_fmap_239[7:0]) +
	( 15'sd 11076) * $signed(input_fmap_240[7:0]) +
	( 14'sd 4482) * $signed(input_fmap_241[7:0]) +
	( 14'sd 6518) * $signed(input_fmap_242[7:0]) +
	( 12'sd 1496) * $signed(input_fmap_243[7:0]) +
	( 16'sd 27218) * $signed(input_fmap_244[7:0]) +
	( 15'sd 10470) * $signed(input_fmap_245[7:0]) +
	( 16'sd 25343) * $signed(input_fmap_246[7:0]) +
	( 8'sd 80) * $signed(input_fmap_247[7:0]) +
	( 10'sd 376) * $signed(input_fmap_248[7:0]) +
	( 15'sd 13595) * $signed(input_fmap_249[7:0]) +
	( 16'sd 32141) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4110) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4139) * $signed(input_fmap_252[7:0]) +
	( 16'sd 20998) * $signed(input_fmap_253[7:0]) +
	( 14'sd 7211) * $signed(input_fmap_254[7:0]) +
	( 16'sd 25381) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_240;
assign conv_mac_240 = 
	( 16'sd 30312) * $signed(input_fmap_0[7:0]) +
	( 16'sd 20869) * $signed(input_fmap_1[7:0]) +
	( 11'sd 840) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9784) * $signed(input_fmap_3[7:0]) +
	( 16'sd 20433) * $signed(input_fmap_4[7:0]) +
	( 16'sd 30781) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25223) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29033) * $signed(input_fmap_7[7:0]) +
	( 16'sd 24336) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30765) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5336) * $signed(input_fmap_10[7:0]) +
	( 15'sd 12555) * $signed(input_fmap_11[7:0]) +
	( 16'sd 24010) * $signed(input_fmap_12[7:0]) +
	( 16'sd 26238) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9446) * $signed(input_fmap_14[7:0]) +
	( 15'sd 9637) * $signed(input_fmap_15[7:0]) +
	( 11'sd 820) * $signed(input_fmap_16[7:0]) +
	( 16'sd 22894) * $signed(input_fmap_17[7:0]) +
	( 13'sd 3652) * $signed(input_fmap_18[7:0]) +
	( 16'sd 18596) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11086) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3879) * $signed(input_fmap_21[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_22[7:0]) +
	( 14'sd 8075) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1050) * $signed(input_fmap_24[7:0]) +
	( 15'sd 13036) * $signed(input_fmap_25[7:0]) +
	( 15'sd 8508) * $signed(input_fmap_26[7:0]) +
	( 16'sd 20163) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10725) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3192) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10597) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4248) * $signed(input_fmap_31[7:0]) +
	( 16'sd 28505) * $signed(input_fmap_32[7:0]) +
	( 16'sd 19552) * $signed(input_fmap_33[7:0]) +
	( 16'sd 18222) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26938) * $signed(input_fmap_35[7:0]) +
	( 16'sd 19125) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6169) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17900) * $signed(input_fmap_39[7:0]) +
	( 14'sd 6969) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11003) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6776) * $signed(input_fmap_42[7:0]) +
	( 16'sd 18019) * $signed(input_fmap_43[7:0]) +
	( 16'sd 26334) * $signed(input_fmap_44[7:0]) +
	( 12'sd 1382) * $signed(input_fmap_45[7:0]) +
	( 13'sd 3233) * $signed(input_fmap_46[7:0]) +
	( 16'sd 25794) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24589) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26157) * $signed(input_fmap_50[7:0]) +
	( 16'sd 27256) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16522) * $signed(input_fmap_52[7:0]) +
	( 16'sd 22097) * $signed(input_fmap_53[7:0]) +
	( 16'sd 21890) * $signed(input_fmap_54[7:0]) +
	( 15'sd 10763) * $signed(input_fmap_55[7:0]) +
	( 16'sd 29749) * $signed(input_fmap_56[7:0]) +
	( 16'sd 20309) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17848) * $signed(input_fmap_58[7:0]) +
	( 14'sd 7585) * $signed(input_fmap_59[7:0]) +
	( 8'sd 85) * $signed(input_fmap_60[7:0]) +
	( 16'sd 24880) * $signed(input_fmap_61[7:0]) +
	( 16'sd 29286) * $signed(input_fmap_62[7:0]) +
	( 16'sd 32288) * $signed(input_fmap_63[7:0]) +
	( 15'sd 13741) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30301) * $signed(input_fmap_65[7:0]) +
	( 15'sd 16342) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7251) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5003) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14368) * $signed(input_fmap_69[7:0]) +
	( 16'sd 22082) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2343) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20198) * $signed(input_fmap_72[7:0]) +
	( 14'sd 6713) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9165) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24623) * $signed(input_fmap_75[7:0]) +
	( 14'sd 8142) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27165) * $signed(input_fmap_77[7:0]) +
	( 15'sd 13779) * $signed(input_fmap_78[7:0]) +
	( 16'sd 25484) * $signed(input_fmap_79[7:0]) +
	( 16'sd 17155) * $signed(input_fmap_80[7:0]) +
	( 16'sd 22490) * $signed(input_fmap_81[7:0]) +
	( 14'sd 4199) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5025) * $signed(input_fmap_83[7:0]) +
	( 15'sd 16135) * $signed(input_fmap_84[7:0]) +
	( 16'sd 31819) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15163) * $signed(input_fmap_86[7:0]) +
	( 14'sd 5092) * $signed(input_fmap_87[7:0]) +
	( 16'sd 19915) * $signed(input_fmap_88[7:0]) +
	( 15'sd 12419) * $signed(input_fmap_89[7:0]) +
	( 16'sd 26683) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11017) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31422) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24747) * $signed(input_fmap_93[7:0]) +
	( 13'sd 3408) * $signed(input_fmap_94[7:0]) +
	( 15'sd 14805) * $signed(input_fmap_95[7:0]) +
	( 14'sd 4661) * $signed(input_fmap_96[7:0]) +
	( 14'sd 4736) * $signed(input_fmap_97[7:0]) +
	( 15'sd 14915) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18546) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30716) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31898) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29067) * $signed(input_fmap_102[7:0]) +
	( 13'sd 3354) * $signed(input_fmap_103[7:0]) +
	( 15'sd 13367) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17998) * $signed(input_fmap_105[7:0]) +
	( 16'sd 21656) * $signed(input_fmap_106[7:0]) +
	( 16'sd 19829) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28971) * $signed(input_fmap_108[7:0]) +
	( 16'sd 32424) * $signed(input_fmap_109[7:0]) +
	( 16'sd 29381) * $signed(input_fmap_110[7:0]) +
	( 16'sd 30955) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4510) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5762) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16142) * $signed(input_fmap_114[7:0]) +
	( 16'sd 20280) * $signed(input_fmap_115[7:0]) +
	( 16'sd 20928) * $signed(input_fmap_116[7:0]) +
	( 16'sd 25588) * $signed(input_fmap_117[7:0]) +
	( 14'sd 8082) * $signed(input_fmap_118[7:0]) +
	( 10'sd 323) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11297) * $signed(input_fmap_120[7:0]) +
	( 16'sd 25096) * $signed(input_fmap_121[7:0]) +
	( 16'sd 26075) * $signed(input_fmap_122[7:0]) +
	( 15'sd 13525) * $signed(input_fmap_123[7:0]) +
	( 15'sd 10727) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27277) * $signed(input_fmap_125[7:0]) +
	( 14'sd 6040) * $signed(input_fmap_126[7:0]) +
	( 14'sd 5227) * $signed(input_fmap_127[7:0]) +
	( 14'sd 4289) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7345) * $signed(input_fmap_129[7:0]) +
	( 15'sd 15509) * $signed(input_fmap_130[7:0]) +
	( 16'sd 29602) * $signed(input_fmap_131[7:0]) +
	( 16'sd 24061) * $signed(input_fmap_132[7:0]) +
	( 16'sd 18512) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1890) * $signed(input_fmap_134[7:0]) +
	( 15'sd 11561) * $signed(input_fmap_135[7:0]) +
	( 16'sd 30030) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6314) * $signed(input_fmap_137[7:0]) +
	( 15'sd 13225) * $signed(input_fmap_138[7:0]) +
	( 15'sd 16041) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9405) * $signed(input_fmap_140[7:0]) +
	( 14'sd 7659) * $signed(input_fmap_141[7:0]) +
	( 16'sd 24702) * $signed(input_fmap_142[7:0]) +
	( 16'sd 25610) * $signed(input_fmap_143[7:0]) +
	( 13'sd 2258) * $signed(input_fmap_144[7:0]) +
	( 13'sd 3645) * $signed(input_fmap_145[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_146[7:0]) +
	( 7'sd 41) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11671) * $signed(input_fmap_148[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_149[7:0]) +
	( 16'sd 16765) * $signed(input_fmap_150[7:0]) +
	( 14'sd 5638) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14996) * $signed(input_fmap_152[7:0]) +
	( 16'sd 16742) * $signed(input_fmap_153[7:0]) +
	( 16'sd 23445) * $signed(input_fmap_154[7:0]) +
	( 16'sd 20906) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20439) * $signed(input_fmap_156[7:0]) +
	( 14'sd 4290) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4228) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6792) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21403) * $signed(input_fmap_160[7:0]) +
	( 15'sd 11318) * $signed(input_fmap_161[7:0]) +
	( 16'sd 22183) * $signed(input_fmap_162[7:0]) +
	( 13'sd 4092) * $signed(input_fmap_163[7:0]) +
	( 16'sd 23663) * $signed(input_fmap_164[7:0]) +
	( 11'sd 972) * $signed(input_fmap_165[7:0]) +
	( 15'sd 11405) * $signed(input_fmap_166[7:0]) +
	( 14'sd 6660) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26053) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26077) * $signed(input_fmap_169[7:0]) +
	( 15'sd 10566) * $signed(input_fmap_170[7:0]) +
	( 16'sd 21785) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22777) * $signed(input_fmap_172[7:0]) +
	( 14'sd 6171) * $signed(input_fmap_173[7:0]) +
	( 15'sd 11056) * $signed(input_fmap_174[7:0]) +
	( 15'sd 9706) * $signed(input_fmap_175[7:0]) +
	( 16'sd 17543) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30616) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32043) * $signed(input_fmap_178[7:0]) +
	( 15'sd 14754) * $signed(input_fmap_179[7:0]) +
	( 16'sd 18281) * $signed(input_fmap_180[7:0]) +
	( 16'sd 17027) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30706) * $signed(input_fmap_182[7:0]) +
	( 16'sd 29981) * $signed(input_fmap_183[7:0]) +
	( 16'sd 17185) * $signed(input_fmap_184[7:0]) +
	( 16'sd 32074) * $signed(input_fmap_185[7:0]) +
	( 16'sd 25386) * $signed(input_fmap_186[7:0]) +
	( 16'sd 21658) * $signed(input_fmap_187[7:0]) +
	( 15'sd 9596) * $signed(input_fmap_188[7:0]) +
	( 14'sd 4766) * $signed(input_fmap_189[7:0]) +
	( 16'sd 26747) * $signed(input_fmap_190[7:0]) +
	( 15'sd 11990) * $signed(input_fmap_191[7:0]) +
	( 14'sd 6729) * $signed(input_fmap_192[7:0]) +
	( 16'sd 17500) * $signed(input_fmap_193[7:0]) +
	( 10'sd 294) * $signed(input_fmap_194[7:0]) +
	( 12'sd 1659) * $signed(input_fmap_195[7:0]) +
	( 13'sd 3357) * $signed(input_fmap_196[7:0]) +
	( 16'sd 24609) * $signed(input_fmap_197[7:0]) +
	( 14'sd 7601) * $signed(input_fmap_198[7:0]) +
	( 13'sd 3174) * $signed(input_fmap_199[7:0]) +
	( 15'sd 11744) * $signed(input_fmap_200[7:0]) +
	( 16'sd 28692) * $signed(input_fmap_201[7:0]) +
	( 16'sd 30721) * $signed(input_fmap_202[7:0]) +
	( 14'sd 7165) * $signed(input_fmap_203[7:0]) +
	( 16'sd 31045) * $signed(input_fmap_204[7:0]) +
	( 15'sd 13702) * $signed(input_fmap_205[7:0]) +
	( 16'sd 16866) * $signed(input_fmap_206[7:0]) +
	( 16'sd 18743) * $signed(input_fmap_207[7:0]) +
	( 16'sd 17980) * $signed(input_fmap_208[7:0]) +
	( 16'sd 25138) * $signed(input_fmap_209[7:0]) +
	( 16'sd 18637) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28888) * $signed(input_fmap_211[7:0]) +
	( 15'sd 14710) * $signed(input_fmap_212[7:0]) +
	( 16'sd 29992) * $signed(input_fmap_213[7:0]) +
	( 16'sd 23338) * $signed(input_fmap_214[7:0]) +
	( 16'sd 24978) * $signed(input_fmap_215[7:0]) +
	( 14'sd 6872) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9168) * $signed(input_fmap_217[7:0]) +
	( 16'sd 16613) * $signed(input_fmap_218[7:0]) +
	( 15'sd 12386) * $signed(input_fmap_219[7:0]) +
	( 15'sd 9999) * $signed(input_fmap_220[7:0]) +
	( 15'sd 12989) * $signed(input_fmap_221[7:0]) +
	( 16'sd 20954) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2206) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25185) * $signed(input_fmap_224[7:0]) +
	( 15'sd 9090) * $signed(input_fmap_225[7:0]) +
	( 12'sd 1325) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5881) * $signed(input_fmap_227[7:0]) +
	( 15'sd 12981) * $signed(input_fmap_228[7:0]) +
	( 15'sd 8967) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18022) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14215) * $signed(input_fmap_231[7:0]) +
	( 16'sd 26030) * $signed(input_fmap_232[7:0]) +
	( 15'sd 10541) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4605) * $signed(input_fmap_234[7:0]) +
	( 11'sd 960) * $signed(input_fmap_235[7:0]) +
	( 16'sd 27073) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28124) * $signed(input_fmap_237[7:0]) +
	( 15'sd 16032) * $signed(input_fmap_238[7:0]) +
	( 14'sd 5178) * $signed(input_fmap_239[7:0]) +
	( 16'sd 16713) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18758) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29771) * $signed(input_fmap_242[7:0]) +
	( 16'sd 28295) * $signed(input_fmap_243[7:0]) +
	( 15'sd 14064) * $signed(input_fmap_244[7:0]) +
	( 16'sd 25111) * $signed(input_fmap_245[7:0]) +
	( 15'sd 12931) * $signed(input_fmap_246[7:0]) +
	( 16'sd 17129) * $signed(input_fmap_247[7:0]) +
	( 16'sd 30666) * $signed(input_fmap_248[7:0]) +
	( 16'sd 21218) * $signed(input_fmap_249[7:0]) +
	( 16'sd 28749) * $signed(input_fmap_250[7:0]) +
	( 15'sd 15705) * $signed(input_fmap_251[7:0]) +
	( 16'sd 30447) * $signed(input_fmap_252[7:0]) +
	( 16'sd 26712) * $signed(input_fmap_253[7:0]) +
	( 16'sd 20413) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26011) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_241;
assign conv_mac_241 = 
	( 11'sd 668) * $signed(input_fmap_0[7:0]) +
	( 15'sd 16379) * $signed(input_fmap_1[7:0]) +
	( 16'sd 28142) * $signed(input_fmap_2[7:0]) +
	( 15'sd 8671) * $signed(input_fmap_3[7:0]) +
	( 15'sd 12891) * $signed(input_fmap_4[7:0]) +
	( 10'sd 501) * $signed(input_fmap_5[7:0]) +
	( 15'sd 12324) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19391) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28161) * $signed(input_fmap_8[7:0]) +
	( 16'sd 25479) * $signed(input_fmap_9[7:0]) +
	( 14'sd 4148) * $signed(input_fmap_10[7:0]) +
	( 16'sd 23162) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1485) * $signed(input_fmap_12[7:0]) +
	( 13'sd 3937) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7323) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28537) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30299) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11696) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15049) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25891) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22848) * $signed(input_fmap_20[7:0]) +
	( 15'sd 10604) * $signed(input_fmap_21[7:0]) +
	( 15'sd 12170) * $signed(input_fmap_22[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_23[7:0]) +
	( 16'sd 32410) * $signed(input_fmap_24[7:0]) +
	( 14'sd 8051) * $signed(input_fmap_25[7:0]) +
	( 16'sd 27665) * $signed(input_fmap_26[7:0]) +
	( 16'sd 18606) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10883) * $signed(input_fmap_28[7:0]) +
	( 16'sd 26759) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10969) * $signed(input_fmap_30[7:0]) +
	( 15'sd 11246) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18334) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8379) * $signed(input_fmap_33[7:0]) +
	( 16'sd 19282) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21293) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22366) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26978) * $signed(input_fmap_37[7:0]) +
	( 15'sd 13887) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30233) * $signed(input_fmap_39[7:0]) +
	( 16'sd 21361) * $signed(input_fmap_40[7:0]) +
	( 16'sd 24529) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3365) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26478) * $signed(input_fmap_43[7:0]) +
	( 15'sd 11484) * $signed(input_fmap_44[7:0]) +
	( 16'sd 27814) * $signed(input_fmap_45[7:0]) +
	( 16'sd 19626) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17753) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24175) * $signed(input_fmap_48[7:0]) +
	( 14'sd 5997) * $signed(input_fmap_49[7:0]) +
	( 16'sd 27424) * $signed(input_fmap_50[7:0]) +
	( 16'sd 25299) * $signed(input_fmap_51[7:0]) +
	( 16'sd 28873) * $signed(input_fmap_52[7:0]) +
	( 15'sd 12622) * $signed(input_fmap_53[7:0]) +
	( 16'sd 29697) * $signed(input_fmap_54[7:0]) +
	( 16'sd 24696) * $signed(input_fmap_55[7:0]) +
	( 14'sd 8165) * $signed(input_fmap_56[7:0]) +
	( 16'sd 27293) * $signed(input_fmap_57[7:0]) +
	( 16'sd 26477) * $signed(input_fmap_58[7:0]) +
	( 16'sd 17672) * $signed(input_fmap_59[7:0]) +
	( 14'sd 7171) * $signed(input_fmap_60[7:0]) +
	( 15'sd 11748) * $signed(input_fmap_61[7:0]) +
	( 13'sd 2378) * $signed(input_fmap_62[7:0]) +
	( 16'sd 24566) * $signed(input_fmap_63[7:0]) +
	( 15'sd 10855) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2551) * $signed(input_fmap_65[7:0]) +
	( 13'sd 3218) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26306) * $signed(input_fmap_67[7:0]) +
	( 14'sd 4436) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20119) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14722) * $signed(input_fmap_70[7:0]) +
	( 16'sd 27715) * $signed(input_fmap_71[7:0]) +
	( 15'sd 12611) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7769) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6570) * $signed(input_fmap_74[7:0]) +
	( 16'sd 30062) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3589) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11355) * $signed(input_fmap_77[7:0]) +
	( 16'sd 24152) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27394) * $signed(input_fmap_79[7:0]) +
	( 15'sd 11031) * $signed(input_fmap_80[7:0]) +
	( 11'sd 638) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24568) * $signed(input_fmap_82[7:0]) +
	( 12'sd 1294) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4753) * $signed(input_fmap_84[7:0]) +
	( 16'sd 24472) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29941) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17586) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17497) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17491) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10535) * $signed(input_fmap_90[7:0]) +
	( 14'sd 5175) * $signed(input_fmap_91[7:0]) +
	( 16'sd 22474) * $signed(input_fmap_92[7:0]) +
	( 16'sd 30290) * $signed(input_fmap_93[7:0]) +
	( 13'sd 2534) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8228) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6954) * $signed(input_fmap_96[7:0]) +
	( 15'sd 15112) * $signed(input_fmap_97[7:0]) +
	( 15'sd 8405) * $signed(input_fmap_98[7:0]) +
	( 16'sd 18755) * $signed(input_fmap_99[7:0]) +
	( 15'sd 12861) * $signed(input_fmap_100[7:0]) +
	( 16'sd 20484) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4698) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10212) * $signed(input_fmap_103[7:0]) +
	( 16'sd 20468) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6690) * $signed(input_fmap_105[7:0]) +
	( 16'sd 18831) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31121) * $signed(input_fmap_107[7:0]) +
	( 12'sd 1110) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9753) * $signed(input_fmap_109[7:0]) +
	( 15'sd 9320) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22329) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29149) * $signed(input_fmap_112[7:0]) +
	( 14'sd 7081) * $signed(input_fmap_113[7:0]) +
	( 15'sd 12230) * $signed(input_fmap_114[7:0]) +
	( 15'sd 15510) * $signed(input_fmap_115[7:0]) +
	( 15'sd 12337) * $signed(input_fmap_116[7:0]) +
	( 11'sd 548) * $signed(input_fmap_117[7:0]) +
	( 14'sd 6162) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31606) * $signed(input_fmap_119[7:0]) +
	( 16'sd 32013) * $signed(input_fmap_120[7:0]) +
	( 16'sd 32423) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19309) * $signed(input_fmap_122[7:0]) +
	( 16'sd 24830) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24812) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30123) * $signed(input_fmap_125[7:0]) +
	( 12'sd 1155) * $signed(input_fmap_126[7:0]) +
	( 16'sd 17569) * $signed(input_fmap_127[7:0]) +
	( 16'sd 27462) * $signed(input_fmap_128[7:0]) +
	( 14'sd 7726) * $signed(input_fmap_129[7:0]) +
	( 16'sd 24814) * $signed(input_fmap_130[7:0]) +
	( 15'sd 14043) * $signed(input_fmap_131[7:0]) +
	( 16'sd 19711) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12538) * $signed(input_fmap_133[7:0]) +
	( 13'sd 3924) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23533) * $signed(input_fmap_135[7:0]) +
	( 16'sd 26928) * $signed(input_fmap_136[7:0]) +
	( 16'sd 16895) * $signed(input_fmap_137[7:0]) +
	( 16'sd 20223) * $signed(input_fmap_138[7:0]) +
	( 16'sd 31952) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9958) * $signed(input_fmap_140[7:0]) +
	( 16'sd 19670) * $signed(input_fmap_141[7:0]) +
	( 14'sd 6617) * $signed(input_fmap_142[7:0]) +
	( 9'sd 160) * $signed(input_fmap_143[7:0]) +
	( 16'sd 16466) * $signed(input_fmap_144[7:0]) +
	( 16'sd 21997) * $signed(input_fmap_145[7:0]) +
	( 16'sd 25110) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13136) * $signed(input_fmap_147[7:0]) +
	( 16'sd 21988) * $signed(input_fmap_148[7:0]) +
	( 13'sd 3563) * $signed(input_fmap_149[7:0]) +
	( 16'sd 28305) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17097) * $signed(input_fmap_151[7:0]) +
	( 16'sd 21456) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11612) * $signed(input_fmap_153[7:0]) +
	( 15'sd 8720) * $signed(input_fmap_154[7:0]) +
	( 14'sd 5987) * $signed(input_fmap_155[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_156[7:0]) +
	( 11'sd 842) * $signed(input_fmap_157[7:0]) +
	( 14'sd 5213) * $signed(input_fmap_158[7:0]) +
	( 16'sd 30639) * $signed(input_fmap_159[7:0]) +
	( 16'sd 22205) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19549) * $signed(input_fmap_161[7:0]) +
	( 13'sd 2665) * $signed(input_fmap_162[7:0]) +
	( 15'sd 10323) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9143) * $signed(input_fmap_164[7:0]) +
	( 16'sd 22544) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30736) * $signed(input_fmap_166[7:0]) +
	( 14'sd 6080) * $signed(input_fmap_167[7:0]) +
	( 13'sd 3625) * $signed(input_fmap_168[7:0]) +
	( 14'sd 8177) * $signed(input_fmap_169[7:0]) +
	( 14'sd 7057) * $signed(input_fmap_170[7:0]) +
	( 16'sd 27528) * $signed(input_fmap_171[7:0]) +
	( 16'sd 22085) * $signed(input_fmap_172[7:0]) +
	( 13'sd 3376) * $signed(input_fmap_173[7:0]) +
	( 16'sd 32718) * $signed(input_fmap_174[7:0]) +
	( 16'sd 29230) * $signed(input_fmap_175[7:0]) +
	( 14'sd 5794) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30487) * $signed(input_fmap_177[7:0]) +
	( 16'sd 18797) * $signed(input_fmap_178[7:0]) +
	( 16'sd 32397) * $signed(input_fmap_179[7:0]) +
	( 16'sd 16878) * $signed(input_fmap_180[7:0]) +
	( 15'sd 13752) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6226) * $signed(input_fmap_182[7:0]) +
	( 15'sd 15885) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8810) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24413) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6837) * $signed(input_fmap_186[7:0]) +
	( 15'sd 11950) * $signed(input_fmap_187[7:0]) +
	( 14'sd 6566) * $signed(input_fmap_188[7:0]) +
	( 14'sd 5653) * $signed(input_fmap_189[7:0]) +
	( 16'sd 18815) * $signed(input_fmap_190[7:0]) +
	( 15'sd 12097) * $signed(input_fmap_191[7:0]) +
	( 16'sd 29716) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29937) * $signed(input_fmap_193[7:0]) +
	( 15'sd 11959) * $signed(input_fmap_194[7:0]) +
	( 13'sd 2744) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7952) * $signed(input_fmap_196[7:0]) +
	( 14'sd 8121) * $signed(input_fmap_197[7:0]) +
	( 16'sd 17555) * $signed(input_fmap_198[7:0]) +
	( 16'sd 23846) * $signed(input_fmap_199[7:0]) +
	( 16'sd 32140) * $signed(input_fmap_200[7:0]) +
	( 14'sd 6195) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18699) * $signed(input_fmap_202[7:0]) +
	( 16'sd 26355) * $signed(input_fmap_203[7:0]) +
	( 16'sd 21473) * $signed(input_fmap_204[7:0]) +
	( 14'sd 6717) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28259) * $signed(input_fmap_206[7:0]) +
	( 16'sd 29402) * $signed(input_fmap_207[7:0]) +
	( 16'sd 31111) * $signed(input_fmap_208[7:0]) +
	( 14'sd 5344) * $signed(input_fmap_209[7:0]) +
	( 16'sd 30921) * $signed(input_fmap_210[7:0]) +
	( 14'sd 6927) * $signed(input_fmap_211[7:0]) +
	( 14'sd 6949) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3707) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30847) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22671) * $signed(input_fmap_215[7:0]) +
	( 13'sd 3120) * $signed(input_fmap_216[7:0]) +
	( 15'sd 16126) * $signed(input_fmap_217[7:0]) +
	( 16'sd 29849) * $signed(input_fmap_218[7:0]) +
	( 12'sd 1474) * $signed(input_fmap_219[7:0]) +
	( 15'sd 9739) * $signed(input_fmap_220[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_221[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2126) * $signed(input_fmap_223[7:0]) +
	( 9'sd 160) * $signed(input_fmap_224[7:0]) +
	( 15'sd 13081) * $signed(input_fmap_225[7:0]) +
	( 15'sd 9116) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22633) * $signed(input_fmap_227[7:0]) +
	( 16'sd 25426) * $signed(input_fmap_228[7:0]) +
	( 15'sd 10750) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18092) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31393) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8450) * $signed(input_fmap_232[7:0]) +
	( 16'sd 29206) * $signed(input_fmap_233[7:0]) +
	( 12'sd 1264) * $signed(input_fmap_234[7:0]) +
	( 16'sd 30166) * $signed(input_fmap_235[7:0]) +
	( 15'sd 14494) * $signed(input_fmap_236[7:0]) +
	( 13'sd 3661) * $signed(input_fmap_237[7:0]) +
	( 16'sd 30319) * $signed(input_fmap_238[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_239[7:0]) +
	( 16'sd 18353) * $signed(input_fmap_240[7:0]) +
	( 16'sd 29858) * $signed(input_fmap_241[7:0]) +
	( 13'sd 2903) * $signed(input_fmap_242[7:0]) +
	( 16'sd 29479) * $signed(input_fmap_243[7:0]) +
	( 16'sd 31182) * $signed(input_fmap_244[7:0]) +
	( 14'sd 4480) * $signed(input_fmap_245[7:0]) +
	( 15'sd 10640) * $signed(input_fmap_246[7:0]) +
	( 15'sd 9775) * $signed(input_fmap_247[7:0]) +
	( 16'sd 23074) * $signed(input_fmap_248[7:0]) +
	( 10'sd 279) * $signed(input_fmap_249[7:0]) +
	( 16'sd 19076) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6993) * $signed(input_fmap_251[7:0]) +
	( 11'sd 746) * $signed(input_fmap_252[7:0]) +
	( 15'sd 15234) * $signed(input_fmap_253[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_254[7:0]) +
	( 14'sd 7256) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_242;
assign conv_mac_242 = 
	( 14'sd 7318) * $signed(input_fmap_0[7:0]) +
	( 16'sd 18037) * $signed(input_fmap_1[7:0]) +
	( 14'sd 7986) * $signed(input_fmap_2[7:0]) +
	( 15'sd 12815) * $signed(input_fmap_3[7:0]) +
	( 15'sd 11590) * $signed(input_fmap_4[7:0]) +
	( 15'sd 13984) * $signed(input_fmap_5[7:0]) +
	( 16'sd 25628) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7388) * $signed(input_fmap_7[7:0]) +
	( 16'sd 17934) * $signed(input_fmap_8[7:0]) +
	( 15'sd 15148) * $signed(input_fmap_9[7:0]) +
	( 16'sd 26387) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11066) * $signed(input_fmap_11[7:0]) +
	( 12'sd 1706) * $signed(input_fmap_12[7:0]) +
	( 16'sd 22732) * $signed(input_fmap_13[7:0]) +
	( 12'sd 1146) * $signed(input_fmap_14[7:0]) +
	( 12'sd 1321) * $signed(input_fmap_15[7:0]) +
	( 16'sd 17745) * $signed(input_fmap_16[7:0]) +
	( 16'sd 27217) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8873) * $signed(input_fmap_18[7:0]) +
	( 16'sd 27839) * $signed(input_fmap_19[7:0]) +
	( 14'sd 8087) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1883) * $signed(input_fmap_21[7:0]) +
	( 16'sd 25708) * $signed(input_fmap_22[7:0]) +
	( 15'sd 14580) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26911) * $signed(input_fmap_24[7:0]) +
	( 15'sd 9559) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20807) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30289) * $signed(input_fmap_27[7:0]) +
	( 16'sd 17918) * $signed(input_fmap_28[7:0]) +
	( 14'sd 7751) * $signed(input_fmap_29[7:0]) +
	( 16'sd 30048) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4692) * $signed(input_fmap_31[7:0]) +
	( 11'sd 582) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29631) * $signed(input_fmap_33[7:0]) +
	( 16'sd 30721) * $signed(input_fmap_34[7:0]) +
	( 16'sd 29370) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29667) * $signed(input_fmap_36[7:0]) +
	( 16'sd 22242) * $signed(input_fmap_37[7:0]) +
	( 14'sd 7112) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17165) * $signed(input_fmap_39[7:0]) +
	( 15'sd 13195) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17053) * $signed(input_fmap_41[7:0]) +
	( 14'sd 4835) * $signed(input_fmap_42[7:0]) +
	( 15'sd 8316) * $signed(input_fmap_43[7:0]) +
	( 16'sd 21798) * $signed(input_fmap_44[7:0]) +
	( 16'sd 17746) * $signed(input_fmap_45[7:0]) +
	( 16'sd 21033) * $signed(input_fmap_46[7:0]) +
	( 15'sd 9755) * $signed(input_fmap_47[7:0]) +
	( 16'sd 22386) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8568) * $signed(input_fmap_49[7:0]) +
	( 16'sd 17215) * $signed(input_fmap_50[7:0]) +
	( 16'sd 26632) * $signed(input_fmap_51[7:0]) +
	( 16'sd 16611) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16043) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16975) * $signed(input_fmap_54[7:0]) +
	( 15'sd 9683) * $signed(input_fmap_55[7:0]) +
	( 12'sd 1744) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23907) * $signed(input_fmap_57[7:0]) +
	( 15'sd 14964) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19785) * $signed(input_fmap_59[7:0]) +
	( 15'sd 9371) * $signed(input_fmap_60[7:0]) +
	( 16'sd 30245) * $signed(input_fmap_61[7:0]) +
	( 16'sd 27065) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23920) * $signed(input_fmap_63[7:0]) +
	( 16'sd 18812) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23208) * $signed(input_fmap_65[7:0]) +
	( 16'sd 29145) * $signed(input_fmap_66[7:0]) +
	( 16'sd 32597) * $signed(input_fmap_67[7:0]) +
	( 15'sd 14898) * $signed(input_fmap_68[7:0]) +
	( 14'sd 7577) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12177) * $signed(input_fmap_70[7:0]) +
	( 16'sd 29735) * $signed(input_fmap_71[7:0]) +
	( 12'sd 1683) * $signed(input_fmap_72[7:0]) +
	( 15'sd 10404) * $signed(input_fmap_73[7:0]) +
	( 14'sd 6200) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24519) * $signed(input_fmap_75[7:0]) +
	( 14'sd 7701) * $signed(input_fmap_76[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_77[7:0]) +
	( 15'sd 11493) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29827) * $signed(input_fmap_79[7:0]) +
	( 16'sd 31525) * $signed(input_fmap_80[7:0]) +
	( 16'sd 18091) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2484) * $signed(input_fmap_82[7:0]) +
	( 16'sd 32472) * $signed(input_fmap_83[7:0]) +
	( 16'sd 28820) * $signed(input_fmap_84[7:0]) +
	( 15'sd 10059) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29529) * $signed(input_fmap_86[7:0]) +
	( 16'sd 23798) * $signed(input_fmap_87[7:0]) +
	( 16'sd 24064) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32303) * $signed(input_fmap_89[7:0]) +
	( 14'sd 6728) * $signed(input_fmap_90[7:0]) +
	( 15'sd 10791) * $signed(input_fmap_91[7:0]) +
	( 16'sd 18426) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24347) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21562) * $signed(input_fmap_94[7:0]) +
	( 15'sd 13517) * $signed(input_fmap_95[7:0]) +
	( 15'sd 15363) * $signed(input_fmap_96[7:0]) +
	( 16'sd 28324) * $signed(input_fmap_97[7:0]) +
	( 13'sd 2625) * $signed(input_fmap_98[7:0]) +
	( 10'sd 295) * $signed(input_fmap_99[7:0]) +
	( 16'sd 24520) * $signed(input_fmap_100[7:0]) +
	( 16'sd 29714) * $signed(input_fmap_101[7:0]) +
	( 16'sd 30529) * $signed(input_fmap_102[7:0]) +
	( 16'sd 29414) * $signed(input_fmap_103[7:0]) +
	( 12'sd 1196) * $signed(input_fmap_104[7:0]) +
	( 16'sd 26369) * $signed(input_fmap_105[7:0]) +
	( 16'sd 24506) * $signed(input_fmap_106[7:0]) +
	( 16'sd 31898) * $signed(input_fmap_107[7:0]) +
	( 15'sd 12678) * $signed(input_fmap_108[7:0]) +
	( 16'sd 30780) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11182) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29918) * $signed(input_fmap_111[7:0]) +
	( 16'sd 22960) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5960) * $signed(input_fmap_113[7:0]) +
	( 13'sd 3955) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31890) * $signed(input_fmap_115[7:0]) +
	( 15'sd 13272) * $signed(input_fmap_116[7:0]) +
	( 16'sd 26230) * $signed(input_fmap_117[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_118[7:0]) +
	( 14'sd 7551) * $signed(input_fmap_119[7:0]) +
	( 15'sd 9823) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30856) * $signed(input_fmap_121[7:0]) +
	( 16'sd 28446) * $signed(input_fmap_122[7:0]) +
	( 16'sd 22610) * $signed(input_fmap_123[7:0]) +
	( 11'sd 869) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25656) * $signed(input_fmap_125[7:0]) +
	( 16'sd 28305) * $signed(input_fmap_126[7:0]) +
	( 16'sd 28334) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23120) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17844) * $signed(input_fmap_129[7:0]) +
	( 16'sd 31505) * $signed(input_fmap_130[7:0]) +
	( 14'sd 4123) * $signed(input_fmap_131[7:0]) +
	( 16'sd 23839) * $signed(input_fmap_132[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_133[7:0]) +
	( 16'sd 31459) * $signed(input_fmap_134[7:0]) +
	( 16'sd 27800) * $signed(input_fmap_135[7:0]) +
	( 15'sd 16193) * $signed(input_fmap_136[7:0]) +
	( 13'sd 3997) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29632) * $signed(input_fmap_138[7:0]) +
	( 16'sd 30258) * $signed(input_fmap_139[7:0]) +
	( 15'sd 8739) * $signed(input_fmap_140[7:0]) +
	( 15'sd 12419) * $signed(input_fmap_141[7:0]) +
	( 16'sd 24970) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20613) * $signed(input_fmap_143[7:0]) +
	( 16'sd 19146) * $signed(input_fmap_144[7:0]) +
	( 16'sd 23969) * $signed(input_fmap_145[7:0]) +
	( 14'sd 6623) * $signed(input_fmap_146[7:0]) +
	( 12'sd 1578) * $signed(input_fmap_147[7:0]) +
	( 11'sd 784) * $signed(input_fmap_148[7:0]) +
	( 16'sd 19960) * $signed(input_fmap_149[7:0]) +
	( 15'sd 9348) * $signed(input_fmap_150[7:0]) +
	( 16'sd 20427) * $signed(input_fmap_151[7:0]) +
	( 16'sd 31640) * $signed(input_fmap_152[7:0]) +
	( 15'sd 11033) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_154[7:0]) +
	( 16'sd 29234) * $signed(input_fmap_155[7:0]) +
	( 16'sd 23876) * $signed(input_fmap_156[7:0]) +
	( 15'sd 8863) * $signed(input_fmap_157[7:0]) +
	( 15'sd 11975) * $signed(input_fmap_158[7:0]) +
	( 16'sd 28869) * $signed(input_fmap_159[7:0]) +
	( 16'sd 19745) * $signed(input_fmap_160[7:0]) +
	( 13'sd 2984) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26799) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2123) * $signed(input_fmap_163[7:0]) +
	( 16'sd 16436) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19059) * $signed(input_fmap_165[7:0]) +
	( 15'sd 14116) * $signed(input_fmap_166[7:0]) +
	( 16'sd 30619) * $signed(input_fmap_167[7:0]) +
	( 15'sd 13012) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30000) * $signed(input_fmap_169[7:0]) +
	( 16'sd 24973) * $signed(input_fmap_170[7:0]) +
	( 7'sd 58) * $signed(input_fmap_171[7:0]) +
	( 15'sd 12663) * $signed(input_fmap_172[7:0]) +
	( 15'sd 8220) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_174[7:0]) +
	( 15'sd 10797) * $signed(input_fmap_175[7:0]) +
	( 16'sd 17985) * $signed(input_fmap_176[7:0]) +
	( 16'sd 25716) * $signed(input_fmap_177[7:0]) +
	( 14'sd 7762) * $signed(input_fmap_178[7:0]) +
	( 16'sd 30986) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32758) * $signed(input_fmap_180[7:0]) +
	( 15'sd 8897) * $signed(input_fmap_181[7:0]) +
	( 15'sd 10256) * $signed(input_fmap_182[7:0]) +
	( 16'sd 20503) * $signed(input_fmap_183[7:0]) +
	( 15'sd 13811) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5396) * $signed(input_fmap_185[7:0]) +
	( 16'sd 18424) * $signed(input_fmap_186[7:0]) +
	( 16'sd 17301) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4651) * $signed(input_fmap_188[7:0]) +
	( 16'sd 28424) * $signed(input_fmap_189[7:0]) +
	( 16'sd 22652) * $signed(input_fmap_190[7:0]) +
	( 15'sd 9153) * $signed(input_fmap_191[7:0]) +
	( 13'sd 2408) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22486) * $signed(input_fmap_193[7:0]) +
	( 16'sd 24168) * $signed(input_fmap_194[7:0]) +
	( 14'sd 5877) * $signed(input_fmap_195[7:0]) +
	( 13'sd 3407) * $signed(input_fmap_196[7:0]) +
	( 16'sd 29676) * $signed(input_fmap_197[7:0]) +
	( 16'sd 30379) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28444) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18957) * $signed(input_fmap_200[7:0]) +
	( 13'sd 4062) * $signed(input_fmap_201[7:0]) +
	( 10'sd 407) * $signed(input_fmap_202[7:0]) +
	( 15'sd 12596) * $signed(input_fmap_203[7:0]) +
	( 15'sd 11394) * $signed(input_fmap_204[7:0]) +
	( 14'sd 5652) * $signed(input_fmap_205[7:0]) +
	( 16'sd 17333) * $signed(input_fmap_206[7:0]) +
	( 16'sd 30934) * $signed(input_fmap_207[7:0]) +
	( 15'sd 12605) * $signed(input_fmap_208[7:0]) +
	( 16'sd 29525) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23026) * $signed(input_fmap_210[7:0]) +
	( 16'sd 22384) * $signed(input_fmap_211[7:0]) +
	( 16'sd 22837) * $signed(input_fmap_212[7:0]) +
	( 15'sd 8689) * $signed(input_fmap_213[7:0]) +
	( 16'sd 24285) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6262) * $signed(input_fmap_215[7:0]) +
	( 16'sd 23856) * $signed(input_fmap_216[7:0]) +
	( 16'sd 18823) * $signed(input_fmap_217[7:0]) +
	( 16'sd 32559) * $signed(input_fmap_218[7:0]) +
	( 15'sd 11729) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24529) * $signed(input_fmap_220[7:0]) +
	( 13'sd 3026) * $signed(input_fmap_221[7:0]) +
	( 14'sd 6696) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12563) * $signed(input_fmap_223[7:0]) +
	( 16'sd 28253) * $signed(input_fmap_224[7:0]) +
	( 14'sd 5129) * $signed(input_fmap_225[7:0]) +
	( 16'sd 30787) * $signed(input_fmap_226[7:0]) +
	( 13'sd 2821) * $signed(input_fmap_227[7:0]) +
	( 16'sd 19633) * $signed(input_fmap_228[7:0]) +
	( 16'sd 24502) * $signed(input_fmap_229[7:0]) +
	( 16'sd 18517) * $signed(input_fmap_230[7:0]) +
	( 14'sd 6363) * $signed(input_fmap_231[7:0]) +
	( 15'sd 16166) * $signed(input_fmap_232[7:0]) +
	( 15'sd 14548) * $signed(input_fmap_233[7:0]) +
	( 16'sd 19763) * $signed(input_fmap_234[7:0]) +
	( 16'sd 17243) * $signed(input_fmap_235[7:0]) +
	( 16'sd 24939) * $signed(input_fmap_236[7:0]) +
	( 16'sd 27851) * $signed(input_fmap_237[7:0]) +
	( 15'sd 9017) * $signed(input_fmap_238[7:0]) +
	( 16'sd 27425) * $signed(input_fmap_239[7:0]) +
	( 15'sd 13186) * $signed(input_fmap_240[7:0]) +
	( 12'sd 2021) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17262) * $signed(input_fmap_242[7:0]) +
	( 10'sd 443) * $signed(input_fmap_243[7:0]) +
	( 16'sd 19990) * $signed(input_fmap_244[7:0]) +
	( 11'sd 706) * $signed(input_fmap_245[7:0]) +
	( 16'sd 20508) * $signed(input_fmap_246[7:0]) +
	( 15'sd 15892) * $signed(input_fmap_247[7:0]) +
	( 14'sd 4528) * $signed(input_fmap_248[7:0]) +
	( 14'sd 7216) * $signed(input_fmap_249[7:0]) +
	( 13'sd 2623) * $signed(input_fmap_250[7:0]) +
	( 15'sd 12403) * $signed(input_fmap_251[7:0]) +
	( 15'sd 9678) * $signed(input_fmap_252[7:0]) +
	( 16'sd 19544) * $signed(input_fmap_253[7:0]) +
	( 15'sd 15636) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24245) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_243;
assign conv_mac_243 = 
	( 13'sd 4062) * $signed(input_fmap_0[7:0]) +
	( 12'sd 1455) * $signed(input_fmap_1[7:0]) +
	( 16'sd 20226) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29857) * $signed(input_fmap_3[7:0]) +
	( 14'sd 6485) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1812) * $signed(input_fmap_5[7:0]) +
	( 16'sd 31287) * $signed(input_fmap_6[7:0]) +
	( 12'sd 1286) * $signed(input_fmap_7[7:0]) +
	( 12'sd 1443) * $signed(input_fmap_8[7:0]) +
	( 12'sd 1111) * $signed(input_fmap_9[7:0]) +
	( 15'sd 15100) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17968) * $signed(input_fmap_11[7:0]) +
	( 16'sd 25671) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11757) * $signed(input_fmap_13[7:0]) +
	( 16'sd 22350) * $signed(input_fmap_14[7:0]) +
	( 16'sd 28075) * $signed(input_fmap_15[7:0]) +
	( 16'sd 28881) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11655) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32399) * $signed(input_fmap_18[7:0]) +
	( 16'sd 25587) * $signed(input_fmap_19[7:0]) +
	( 14'sd 4831) * $signed(input_fmap_20[7:0]) +
	( 16'sd 31133) * $signed(input_fmap_21[7:0]) +
	( 16'sd 23125) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4458) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27727) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14032) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21865) * $signed(input_fmap_26[7:0]) +
	( 8'sd 98) * $signed(input_fmap_27[7:0]) +
	( 16'sd 16607) * $signed(input_fmap_28[7:0]) +
	( 12'sd 1461) * $signed(input_fmap_29[7:0]) +
	( 16'sd 20421) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18554) * $signed(input_fmap_31[7:0]) +
	( 16'sd 20817) * $signed(input_fmap_32[7:0]) +
	( 16'sd 18923) * $signed(input_fmap_33[7:0]) +
	( 16'sd 29457) * $signed(input_fmap_34[7:0]) +
	( 16'sd 24444) * $signed(input_fmap_35[7:0]) +
	( 16'sd 22761) * $signed(input_fmap_36[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_37[7:0]) +
	( 16'sd 30593) * $signed(input_fmap_38[7:0]) +
	( 14'sd 6946) * $signed(input_fmap_39[7:0]) +
	( 13'sd 3531) * $signed(input_fmap_40[7:0]) +
	( 16'sd 21579) * $signed(input_fmap_41[7:0]) +
	( 16'sd 19902) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23476) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17400) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11579) * $signed(input_fmap_45[7:0]) +
	( 15'sd 8414) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3666) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14026) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27441) * $signed(input_fmap_49[7:0]) +
	( 16'sd 30372) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15663) * $signed(input_fmap_51[7:0]) +
	( 16'sd 26531) * $signed(input_fmap_52[7:0]) +
	( 16'sd 31847) * $signed(input_fmap_53[7:0]) +
	( 16'sd 26880) * $signed(input_fmap_54[7:0]) +
	( 13'sd 4008) * $signed(input_fmap_55[7:0]) +
	( 16'sd 31470) * $signed(input_fmap_56[7:0]) +
	( 14'sd 8040) * $signed(input_fmap_57[7:0]) +
	( 13'sd 3086) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26589) * $signed(input_fmap_59[7:0]) +
	( 15'sd 16089) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25746) * $signed(input_fmap_61[7:0]) +
	( 16'sd 26301) * $signed(input_fmap_62[7:0]) +
	( 14'sd 4685) * $signed(input_fmap_63[7:0]) +
	( 14'sd 6166) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10758) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27411) * $signed(input_fmap_66[7:0]) +
	( 16'sd 16995) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5784) * $signed(input_fmap_68[7:0]) +
	( 13'sd 3560) * $signed(input_fmap_69[7:0]) +
	( 14'sd 6505) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30951) * $signed(input_fmap_71[7:0]) +
	( 13'sd 3345) * $signed(input_fmap_72[7:0]) +
	( 15'sd 14527) * $signed(input_fmap_73[7:0]) +
	( 16'sd 28001) * $signed(input_fmap_74[7:0]) +
	( 15'sd 8391) * $signed(input_fmap_75[7:0]) +
	( 16'sd 25003) * $signed(input_fmap_76[7:0]) +
	( 14'sd 7315) * $signed(input_fmap_77[7:0]) +
	( 13'sd 3405) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22366) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19778) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28048) * $signed(input_fmap_81[7:0]) +
	( 16'sd 24204) * $signed(input_fmap_82[7:0]) +
	( 16'sd 23365) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5053) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22094) * $signed(input_fmap_85[7:0]) +
	( 15'sd 11442) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26807) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9036) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2812) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28252) * $signed(input_fmap_90[7:0]) +
	( 11'sd 731) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9446) * $signed(input_fmap_92[7:0]) +
	( 16'sd 31752) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12493) * $signed(input_fmap_94[7:0]) +
	( 14'sd 6971) * $signed(input_fmap_95[7:0]) +
	( 16'sd 16824) * $signed(input_fmap_96[7:0]) +
	( 16'sd 22637) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7958) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29458) * $signed(input_fmap_99[7:0]) +
	( 15'sd 13605) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17160) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27018) * $signed(input_fmap_102[7:0]) +
	( 16'sd 27104) * $signed(input_fmap_103[7:0]) +
	( 13'sd 3227) * $signed(input_fmap_104[7:0]) +
	( 15'sd 13564) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6335) * $signed(input_fmap_106[7:0]) +
	( 15'sd 14476) * $signed(input_fmap_107[7:0]) +
	( 16'sd 22796) * $signed(input_fmap_108[7:0]) +
	( 12'sd 2046) * $signed(input_fmap_109[7:0]) +
	( 12'sd 2022) * $signed(input_fmap_110[7:0]) +
	( 16'sd 17479) * $signed(input_fmap_111[7:0]) +
	( 15'sd 10073) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8709) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11225) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31041) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27637) * $signed(input_fmap_116[7:0]) +
	( 15'sd 15339) * $signed(input_fmap_117[7:0]) +
	( 16'sd 24417) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15444) * $signed(input_fmap_119[7:0]) +
	( 14'sd 6095) * $signed(input_fmap_120[7:0]) +
	( 16'sd 30959) * $signed(input_fmap_121[7:0]) +
	( 16'sd 25505) * $signed(input_fmap_122[7:0]) +
	( 15'sd 10015) * $signed(input_fmap_123[7:0]) +
	( 14'sd 5315) * $signed(input_fmap_124[7:0]) +
	( 16'sd 22753) * $signed(input_fmap_125[7:0]) +
	( 11'sd 920) * $signed(input_fmap_126[7:0]) +
	( 11'sd 647) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15562) * $signed(input_fmap_128[7:0]) +
	( 16'sd 32683) * $signed(input_fmap_129[7:0]) +
	( 16'sd 25052) * $signed(input_fmap_130[7:0]) +
	( 16'sd 21163) * $signed(input_fmap_131[7:0]) +
	( 16'sd 30145) * $signed(input_fmap_132[7:0]) +
	( 13'sd 3825) * $signed(input_fmap_133[7:0]) +
	( 16'sd 22251) * $signed(input_fmap_134[7:0]) +
	( 14'sd 6996) * $signed(input_fmap_135[7:0]) +
	( 14'sd 7955) * $signed(input_fmap_136[7:0]) +
	( 15'sd 10247) * $signed(input_fmap_137[7:0]) +
	( 16'sd 22839) * $signed(input_fmap_138[7:0]) +
	( 16'sd 28841) * $signed(input_fmap_139[7:0]) +
	( 14'sd 6877) * $signed(input_fmap_140[7:0]) +
	( 16'sd 30829) * $signed(input_fmap_141[7:0]) +
	( 12'sd 1785) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31072) * $signed(input_fmap_143[7:0]) +
	( 16'sd 28480) * $signed(input_fmap_144[7:0]) +
	( 15'sd 15535) * $signed(input_fmap_145[7:0]) +
	( 15'sd 15675) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11155) * $signed(input_fmap_147[7:0]) +
	( 16'sd 20732) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25714) * $signed(input_fmap_149[7:0]) +
	( 16'sd 26719) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17201) * $signed(input_fmap_151[7:0]) +
	( 14'sd 4633) * $signed(input_fmap_152[7:0]) +
	( 12'sd 1116) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31160) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30896) * $signed(input_fmap_155[7:0]) +
	( 15'sd 9464) * $signed(input_fmap_156[7:0]) +
	( 16'sd 27863) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20379) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20886) * $signed(input_fmap_159[7:0]) +
	( 16'sd 25860) * $signed(input_fmap_160[7:0]) +
	( 14'sd 7507) * $signed(input_fmap_161[7:0]) +
	( 15'sd 12489) * $signed(input_fmap_162[7:0]) +
	( 14'sd 5827) * $signed(input_fmap_163[7:0]) +
	( 12'sd 1810) * $signed(input_fmap_164[7:0]) +
	( 16'sd 19424) * $signed(input_fmap_165[7:0]) +
	( 16'sd 19152) * $signed(input_fmap_166[7:0]) +
	( 16'sd 29489) * $signed(input_fmap_167[7:0]) +
	( 14'sd 6253) * $signed(input_fmap_168[7:0]) +
	( 15'sd 9106) * $signed(input_fmap_169[7:0]) +
	( 16'sd 20272) * $signed(input_fmap_170[7:0]) +
	( 16'sd 26847) * $signed(input_fmap_171[7:0]) +
	( 16'sd 30742) * $signed(input_fmap_172[7:0]) +
	( 15'sd 13556) * $signed(input_fmap_173[7:0]) +
	( 11'sd 771) * $signed(input_fmap_174[7:0]) +
	( 16'sd 28224) * $signed(input_fmap_175[7:0]) +
	( 16'sd 29355) * $signed(input_fmap_176[7:0]) +
	( 13'sd 2520) * $signed(input_fmap_177[7:0]) +
	( 14'sd 6604) * $signed(input_fmap_178[7:0]) +
	( 14'sd 7021) * $signed(input_fmap_179[7:0]) +
	( 16'sd 17948) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28578) * $signed(input_fmap_181[7:0]) +
	( 15'sd 12881) * $signed(input_fmap_182[7:0]) +
	( 15'sd 8263) * $signed(input_fmap_183[7:0]) +
	( 16'sd 16997) * $signed(input_fmap_184[7:0]) +
	( 16'sd 24450) * $signed(input_fmap_185[7:0]) +
	( 16'sd 30052) * $signed(input_fmap_186[7:0]) +
	( 14'sd 6588) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17668) * $signed(input_fmap_188[7:0]) +
	( 14'sd 6039) * $signed(input_fmap_189[7:0]) +
	( 13'sd 3777) * $signed(input_fmap_190[7:0]) +
	( 16'sd 19028) * $signed(input_fmap_191[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_192[7:0]) +
	( 15'sd 15222) * $signed(input_fmap_193[7:0]) +
	( 16'sd 24219) * $signed(input_fmap_194[7:0]) +
	( 16'sd 20237) * $signed(input_fmap_195[7:0]) +
	( 15'sd 9739) * $signed(input_fmap_196[7:0]) +
	( 16'sd 23996) * $signed(input_fmap_197[7:0]) +
	( 16'sd 26781) * $signed(input_fmap_198[7:0]) +
	( 15'sd 12364) * $signed(input_fmap_199[7:0]) +
	( 16'sd 29088) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15948) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18731) * $signed(input_fmap_202[7:0]) +
	( 14'sd 4445) * $signed(input_fmap_203[7:0]) +
	( 14'sd 5804) * $signed(input_fmap_204[7:0]) +
	( 13'sd 3644) * $signed(input_fmap_205[7:0]) +
	( 16'sd 31294) * $signed(input_fmap_206[7:0]) +
	( 16'sd 24925) * $signed(input_fmap_207[7:0]) +
	( 14'sd 4711) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26318) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5439) * $signed(input_fmap_210[7:0]) +
	( 15'sd 10450) * $signed(input_fmap_211[7:0]) +
	( 12'sd 1310) * $signed(input_fmap_212[7:0]) +
	( 16'sd 30582) * $signed(input_fmap_213[7:0]) +
	( 16'sd 19628) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6592) * $signed(input_fmap_215[7:0]) +
	( 16'sd 17481) * $signed(input_fmap_216[7:0]) +
	( 16'sd 29509) * $signed(input_fmap_217[7:0]) +
	( 16'sd 26610) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19545) * $signed(input_fmap_219[7:0]) +
	( 16'sd 30135) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27046) * $signed(input_fmap_221[7:0]) +
	( 15'sd 14849) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8645) * $signed(input_fmap_223[7:0]) +
	( 16'sd 30699) * $signed(input_fmap_224[7:0]) +
	( 15'sd 12104) * $signed(input_fmap_225[7:0]) +
	( 13'sd 3644) * $signed(input_fmap_226[7:0]) +
	( 15'sd 8853) * $signed(input_fmap_227[7:0]) +
	( 15'sd 12752) * $signed(input_fmap_228[7:0]) +
	( 14'sd 7891) * $signed(input_fmap_229[7:0]) +
	( 14'sd 4750) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14798) * $signed(input_fmap_231[7:0]) +
	( 16'sd 30894) * $signed(input_fmap_232[7:0]) +
	( 14'sd 5034) * $signed(input_fmap_233[7:0]) +
	( 15'sd 16227) * $signed(input_fmap_234[7:0]) +
	( 15'sd 12547) * $signed(input_fmap_235[7:0]) +
	( 15'sd 12357) * $signed(input_fmap_236[7:0]) +
	( 16'sd 31523) * $signed(input_fmap_237[7:0]) +
	( 16'sd 24651) * $signed(input_fmap_238[7:0]) +
	( 16'sd 32061) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22732) * $signed(input_fmap_240[7:0]) +
	( 9'sd 207) * $signed(input_fmap_241[7:0]) +
	( 16'sd 20486) * $signed(input_fmap_242[7:0]) +
	( 16'sd 21507) * $signed(input_fmap_243[7:0]) +
	( 16'sd 25992) * $signed(input_fmap_244[7:0]) +
	( 16'sd 29947) * $signed(input_fmap_245[7:0]) +
	( 15'sd 15468) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3317) * $signed(input_fmap_247[7:0]) +
	( 16'sd 26510) * $signed(input_fmap_248[7:0]) +
	( 16'sd 19233) * $signed(input_fmap_249[7:0]) +
	( 15'sd 16033) * $signed(input_fmap_250[7:0]) +
	( 16'sd 21633) * $signed(input_fmap_251[7:0]) +
	( 16'sd 17646) * $signed(input_fmap_252[7:0]) +
	( 15'sd 11946) * $signed(input_fmap_253[7:0]) +
	( 16'sd 27241) * $signed(input_fmap_254[7:0]) +
	( 16'sd 21398) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_244;
assign conv_mac_244 = 
	( 13'sd 2602) * $signed(input_fmap_0[7:0]) +
	( 15'sd 13794) * $signed(input_fmap_1[7:0]) +
	( 13'sd 3544) * $signed(input_fmap_2[7:0]) +
	( 14'sd 7123) * $signed(input_fmap_3[7:0]) +
	( 16'sd 22430) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27968) * $signed(input_fmap_5[7:0]) +
	( 16'sd 30596) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20160) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7084) * $signed(input_fmap_8[7:0]) +
	( 16'sd 30293) * $signed(input_fmap_9[7:0]) +
	( 16'sd 31245) * $signed(input_fmap_10[7:0]) +
	( 16'sd 27168) * $signed(input_fmap_11[7:0]) +
	( 16'sd 30235) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28171) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18526) * $signed(input_fmap_14[7:0]) +
	( 13'sd 3959) * $signed(input_fmap_15[7:0]) +
	( 13'sd 3760) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23054) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7907) * $signed(input_fmap_18[7:0]) +
	( 16'sd 21095) * $signed(input_fmap_19[7:0]) +
	( 15'sd 9740) * $signed(input_fmap_20[7:0]) +
	( 16'sd 25990) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_22[7:0]) +
	( 14'sd 5850) * $signed(input_fmap_23[7:0]) +
	( 12'sd 1861) * $signed(input_fmap_24[7:0]) +
	( 15'sd 14334) * $signed(input_fmap_25[7:0]) +
	( 15'sd 13240) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8492) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10616) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21483) * $signed(input_fmap_29[7:0]) +
	( 15'sd 12616) * $signed(input_fmap_30[7:0]) +
	( 16'sd 27551) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1424) * $signed(input_fmap_32[7:0]) +
	( 15'sd 12865) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24858) * $signed(input_fmap_34[7:0]) +
	( 15'sd 8572) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30185) * $signed(input_fmap_36[7:0]) +
	( 14'sd 7937) * $signed(input_fmap_37[7:0]) +
	( 16'sd 24522) * $signed(input_fmap_38[7:0]) +
	( 12'sd 2013) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18614) * $signed(input_fmap_40[7:0]) +
	( 16'sd 26163) * $signed(input_fmap_41[7:0]) +
	( 14'sd 6320) * $signed(input_fmap_42[7:0]) +
	( 16'sd 25509) * $signed(input_fmap_43[7:0]) +
	( 16'sd 32381) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4160) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24711) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28204) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28351) * $signed(input_fmap_48[7:0]) +
	( 16'sd 27140) * $signed(input_fmap_49[7:0]) +
	( 14'sd 6809) * $signed(input_fmap_50[7:0]) +
	( 15'sd 15206) * $signed(input_fmap_51[7:0]) +
	( 15'sd 9721) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15912) * $signed(input_fmap_53[7:0]) +
	( 16'sd 28950) * $signed(input_fmap_54[7:0]) +
	( 16'sd 17535) * $signed(input_fmap_55[7:0]) +
	( 16'sd 18506) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13367) * $signed(input_fmap_57[7:0]) +
	( 15'sd 11277) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26565) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30216) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14031) * $signed(input_fmap_61[7:0]) +
	( 16'sd 23438) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13569) * $signed(input_fmap_63[7:0]) +
	( 16'sd 25444) * $signed(input_fmap_64[7:0]) +
	( 16'sd 19263) * $signed(input_fmap_65[7:0]) +
	( 16'sd 25530) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13578) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5953) * $signed(input_fmap_68[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_69[7:0]) +
	( 16'sd 21210) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6033) * $signed(input_fmap_71[7:0]) +
	( 13'sd 2786) * $signed(input_fmap_72[7:0]) +
	( 16'sd 27047) * $signed(input_fmap_73[7:0]) +
	( 16'sd 21159) * $signed(input_fmap_74[7:0]) +
	( 15'sd 13121) * $signed(input_fmap_75[7:0]) +
	( 16'sd 30534) * $signed(input_fmap_76[7:0]) +
	( 16'sd 16504) * $signed(input_fmap_77[7:0]) +
	( 16'sd 31928) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11259) * $signed(input_fmap_79[7:0]) +
	( 16'sd 27298) * $signed(input_fmap_80[7:0]) +
	( 16'sd 19348) * $signed(input_fmap_81[7:0]) +
	( 16'sd 28374) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18547) * $signed(input_fmap_83[7:0]) +
	( 13'sd 3110) * $signed(input_fmap_84[7:0]) +
	( 10'sd 257) * $signed(input_fmap_85[7:0]) +
	( 16'sd 29923) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16923) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5797) * $signed(input_fmap_88[7:0]) +
	( 16'sd 28968) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28567) * $signed(input_fmap_90[7:0]) +
	( 15'sd 13423) * $signed(input_fmap_91[7:0]) +
	( 16'sd 20547) * $signed(input_fmap_92[7:0]) +
	( 16'sd 16800) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14651) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12887) * $signed(input_fmap_95[7:0]) +
	( 15'sd 13155) * $signed(input_fmap_96[7:0]) +
	( 11'sd 860) * $signed(input_fmap_97[7:0]) +
	( 13'sd 3261) * $signed(input_fmap_98[7:0]) +
	( 15'sd 11581) * $signed(input_fmap_99[7:0]) +
	( 14'sd 7555) * $signed(input_fmap_100[7:0]) +
	( 15'sd 8293) * $signed(input_fmap_101[7:0]) +
	( 14'sd 6614) * $signed(input_fmap_102[7:0]) +
	( 15'sd 16001) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12169) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6429) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2320) * $signed(input_fmap_106[7:0]) +
	( 15'sd 16124) * $signed(input_fmap_107[7:0]) +
	( 14'sd 5404) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6958) * $signed(input_fmap_109[7:0]) +
	( 15'sd 12689) * $signed(input_fmap_110[7:0]) +
	( 14'sd 4745) * $signed(input_fmap_111[7:0]) +
	( 14'sd 5500) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4311) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32063) * $signed(input_fmap_114[7:0]) +
	( 16'sd 21927) * $signed(input_fmap_115[7:0]) +
	( 16'sd 22186) * $signed(input_fmap_116[7:0]) +
	( 16'sd 17537) * $signed(input_fmap_117[7:0]) +
	( 13'sd 3511) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17374) * $signed(input_fmap_119[7:0]) +
	( 3'sd 3) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14088) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22918) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20273) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23597) * $signed(input_fmap_124[7:0]) +
	( 16'sd 27020) * $signed(input_fmap_125[7:0]) +
	( 16'sd 29409) * $signed(input_fmap_126[7:0]) +
	( 16'sd 18745) * $signed(input_fmap_127[7:0]) +
	( 12'sd 1851) * $signed(input_fmap_128[7:0]) +
	( 16'sd 26648) * $signed(input_fmap_129[7:0]) +
	( 16'sd 21607) * $signed(input_fmap_130[7:0]) +
	( 16'sd 31744) * $signed(input_fmap_131[7:0]) +
	( 15'sd 12220) * $signed(input_fmap_132[7:0]) +
	( 16'sd 31843) * $signed(input_fmap_133[7:0]) +
	( 13'sd 2735) * $signed(input_fmap_134[7:0]) +
	( 16'sd 25466) * $signed(input_fmap_135[7:0]) +
	( 16'sd 23479) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6356) * $signed(input_fmap_137[7:0]) +
	( 16'sd 28377) * $signed(input_fmap_138[7:0]) +
	( 13'sd 2870) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24797) * $signed(input_fmap_140[7:0]) +
	( 16'sd 22747) * $signed(input_fmap_141[7:0]) +
	( 15'sd 14536) * $signed(input_fmap_142[7:0]) +
	( 13'sd 2533) * $signed(input_fmap_143[7:0]) +
	( 16'sd 24717) * $signed(input_fmap_144[7:0]) +
	( 15'sd 14121) * $signed(input_fmap_145[7:0]) +
	( 15'sd 9769) * $signed(input_fmap_146[7:0]) +
	( 14'sd 4895) * $signed(input_fmap_147[7:0]) +
	( 15'sd 9518) * $signed(input_fmap_148[7:0]) +
	( 12'sd 1295) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23094) * $signed(input_fmap_150[7:0]) +
	( 16'sd 26455) * $signed(input_fmap_151[7:0]) +
	( 16'sd 30987) * $signed(input_fmap_152[7:0]) +
	( 15'sd 10806) * $signed(input_fmap_153[7:0]) +
	( 15'sd 8811) * $signed(input_fmap_154[7:0]) +
	( 16'sd 23548) * $signed(input_fmap_155[7:0]) +
	( 16'sd 17292) * $signed(input_fmap_156[7:0]) +
	( 15'sd 13856) * $signed(input_fmap_157[7:0]) +
	( 15'sd 10263) * $signed(input_fmap_158[7:0]) +
	( 16'sd 27800) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26524) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23043) * $signed(input_fmap_161[7:0]) +
	( 16'sd 25670) * $signed(input_fmap_162[7:0]) +
	( 16'sd 18747) * $signed(input_fmap_163[7:0]) +
	( 15'sd 15462) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9965) * $signed(input_fmap_165[7:0]) +
	( 14'sd 7860) * $signed(input_fmap_166[7:0]) +
	( 15'sd 10956) * $signed(input_fmap_167[7:0]) +
	( 15'sd 9741) * $signed(input_fmap_168[7:0]) +
	( 16'sd 25730) * $signed(input_fmap_169[7:0]) +
	( 13'sd 2875) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31969) * $signed(input_fmap_171[7:0]) +
	( 16'sd 30525) * $signed(input_fmap_172[7:0]) +
	( 15'sd 8729) * $signed(input_fmap_173[7:0]) +
	( 14'sd 6503) * $signed(input_fmap_174[7:0]) +
	( 12'sd 1098) * $signed(input_fmap_175[7:0]) +
	( 15'sd 14551) * $signed(input_fmap_176[7:0]) +
	( 15'sd 8415) * $signed(input_fmap_177[7:0]) +
	( 16'sd 26088) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22424) * $signed(input_fmap_179[7:0]) +
	( 15'sd 8589) * $signed(input_fmap_180[7:0]) +
	( 11'sd 557) * $signed(input_fmap_181[7:0]) +
	( 16'sd 19936) * $signed(input_fmap_182[7:0]) +
	( 15'sd 8416) * $signed(input_fmap_183[7:0]) +
	( 15'sd 15778) * $signed(input_fmap_184[7:0]) +
	( 16'sd 25662) * $signed(input_fmap_185[7:0]) +
	( 15'sd 16107) * $signed(input_fmap_186[7:0]) +
	( 15'sd 9725) * $signed(input_fmap_187[7:0]) +
	( 14'sd 4416) * $signed(input_fmap_188[7:0]) +
	( 16'sd 18210) * $signed(input_fmap_189[7:0]) +
	( 16'sd 17594) * $signed(input_fmap_190[7:0]) +
	( 15'sd 8636) * $signed(input_fmap_191[7:0]) +
	( 16'sd 31216) * $signed(input_fmap_192[7:0]) +
	( 15'sd 11199) * $signed(input_fmap_193[7:0]) +
	( 15'sd 14412) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22432) * $signed(input_fmap_195[7:0]) +
	( 16'sd 27014) * $signed(input_fmap_196[7:0]) +
	( 15'sd 13002) * $signed(input_fmap_197[7:0]) +
	( 16'sd 27419) * $signed(input_fmap_198[7:0]) +
	( 15'sd 11828) * $signed(input_fmap_199[7:0]) +
	( 16'sd 18825) * $signed(input_fmap_200[7:0]) +
	( 16'sd 23719) * $signed(input_fmap_201[7:0]) +
	( 16'sd 30772) * $signed(input_fmap_202[7:0]) +
	( 16'sd 24833) * $signed(input_fmap_203[7:0]) +
	( 13'sd 2966) * $signed(input_fmap_204[7:0]) +
	( 16'sd 27141) * $signed(input_fmap_205[7:0]) +
	( 15'sd 13222) * $signed(input_fmap_206[7:0]) +
	( 15'sd 8773) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22180) * $signed(input_fmap_208[7:0]) +
	( 15'sd 11610) * $signed(input_fmap_209[7:0]) +
	( 16'sd 29760) * $signed(input_fmap_210[7:0]) +
	( 16'sd 27240) * $signed(input_fmap_211[7:0]) +
	( 16'sd 26266) * $signed(input_fmap_212[7:0]) +
	( 14'sd 6244) * $signed(input_fmap_213[7:0]) +
	( 15'sd 9568) * $signed(input_fmap_214[7:0]) +
	( 15'sd 14863) * $signed(input_fmap_215[7:0]) +
	( 16'sd 22230) * $signed(input_fmap_216[7:0]) +
	( 14'sd 4119) * $signed(input_fmap_217[7:0]) +
	( 14'sd 6604) * $signed(input_fmap_218[7:0]) +
	( 16'sd 32044) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14264) * $signed(input_fmap_220[7:0]) +
	( 15'sd 11675) * $signed(input_fmap_221[7:0]) +
	( 16'sd 27595) * $signed(input_fmap_222[7:0]) +
	( 16'sd 29941) * $signed(input_fmap_223[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_224[7:0]) +
	( 15'sd 10149) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22955) * $signed(input_fmap_226[7:0]) +
	( 16'sd 31311) * $signed(input_fmap_227[7:0]) +
	( 16'sd 28194) * $signed(input_fmap_228[7:0]) +
	( 16'sd 30300) * $signed(input_fmap_229[7:0]) +
	( 16'sd 22342) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1940) * $signed(input_fmap_231[7:0]) +
	( 14'sd 5562) * $signed(input_fmap_232[7:0]) +
	( 16'sd 17589) * $signed(input_fmap_233[7:0]) +
	( 16'sd 29314) * $signed(input_fmap_234[7:0]) +
	( 15'sd 15820) * $signed(input_fmap_235[7:0]) +
	( 16'sd 20058) * $signed(input_fmap_236[7:0]) +
	( 10'sd 423) * $signed(input_fmap_237[7:0]) +
	( 16'sd 26152) * $signed(input_fmap_238[7:0]) +
	( 10'sd 410) * $signed(input_fmap_239[7:0]) +
	( 16'sd 20619) * $signed(input_fmap_240[7:0]) +
	( 16'sd 25475) * $signed(input_fmap_241[7:0]) +
	( 16'sd 16701) * $signed(input_fmap_242[7:0]) +
	( 16'sd 18293) * $signed(input_fmap_243[7:0]) +
	( 15'sd 15608) * $signed(input_fmap_244[7:0]) +
	( 15'sd 14043) * $signed(input_fmap_245[7:0]) +
	( 16'sd 19661) * $signed(input_fmap_246[7:0]) +
	( 16'sd 26137) * $signed(input_fmap_247[7:0]) +
	( 14'sd 6391) * $signed(input_fmap_248[7:0]) +
	( 13'sd 2210) * $signed(input_fmap_249[7:0]) +
	( 15'sd 15001) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22121) * $signed(input_fmap_251[7:0]) +
	( 16'sd 25480) * $signed(input_fmap_252[7:0]) +
	( 14'sd 4368) * $signed(input_fmap_253[7:0]) +
	( 16'sd 18792) * $signed(input_fmap_254[7:0]) +
	( 15'sd 12888) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_245;
assign conv_mac_245 = 
	( 16'sd 18559) * $signed(input_fmap_0[7:0]) +
	( 15'sd 9401) * $signed(input_fmap_1[7:0]) +
	( 16'sd 27096) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5165) * $signed(input_fmap_3[7:0]) +
	( 15'sd 13549) * $signed(input_fmap_4[7:0]) +
	( 16'sd 18698) * $signed(input_fmap_5[7:0]) +
	( 15'sd 9022) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20445) * $signed(input_fmap_7[7:0]) +
	( 16'sd 28341) * $signed(input_fmap_8[7:0]) +
	( 16'sd 31645) * $signed(input_fmap_9[7:0]) +
	( 16'sd 19178) * $signed(input_fmap_10[7:0]) +
	( 13'sd 2577) * $signed(input_fmap_11[7:0]) +
	( 15'sd 8799) * $signed(input_fmap_12[7:0]) +
	( 15'sd 10381) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9963) * $signed(input_fmap_14[7:0]) +
	( 16'sd 21963) * $signed(input_fmap_15[7:0]) +
	( 16'sd 30912) * $signed(input_fmap_16[7:0]) +
	( 16'sd 21398) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8256) * $signed(input_fmap_18[7:0]) +
	( 16'sd 19009) * $signed(input_fmap_19[7:0]) +
	( 16'sd 27457) * $signed(input_fmap_20[7:0]) +
	( 16'sd 26851) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19813) * $signed(input_fmap_22[7:0]) +
	( 15'sd 10547) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14061) * $signed(input_fmap_24[7:0]) +
	( 14'sd 6543) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28421) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30204) * $signed(input_fmap_27[7:0]) +
	( 13'sd 2411) * $signed(input_fmap_28[7:0]) +
	( 16'sd 22532) * $signed(input_fmap_29[7:0]) +
	( 11'sd 604) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5184) * $signed(input_fmap_31[7:0]) +
	( 15'sd 8280) * $signed(input_fmap_32[7:0]) +
	( 16'sd 29116) * $signed(input_fmap_33[7:0]) +
	( 16'sd 23730) * $signed(input_fmap_34[7:0]) +
	( 15'sd 13710) * $signed(input_fmap_35[7:0]) +
	( 16'sd 18989) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13773) * $signed(input_fmap_37[7:0]) +
	( 16'sd 29366) * $signed(input_fmap_38[7:0]) +
	( 16'sd 17798) * $signed(input_fmap_39[7:0]) +
	( 16'sd 17432) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28708) * $signed(input_fmap_41[7:0]) +
	( 16'sd 18964) * $signed(input_fmap_42[7:0]) +
	( 16'sd 31385) * $signed(input_fmap_43[7:0]) +
	( 13'sd 3712) * $signed(input_fmap_44[7:0]) +
	( 14'sd 4197) * $signed(input_fmap_45[7:0]) +
	( 16'sd 24444) * $signed(input_fmap_46[7:0]) +
	( 16'sd 24459) * $signed(input_fmap_47[7:0]) +
	( 11'sd 634) * $signed(input_fmap_48[7:0]) +
	( 13'sd 2472) * $signed(input_fmap_49[7:0]) +
	( 16'sd 32101) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2066) * $signed(input_fmap_51[7:0]) +
	( 12'sd 1987) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24253) * $signed(input_fmap_53[7:0]) +
	( 15'sd 15111) * $signed(input_fmap_54[7:0]) +
	( 15'sd 15267) * $signed(input_fmap_55[7:0]) +
	( 13'sd 2335) * $signed(input_fmap_56[7:0]) +
	( 16'sd 24164) * $signed(input_fmap_57[7:0]) +
	( 16'sd 20400) * $signed(input_fmap_58[7:0]) +
	( 15'sd 12411) * $signed(input_fmap_59[7:0]) +
	( 16'sd 30787) * $signed(input_fmap_60[7:0]) +
	( 16'sd 28155) * $signed(input_fmap_61[7:0]) +
	( 11'sd 688) * $signed(input_fmap_62[7:0]) +
	( 16'sd 29520) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24613) * $signed(input_fmap_64[7:0]) +
	( 16'sd 32158) * $signed(input_fmap_65[7:0]) +
	( 15'sd 10499) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7943) * $signed(input_fmap_67[7:0]) +
	( 16'sd 23072) * $signed(input_fmap_68[7:0]) +
	( 13'sd 2416) * $signed(input_fmap_69[7:0]) +
	( 16'sd 19915) * $signed(input_fmap_70[7:0]) +
	( 13'sd 2889) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26986) * $signed(input_fmap_72[7:0]) +
	( 14'sd 8136) * $signed(input_fmap_73[7:0]) +
	( 16'sd 26913) * $signed(input_fmap_74[7:0]) +
	( 16'sd 25804) * $signed(input_fmap_75[7:0]) +
	( 15'sd 15213) * $signed(input_fmap_76[7:0]) +
	( 13'sd 3698) * $signed(input_fmap_77[7:0]) +
	( 11'sd 906) * $signed(input_fmap_78[7:0]) +
	( 15'sd 11184) * $signed(input_fmap_79[7:0]) +
	( 16'sd 21817) * $signed(input_fmap_80[7:0]) +
	( 11'sd 729) * $signed(input_fmap_81[7:0]) +
	( 13'sd 2113) * $signed(input_fmap_82[7:0]) +
	( 14'sd 5666) * $signed(input_fmap_83[7:0]) +
	( 14'sd 6101) * $signed(input_fmap_84[7:0]) +
	( 15'sd 14937) * $signed(input_fmap_85[7:0]) +
	( 15'sd 8761) * $signed(input_fmap_86[7:0]) +
	( 16'sd 26332) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31793) * $signed(input_fmap_88[7:0]) +
	( 15'sd 13712) * $signed(input_fmap_89[7:0]) +
	( 14'sd 5784) * $signed(input_fmap_90[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_91[7:0]) +
	( 15'sd 15493) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24203) * $signed(input_fmap_93[7:0]) +
	( 15'sd 15483) * $signed(input_fmap_94[7:0]) +
	( 15'sd 12432) * $signed(input_fmap_95[7:0]) +
	( 15'sd 8281) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1964) * $signed(input_fmap_97[7:0]) +
	( 16'sd 21980) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22231) * $signed(input_fmap_99[7:0]) +
	( 6'sd 29) * $signed(input_fmap_100[7:0]) +
	( 14'sd 6655) * $signed(input_fmap_101[7:0]) +
	( 15'sd 16005) * $signed(input_fmap_102[7:0]) +
	( 14'sd 4264) * $signed(input_fmap_103[7:0]) +
	( 15'sd 12765) * $signed(input_fmap_104[7:0]) +
	( 16'sd 17600) * $signed(input_fmap_105[7:0]) +
	( 14'sd 4698) * $signed(input_fmap_106[7:0]) +
	( 16'sd 23297) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9361) * $signed(input_fmap_108[7:0]) +
	( 16'sd 29248) * $signed(input_fmap_109[7:0]) +
	( 16'sd 21401) * $signed(input_fmap_110[7:0]) +
	( 16'sd 29109) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24151) * $signed(input_fmap_112[7:0]) +
	( 16'sd 19926) * $signed(input_fmap_113[7:0]) +
	( 16'sd 32265) * $signed(input_fmap_114[7:0]) +
	( 16'sd 19212) * $signed(input_fmap_115[7:0]) +
	( 16'sd 27080) * $signed(input_fmap_116[7:0]) +
	( 11'sd 992) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27238) * $signed(input_fmap_118[7:0]) +
	( 13'sd 2340) * $signed(input_fmap_119[7:0]) +
	( 12'sd 1135) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9218) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1898) * $signed(input_fmap_122[7:0]) +
	( 15'sd 12638) * $signed(input_fmap_123[7:0]) +
	( 15'sd 11554) * $signed(input_fmap_124[7:0]) +
	( 16'sd 28667) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27068) * $signed(input_fmap_126[7:0]) +
	( 16'sd 29291) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13235) * $signed(input_fmap_128[7:0]) +
	( 13'sd 2710) * $signed(input_fmap_129[7:0]) +
	( 14'sd 6428) * $signed(input_fmap_130[7:0]) +
	( 10'sd 335) * $signed(input_fmap_131[7:0]) +
	( 16'sd 25481) * $signed(input_fmap_132[7:0]) +
	( 16'sd 24318) * $signed(input_fmap_133[7:0]) +
	( 15'sd 10079) * $signed(input_fmap_134[7:0]) +
	( 16'sd 30207) * $signed(input_fmap_135[7:0]) +
	( 16'sd 18080) * $signed(input_fmap_136[7:0]) +
	( 14'sd 5791) * $signed(input_fmap_137[7:0]) +
	( 16'sd 29853) * $signed(input_fmap_138[7:0]) +
	( 16'sd 32521) * $signed(input_fmap_139[7:0]) +
	( 16'sd 16447) * $signed(input_fmap_140[7:0]) +
	( 14'sd 4110) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8678) * $signed(input_fmap_142[7:0]) +
	( 16'sd 17135) * $signed(input_fmap_143[7:0]) +
	( 16'sd 31631) * $signed(input_fmap_144[7:0]) +
	( 15'sd 8902) * $signed(input_fmap_145[7:0]) +
	( 14'sd 5861) * $signed(input_fmap_146[7:0]) +
	( 16'sd 30243) * $signed(input_fmap_147[7:0]) +
	( 15'sd 11083) * $signed(input_fmap_148[7:0]) +
	( 16'sd 18757) * $signed(input_fmap_149[7:0]) +
	( 16'sd 18672) * $signed(input_fmap_150[7:0]) +
	( 16'sd 20523) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7854) * $signed(input_fmap_152[7:0]) +
	( 16'sd 20988) * $signed(input_fmap_153[7:0]) +
	( 16'sd 17942) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10551) * $signed(input_fmap_155[7:0]) +
	( 16'sd 18124) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23941) * $signed(input_fmap_157[7:0]) +
	( 16'sd 23129) * $signed(input_fmap_158[7:0]) +
	( 16'sd 29122) * $signed(input_fmap_159[7:0]) +
	( 15'sd 8590) * $signed(input_fmap_160[7:0]) +
	( 15'sd 8489) * $signed(input_fmap_161[7:0]) +
	( 16'sd 26052) * $signed(input_fmap_162[7:0]) +
	( 15'sd 11584) * $signed(input_fmap_163[7:0]) +
	( 15'sd 8528) * $signed(input_fmap_164[7:0]) +
	( 15'sd 9815) * $signed(input_fmap_165[7:0]) +
	( 13'sd 3692) * $signed(input_fmap_166[7:0]) +
	( 16'sd 24731) * $signed(input_fmap_167[7:0]) +
	( 14'sd 5520) * $signed(input_fmap_168[7:0]) +
	( 16'sd 29874) * $signed(input_fmap_169[7:0]) +
	( 16'sd 32021) * $signed(input_fmap_170[7:0]) +
	( 13'sd 4058) * $signed(input_fmap_171[7:0]) +
	( 16'sd 24250) * $signed(input_fmap_172[7:0]) +
	( 14'sd 6036) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7336) * $signed(input_fmap_174[7:0]) +
	( 15'sd 13908) * $signed(input_fmap_175[7:0]) +
	( 14'sd 4700) * $signed(input_fmap_176[7:0]) +
	( 16'sd 28868) * $signed(input_fmap_177[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_178[7:0]) +
	( 13'sd 3864) * $signed(input_fmap_179[7:0]) +
	( 15'sd 14527) * $signed(input_fmap_180[7:0]) +
	( 16'sd 30287) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26347) * $signed(input_fmap_182[7:0]) +
	( 12'sd 1537) * $signed(input_fmap_183[7:0]) +
	( 16'sd 21892) * $signed(input_fmap_184[7:0]) +
	( 16'sd 31290) * $signed(input_fmap_185[7:0]) +
	( 16'sd 16526) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5400) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32214) * $signed(input_fmap_188[7:0]) +
	( 16'sd 25228) * $signed(input_fmap_189[7:0]) +
	( 16'sd 28000) * $signed(input_fmap_190[7:0]) +
	( 16'sd 29131) * $signed(input_fmap_191[7:0]) +
	( 13'sd 3716) * $signed(input_fmap_192[7:0]) +
	( 16'sd 27800) * $signed(input_fmap_193[7:0]) +
	( 14'sd 8110) * $signed(input_fmap_194[7:0]) +
	( 3'sd 3) * $signed(input_fmap_195[7:0]) +
	( 16'sd 16957) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26421) * $signed(input_fmap_197[7:0]) +
	( 15'sd 11277) * $signed(input_fmap_198[7:0]) +
	( 15'sd 8777) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3656) * $signed(input_fmap_200[7:0]) +
	( 16'sd 16634) * $signed(input_fmap_201[7:0]) +
	( 15'sd 10235) * $signed(input_fmap_202[7:0]) +
	( 16'sd 17446) * $signed(input_fmap_203[7:0]) +
	( 16'sd 29484) * $signed(input_fmap_204[7:0]) +
	( 15'sd 9909) * $signed(input_fmap_205[7:0]) +
	( 15'sd 9109) * $signed(input_fmap_206[7:0]) +
	( 15'sd 10794) * $signed(input_fmap_207[7:0]) +
	( 16'sd 32668) * $signed(input_fmap_208[7:0]) +
	( 11'sd 834) * $signed(input_fmap_209[7:0]) +
	( 16'sd 32165) * $signed(input_fmap_210[7:0]) +
	( 15'sd 9978) * $signed(input_fmap_211[7:0]) +
	( 13'sd 3402) * $signed(input_fmap_212[7:0]) +
	( 14'sd 8120) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30213) * $signed(input_fmap_214[7:0]) +
	( 14'sd 7435) * $signed(input_fmap_215[7:0]) +
	( 16'sd 19954) * $signed(input_fmap_216[7:0]) +
	( 16'sd 32044) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22774) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5390) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14437) * $signed(input_fmap_220[7:0]) +
	( 15'sd 14915) * $signed(input_fmap_221[7:0]) +
	( 16'sd 29873) * $signed(input_fmap_222[7:0]) +
	( 15'sd 8388) * $signed(input_fmap_223[7:0]) +
	( 15'sd 15960) * $signed(input_fmap_224[7:0]) +
	( 16'sd 24412) * $signed(input_fmap_225[7:0]) +
	( 14'sd 7051) * $signed(input_fmap_226[7:0]) +
	( 16'sd 22276) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26703) * $signed(input_fmap_228[7:0]) +
	( 16'sd 27921) * $signed(input_fmap_229[7:0]) +
	( 14'sd 8079) * $signed(input_fmap_230[7:0]) +
	( 16'sd 31075) * $signed(input_fmap_231[7:0]) +
	( 16'sd 27477) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21637) * $signed(input_fmap_233[7:0]) +
	( 16'sd 17540) * $signed(input_fmap_234[7:0]) +
	( 16'sd 19936) * $signed(input_fmap_235[7:0]) +
	( 16'sd 30784) * $signed(input_fmap_236[7:0]) +
	( 13'sd 2642) * $signed(input_fmap_237[7:0]) +
	( 11'sd 651) * $signed(input_fmap_238[7:0]) +
	( 16'sd 17637) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22845) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7515) * $signed(input_fmap_241[7:0]) +
	( 16'sd 30458) * $signed(input_fmap_242[7:0]) +
	( 15'sd 9734) * $signed(input_fmap_243[7:0]) +
	( 10'sd 288) * $signed(input_fmap_244[7:0]) +
	( 16'sd 31564) * $signed(input_fmap_245[7:0]) +
	( 15'sd 8697) * $signed(input_fmap_246[7:0]) +
	( 15'sd 11501) * $signed(input_fmap_247[7:0]) +
	( 16'sd 21022) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28415) * $signed(input_fmap_249[7:0]) +
	( 16'sd 25865) * $signed(input_fmap_250[7:0]) +
	( 16'sd 27060) * $signed(input_fmap_251[7:0]) +
	( 16'sd 18151) * $signed(input_fmap_252[7:0]) +
	( 14'sd 5867) * $signed(input_fmap_253[7:0]) +
	( 16'sd 23045) * $signed(input_fmap_254[7:0]) +
	( 10'sd 511) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_246;
assign conv_mac_246 = 
	( 16'sd 25276) * $signed(input_fmap_0[7:0]) +
	( 15'sd 14105) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31530) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28019) * $signed(input_fmap_3[7:0]) +
	( 16'sd 24270) * $signed(input_fmap_4[7:0]) +
	( 16'sd 19990) * $signed(input_fmap_5[7:0]) +
	( 16'sd 23556) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19247) * $signed(input_fmap_7[7:0]) +
	( 16'sd 27773) * $signed(input_fmap_8[7:0]) +
	( 16'sd 29638) * $signed(input_fmap_9[7:0]) +
	( 15'sd 8345) * $signed(input_fmap_10[7:0]) +
	( 14'sd 6212) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5270) * $signed(input_fmap_12[7:0]) +
	( 16'sd 23164) * $signed(input_fmap_13[7:0]) +
	( 16'sd 18865) * $signed(input_fmap_14[7:0]) +
	( 14'sd 7704) * $signed(input_fmap_15[7:0]) +
	( 16'sd 25759) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26383) * $signed(input_fmap_17[7:0]) +
	( 16'sd 31296) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5686) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31854) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1794) * $signed(input_fmap_21[7:0]) +
	( 15'sd 13121) * $signed(input_fmap_22[7:0]) +
	( 15'sd 15506) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4407) * $signed(input_fmap_24[7:0]) +
	( 16'sd 17543) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15706) * $signed(input_fmap_26[7:0]) +
	( 16'sd 30581) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14506) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23998) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19780) * $signed(input_fmap_30[7:0]) +
	( 16'sd 21334) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9860) * $signed(input_fmap_32[7:0]) +
	( 16'sd 24336) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3401) * $signed(input_fmap_34[7:0]) +
	( 15'sd 15428) * $signed(input_fmap_35[7:0]) +
	( 16'sd 31579) * $signed(input_fmap_36[7:0]) +
	( 14'sd 5706) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18855) * $signed(input_fmap_38[7:0]) +
	( 16'sd 25706) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25381) * $signed(input_fmap_40[7:0]) +
	( 15'sd 15267) * $signed(input_fmap_41[7:0]) +
	( 16'sd 26392) * $signed(input_fmap_42[7:0]) +
	( 13'sd 3027) * $signed(input_fmap_43[7:0]) +
	( 11'sd 799) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11956) * $signed(input_fmap_45[7:0]) +
	( 16'sd 25335) * $signed(input_fmap_46[7:0]) +
	( 16'sd 31719) * $signed(input_fmap_47[7:0]) +
	( 13'sd 3797) * $signed(input_fmap_48[7:0]) +
	( 16'sd 19433) * $signed(input_fmap_49[7:0]) +
	( 15'sd 15030) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32412) * $signed(input_fmap_51[7:0]) +
	( 15'sd 8631) * $signed(input_fmap_52[7:0]) +
	( 16'sd 30298) * $signed(input_fmap_53[7:0]) +
	( 15'sd 13730) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19585) * $signed(input_fmap_55[7:0]) +
	( 14'sd 5924) * $signed(input_fmap_56[7:0]) +
	( 16'sd 21773) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19895) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26841) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11850) * $signed(input_fmap_60[7:0]) +
	( 16'sd 19715) * $signed(input_fmap_61[7:0]) +
	( 15'sd 9027) * $signed(input_fmap_62[7:0]) +
	( 15'sd 10446) * $signed(input_fmap_63[7:0]) +
	( 16'sd 20782) * $signed(input_fmap_64[7:0]) +
	( 16'sd 23071) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14943) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13619) * $signed(input_fmap_67[7:0]) +
	( 13'sd 3722) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8919) * $signed(input_fmap_69[7:0]) +
	( 15'sd 12731) * $signed(input_fmap_70[7:0]) +
	( 16'sd 25948) * $signed(input_fmap_71[7:0]) +
	( 16'sd 26613) * $signed(input_fmap_72[7:0]) +
	( 14'sd 4210) * $signed(input_fmap_73[7:0]) +
	( 16'sd 31963) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29020) * $signed(input_fmap_75[7:0]) +
	( 15'sd 12194) * $signed(input_fmap_76[7:0]) +
	( 15'sd 9567) * $signed(input_fmap_77[7:0]) +
	( 16'sd 22843) * $signed(input_fmap_78[7:0]) +
	( 14'sd 4730) * $signed(input_fmap_79[7:0]) +
	( 8'sd 114) * $signed(input_fmap_80[7:0]) +
	( 12'sd 1648) * $signed(input_fmap_81[7:0]) +
	( 14'sd 6235) * $signed(input_fmap_82[7:0]) +
	( 15'sd 9699) * $signed(input_fmap_83[7:0]) +
	( 14'sd 4399) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21392) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20732) * $signed(input_fmap_86[7:0]) +
	( 16'sd 18969) * $signed(input_fmap_87[7:0]) +
	( 16'sd 17686) * $signed(input_fmap_88[7:0]) +
	( 16'sd 17618) * $signed(input_fmap_89[7:0]) +
	( 16'sd 23359) * $signed(input_fmap_90[7:0]) +
	( 15'sd 11106) * $signed(input_fmap_91[7:0]) +
	( 15'sd 9225) * $signed(input_fmap_92[7:0]) +
	( 16'sd 21198) * $signed(input_fmap_93[7:0]) +
	( 16'sd 32612) * $signed(input_fmap_94[7:0]) +
	( 15'sd 15915) * $signed(input_fmap_95[7:0]) +
	( 13'sd 2637) * $signed(input_fmap_96[7:0]) +
	( 16'sd 17078) * $signed(input_fmap_97[7:0]) +
	( 15'sd 15731) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7321) * $signed(input_fmap_99[7:0]) +
	( 15'sd 16299) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16772) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23749) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15379) * $signed(input_fmap_103[7:0]) +
	( 14'sd 8039) * $signed(input_fmap_104[7:0]) +
	( 16'sd 31379) * $signed(input_fmap_105[7:0]) +
	( 15'sd 13988) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7348) * $signed(input_fmap_107[7:0]) +
	( 16'sd 27202) * $signed(input_fmap_108[7:0]) +
	( 16'sd 19538) * $signed(input_fmap_109[7:0]) +
	( 14'sd 8179) * $signed(input_fmap_110[7:0]) +
	( 16'sd 23950) * $signed(input_fmap_111[7:0]) +
	( 14'sd 4944) * $signed(input_fmap_112[7:0]) +
	( 16'sd 31174) * $signed(input_fmap_113[7:0]) +
	( 16'sd 27282) * $signed(input_fmap_114[7:0]) +
	( 15'sd 11068) * $signed(input_fmap_115[7:0]) +
	( 16'sd 23214) * $signed(input_fmap_116[7:0]) +
	( 15'sd 13742) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20840) * $signed(input_fmap_118[7:0]) +
	( 15'sd 8584) * $signed(input_fmap_119[7:0]) +
	( 16'sd 28617) * $signed(input_fmap_120[7:0]) +
	( 15'sd 9149) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27113) * $signed(input_fmap_122[7:0]) +
	( 11'sd 902) * $signed(input_fmap_123[7:0]) +
	( 16'sd 24097) * $signed(input_fmap_124[7:0]) +
	( 15'sd 13751) * $signed(input_fmap_125[7:0]) +
	( 10'sd 376) * $signed(input_fmap_126[7:0]) +
	( 15'sd 13366) * $signed(input_fmap_127[7:0]) +
	( 16'sd 23680) * $signed(input_fmap_128[7:0]) +
	( 14'sd 6071) * $signed(input_fmap_129[7:0]) +
	( 15'sd 15130) * $signed(input_fmap_130[7:0]) +
	( 13'sd 2534) * $signed(input_fmap_131[7:0]) +
	( 9'sd 251) * $signed(input_fmap_132[7:0]) +
	( 16'sd 32606) * $signed(input_fmap_133[7:0]) +
	( 16'sd 23673) * $signed(input_fmap_134[7:0]) +
	( 16'sd 21730) * $signed(input_fmap_135[7:0]) +
	( 16'sd 25336) * $signed(input_fmap_136[7:0]) +
	( 16'sd 26467) * $signed(input_fmap_137[7:0]) +
	( 14'sd 6135) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14245) * $signed(input_fmap_139[7:0]) +
	( 16'sd 20127) * $signed(input_fmap_140[7:0]) +
	( 16'sd 18346) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19880) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31231) * $signed(input_fmap_143[7:0]) +
	( 12'sd 1647) * $signed(input_fmap_144[7:0]) +
	( 15'sd 13851) * $signed(input_fmap_145[7:0]) +
	( 16'sd 16717) * $signed(input_fmap_146[7:0]) +
	( 15'sd 8732) * $signed(input_fmap_147[7:0]) +
	( 14'sd 5957) * $signed(input_fmap_148[7:0]) +
	( 14'sd 6287) * $signed(input_fmap_149[7:0]) +
	( 16'sd 29097) * $signed(input_fmap_150[7:0]) +
	( 14'sd 4524) * $signed(input_fmap_151[7:0]) +
	( 15'sd 14529) * $signed(input_fmap_152[7:0]) +
	( 16'sd 20791) * $signed(input_fmap_153[7:0]) +
	( 16'sd 20172) * $signed(input_fmap_154[7:0]) +
	( 16'sd 22893) * $signed(input_fmap_155[7:0]) +
	( 13'sd 2570) * $signed(input_fmap_156[7:0]) +
	( 15'sd 11440) * $signed(input_fmap_157[7:0]) +
	( 15'sd 14025) * $signed(input_fmap_158[7:0]) +
	( 16'sd 31184) * $signed(input_fmap_159[7:0]) +
	( 16'sd 21270) * $signed(input_fmap_160[7:0]) +
	( 13'sd 4075) * $signed(input_fmap_161[7:0]) +
	( 14'sd 6275) * $signed(input_fmap_162[7:0]) +
	( 16'sd 26704) * $signed(input_fmap_163[7:0]) +
	( 16'sd 24064) * $signed(input_fmap_164[7:0]) +
	( 16'sd 16411) * $signed(input_fmap_165[7:0]) +
	( 16'sd 17378) * $signed(input_fmap_166[7:0]) +
	( 16'sd 26851) * $signed(input_fmap_167[7:0]) +
	( 15'sd 15812) * $signed(input_fmap_168[7:0]) +
	( 15'sd 16277) * $signed(input_fmap_169[7:0]) +
	( 16'sd 27532) * $signed(input_fmap_170[7:0]) +
	( 14'sd 4936) * $signed(input_fmap_171[7:0]) +
	( 15'sd 10925) * $signed(input_fmap_172[7:0]) +
	( 16'sd 24209) * $signed(input_fmap_173[7:0]) +
	( 16'sd 26514) * $signed(input_fmap_174[7:0]) +
	( 14'sd 4196) * $signed(input_fmap_175[7:0]) +
	( 16'sd 24665) * $signed(input_fmap_176[7:0]) +
	( 16'sd 27493) * $signed(input_fmap_177[7:0]) +
	( 12'sd 1835) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25867) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32036) * $signed(input_fmap_180[7:0]) +
	( 15'sd 11828) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30416) * $signed(input_fmap_182[7:0]) +
	( 14'sd 7196) * $signed(input_fmap_183[7:0]) +
	( 15'sd 8321) * $signed(input_fmap_184[7:0]) +
	( 15'sd 11917) * $signed(input_fmap_185[7:0]) +
	( 14'sd 6793) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4162) * $signed(input_fmap_187[7:0]) +
	( 16'sd 25101) * $signed(input_fmap_188[7:0]) +
	( 13'sd 2332) * $signed(input_fmap_189[7:0]) +
	( 15'sd 15062) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20961) * $signed(input_fmap_191[7:0]) +
	( 16'sd 24356) * $signed(input_fmap_192[7:0]) +
	( 16'sd 20438) * $signed(input_fmap_193[7:0]) +
	( 11'sd 539) * $signed(input_fmap_194[7:0]) +
	( 16'sd 25754) * $signed(input_fmap_195[7:0]) +
	( 16'sd 31370) * $signed(input_fmap_196[7:0]) +
	( 15'sd 10570) * $signed(input_fmap_197[7:0]) +
	( 16'sd 20542) * $signed(input_fmap_198[7:0]) +
	( 16'sd 28303) * $signed(input_fmap_199[7:0]) +
	( 12'sd 1443) * $signed(input_fmap_200[7:0]) +
	( 15'sd 8614) * $signed(input_fmap_201[7:0]) +
	( 16'sd 18135) * $signed(input_fmap_202[7:0]) +
	( 12'sd 1436) * $signed(input_fmap_203[7:0]) +
	( 16'sd 32221) * $signed(input_fmap_204[7:0]) +
	( 15'sd 12720) * $signed(input_fmap_205[7:0]) +
	( 16'sd 17612) * $signed(input_fmap_206[7:0]) +
	( 16'sd 21621) * $signed(input_fmap_207[7:0]) +
	( 16'sd 22974) * $signed(input_fmap_208[7:0]) +
	( 16'sd 28391) * $signed(input_fmap_209[7:0]) +
	( 15'sd 11000) * $signed(input_fmap_210[7:0]) +
	( 15'sd 13459) * $signed(input_fmap_211[7:0]) +
	( 15'sd 12747) * $signed(input_fmap_212[7:0]) +
	( 15'sd 11606) * $signed(input_fmap_213[7:0]) +
	( 15'sd 10292) * $signed(input_fmap_214[7:0]) +
	( 12'sd 1928) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24328) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9549) * $signed(input_fmap_217[7:0]) +
	( 16'sd 20457) * $signed(input_fmap_218[7:0]) +
	( 16'sd 30949) * $signed(input_fmap_219[7:0]) +
	( 12'sd 1184) * $signed(input_fmap_220[7:0]) +
	( 16'sd 24874) * $signed(input_fmap_221[7:0]) +
	( 16'sd 31142) * $signed(input_fmap_222[7:0]) +
	( 15'sd 14618) * $signed(input_fmap_223[7:0]) +
	( 16'sd 23686) * $signed(input_fmap_224[7:0]) +
	( 14'sd 6191) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22210) * $signed(input_fmap_226[7:0]) +
	( 16'sd 31901) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1178) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20768) * $signed(input_fmap_229[7:0]) +
	( 16'sd 30193) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17140) * $signed(input_fmap_231[7:0]) +
	( 16'sd 28019) * $signed(input_fmap_232[7:0]) +
	( 16'sd 24526) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15452) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3180) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28049) * $signed(input_fmap_236[7:0]) +
	( 10'sd 286) * $signed(input_fmap_237[7:0]) +
	( 16'sd 31282) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19325) * $signed(input_fmap_239[7:0]) +
	( 16'sd 20816) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18647) * $signed(input_fmap_241[7:0]) +
	( 16'sd 29828) * $signed(input_fmap_242[7:0]) +
	( 14'sd 4579) * $signed(input_fmap_243[7:0]) +
	( 16'sd 26663) * $signed(input_fmap_244[7:0]) +
	( 13'sd 2700) * $signed(input_fmap_245[7:0]) +
	( 16'sd 23616) * $signed(input_fmap_246[7:0]) +
	( 16'sd 30705) * $signed(input_fmap_247[7:0]) +
	( 16'sd 22350) * $signed(input_fmap_248[7:0]) +
	( 15'sd 12675) * $signed(input_fmap_249[7:0]) +
	( 15'sd 12505) * $signed(input_fmap_250[7:0]) +
	( 12'sd 1931) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5239) * $signed(input_fmap_252[7:0]) +
	( 16'sd 19974) * $signed(input_fmap_253[7:0]) +
	( 16'sd 31909) * $signed(input_fmap_254[7:0]) +
	( 16'sd 24829) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_247;
assign conv_mac_247 = 
	( 7'sd 63) * $signed(input_fmap_0[7:0]) +
	( 15'sd 10371) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25164) * $signed(input_fmap_2[7:0]) +
	( 16'sd 16653) * $signed(input_fmap_3[7:0]) +
	( 16'sd 21339) * $signed(input_fmap_4[7:0]) +
	( 14'sd 7238) * $signed(input_fmap_5[7:0]) +
	( 15'sd 8931) * $signed(input_fmap_6[7:0]) +
	( 16'sd 20678) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18516) * $signed(input_fmap_8[7:0]) +
	( 16'sd 20200) * $signed(input_fmap_9[7:0]) +
	( 14'sd 5095) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14363) * $signed(input_fmap_11[7:0]) +
	( 11'sd 921) * $signed(input_fmap_12[7:0]) +
	( 16'sd 20572) * $signed(input_fmap_13[7:0]) +
	( 15'sd 12531) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29396) * $signed(input_fmap_15[7:0]) +
	( 14'sd 5818) * $signed(input_fmap_16[7:0]) +
	( 16'sd 25369) * $signed(input_fmap_17[7:0]) +
	( 15'sd 8507) * $signed(input_fmap_18[7:0]) +
	( 16'sd 23902) * $signed(input_fmap_19[7:0]) +
	( 16'sd 26958) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12093) * $signed(input_fmap_21[7:0]) +
	( 16'sd 19538) * $signed(input_fmap_22[7:0]) +
	( 15'sd 9913) * $signed(input_fmap_23[7:0]) +
	( 16'sd 24507) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12217) * $signed(input_fmap_25[7:0]) +
	( 16'sd 18092) * $signed(input_fmap_26[7:0]) +
	( 14'sd 6994) * $signed(input_fmap_27[7:0]) +
	( 15'sd 10372) * $signed(input_fmap_28[7:0]) +
	( 16'sd 25086) * $signed(input_fmap_29[7:0]) +
	( 15'sd 8538) * $signed(input_fmap_30[7:0]) +
	( 16'sd 16698) * $signed(input_fmap_31[7:0]) +
	( 16'sd 29646) * $signed(input_fmap_32[7:0]) +
	( 12'sd 1944) * $signed(input_fmap_33[7:0]) +
	( 11'sd 693) * $signed(input_fmap_34[7:0]) +
	( 15'sd 9671) * $signed(input_fmap_35[7:0]) +
	( 11'sd 546) * $signed(input_fmap_36[7:0]) +
	( 16'sd 25154) * $signed(input_fmap_37[7:0]) +
	( 16'sd 18899) * $signed(input_fmap_38[7:0]) +
	( 16'sd 30377) * $signed(input_fmap_39[7:0]) +
	( 16'sd 24568) * $signed(input_fmap_40[7:0]) +
	( 14'sd 4944) * $signed(input_fmap_41[7:0]) +
	( 16'sd 30546) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26894) * $signed(input_fmap_43[7:0]) +
	( 16'sd 29737) * $signed(input_fmap_44[7:0]) +
	( 15'sd 15107) * $signed(input_fmap_45[7:0]) +
	( 14'sd 5924) * $signed(input_fmap_46[7:0]) +
	( 16'sd 29371) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19248) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8688) * $signed(input_fmap_49[7:0]) +
	( 14'sd 5204) * $signed(input_fmap_50[7:0]) +
	( 15'sd 12745) * $signed(input_fmap_51[7:0]) +
	( 14'sd 5410) * $signed(input_fmap_52[7:0]) +
	( 14'sd 7271) * $signed(input_fmap_53[7:0]) +
	( 14'sd 6574) * $signed(input_fmap_54[7:0]) +
	( 16'sd 31323) * $signed(input_fmap_55[7:0]) +
	( 11'sd 607) * $signed(input_fmap_56[7:0]) +
	( 16'sd 29696) * $signed(input_fmap_57[7:0]) +
	( 16'sd 18421) * $signed(input_fmap_58[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_59[7:0]) +
	( 16'sd 27974) * $signed(input_fmap_60[7:0]) +
	( 15'sd 14187) * $signed(input_fmap_61[7:0]) +
	( 16'sd 17888) * $signed(input_fmap_62[7:0]) +
	( 15'sd 9067) * $signed(input_fmap_63[7:0]) +
	( 16'sd 19943) * $signed(input_fmap_64[7:0]) +
	( 14'sd 6819) * $signed(input_fmap_65[7:0]) +
	( 16'sd 26051) * $signed(input_fmap_66[7:0]) +
	( 15'sd 12761) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9413) * $signed(input_fmap_68[7:0]) +
	( 15'sd 8302) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5584) * $signed(input_fmap_70[7:0]) +
	( 16'sd 19107) * $signed(input_fmap_71[7:0]) +
	( 16'sd 17889) * $signed(input_fmap_72[7:0]) +
	( 16'sd 32562) * $signed(input_fmap_73[7:0]) +
	( 16'sd 17418) * $signed(input_fmap_74[7:0]) +
	( 12'sd 1291) * $signed(input_fmap_75[7:0]) +
	( 15'sd 10807) * $signed(input_fmap_76[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_77[7:0]) +
	( 16'sd 18157) * $signed(input_fmap_78[7:0]) +
	( 16'sd 22609) * $signed(input_fmap_79[7:0]) +
	( 13'sd 2127) * $signed(input_fmap_80[7:0]) +
	( 16'sd 23611) * $signed(input_fmap_81[7:0]) +
	( 14'sd 7705) * $signed(input_fmap_82[7:0]) +
	( 16'sd 19549) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15407) * $signed(input_fmap_84[7:0]) +
	( 16'sd 25488) * $signed(input_fmap_85[7:0]) +
	( 13'sd 4035) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17686) * $signed(input_fmap_87[7:0]) +
	( 16'sd 31700) * $signed(input_fmap_88[7:0]) +
	( 14'sd 7230) * $signed(input_fmap_89[7:0]) +
	( 16'sd 22035) * $signed(input_fmap_90[7:0]) +
	( 15'sd 9401) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16448) * $signed(input_fmap_92[7:0]) +
	( 15'sd 15878) * $signed(input_fmap_93[7:0]) +
	( 16'sd 16770) * $signed(input_fmap_94[7:0]) +
	( 11'sd 834) * $signed(input_fmap_95[7:0]) +
	( 16'sd 32266) * $signed(input_fmap_96[7:0]) +
	( 15'sd 14151) * $signed(input_fmap_97[7:0]) +
	( 16'sd 28223) * $signed(input_fmap_98[7:0]) +
	( 16'sd 22706) * $signed(input_fmap_99[7:0]) +
	( 16'sd 17335) * $signed(input_fmap_100[7:0]) +
	( 16'sd 30247) * $signed(input_fmap_101[7:0]) +
	( 16'sd 29873) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19239) * $signed(input_fmap_103[7:0]) +
	( 10'sd 466) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27878) * $signed(input_fmap_105[7:0]) +
	( 16'sd 27302) * $signed(input_fmap_106[7:0]) +
	( 16'sd 28887) * $signed(input_fmap_107[7:0]) +
	( 16'sd 23333) * $signed(input_fmap_108[7:0]) +
	( 15'sd 9743) * $signed(input_fmap_109[7:0]) +
	( 8'sd 77) * $signed(input_fmap_110[7:0]) +
	( 12'sd 1118) * $signed(input_fmap_111[7:0]) +
	( 14'sd 6050) * $signed(input_fmap_112[7:0]) +
	( 15'sd 10221) * $signed(input_fmap_113[7:0]) +
	( 14'sd 5763) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23168) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21837) * $signed(input_fmap_116[7:0]) +
	( 16'sd 27542) * $signed(input_fmap_117[7:0]) +
	( 16'sd 20441) * $signed(input_fmap_118[7:0]) +
	( 15'sd 12063) * $signed(input_fmap_119[7:0]) +
	( 16'sd 25122) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19011) * $signed(input_fmap_121[7:0]) +
	( 14'sd 5382) * $signed(input_fmap_122[7:0]) +
	( 15'sd 11474) * $signed(input_fmap_123[7:0]) +
	( 16'sd 32626) * $signed(input_fmap_124[7:0]) +
	( 15'sd 9519) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4274) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12029) * $signed(input_fmap_127[7:0]) +
	( 15'sd 11803) * $signed(input_fmap_128[7:0]) +
	( 15'sd 9008) * $signed(input_fmap_129[7:0]) +
	( 16'sd 24324) * $signed(input_fmap_130[7:0]) +
	( 16'sd 22849) * $signed(input_fmap_131[7:0]) +
	( 14'sd 7390) * $signed(input_fmap_132[7:0]) +
	( 16'sd 21013) * $signed(input_fmap_133[7:0]) +
	( 12'sd 1202) * $signed(input_fmap_134[7:0]) +
	( 16'sd 22705) * $signed(input_fmap_135[7:0]) +
	( 15'sd 14499) * $signed(input_fmap_136[7:0]) +
	( 14'sd 6732) * $signed(input_fmap_137[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_138[7:0]) +
	( 10'sd 457) * $signed(input_fmap_139[7:0]) +
	( 16'sd 26358) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29290) * $signed(input_fmap_141[7:0]) +
	( 16'sd 28764) * $signed(input_fmap_142[7:0]) +
	( 14'sd 7538) * $signed(input_fmap_143[7:0]) +
	( 16'sd 18024) * $signed(input_fmap_144[7:0]) +
	( 16'sd 20002) * $signed(input_fmap_145[7:0]) +
	( 13'sd 3284) * $signed(input_fmap_146[7:0]) +
	( 16'sd 28833) * $signed(input_fmap_147[7:0]) +
	( 16'sd 22703) * $signed(input_fmap_148[7:0]) +
	( 14'sd 4680) * $signed(input_fmap_149[7:0]) +
	( 16'sd 27830) * $signed(input_fmap_150[7:0]) +
	( 15'sd 12891) * $signed(input_fmap_151[7:0]) +
	( 15'sd 10262) * $signed(input_fmap_152[7:0]) +
	( 16'sd 17221) * $signed(input_fmap_153[7:0]) +
	( 15'sd 11494) * $signed(input_fmap_154[7:0]) +
	( 13'sd 3171) * $signed(input_fmap_155[7:0]) +
	( 15'sd 12903) * $signed(input_fmap_156[7:0]) +
	( 16'sd 19412) * $signed(input_fmap_157[7:0]) +
	( 14'sd 5456) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20736) * $signed(input_fmap_159[7:0]) +
	( 16'sd 20991) * $signed(input_fmap_160[7:0]) +
	( 16'sd 23721) * $signed(input_fmap_161[7:0]) +
	( 15'sd 8766) * $signed(input_fmap_162[7:0]) +
	( 15'sd 8778) * $signed(input_fmap_163[7:0]) +
	( 14'sd 6877) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23479) * $signed(input_fmap_165[7:0]) +
	( 16'sd 21835) * $signed(input_fmap_166[7:0]) +
	( 13'sd 2510) * $signed(input_fmap_167[7:0]) +
	( 16'sd 23974) * $signed(input_fmap_168[7:0]) +
	( 16'sd 16800) * $signed(input_fmap_169[7:0]) +
	( 16'sd 28681) * $signed(input_fmap_170[7:0]) +
	( 15'sd 10600) * $signed(input_fmap_171[7:0]) +
	( 16'sd 21899) * $signed(input_fmap_172[7:0]) +
	( 15'sd 11515) * $signed(input_fmap_173[7:0]) +
	( 14'sd 4130) * $signed(input_fmap_174[7:0]) +
	( 16'sd 22474) * $signed(input_fmap_175[7:0]) +
	( 15'sd 12899) * $signed(input_fmap_176[7:0]) +
	( 15'sd 14323) * $signed(input_fmap_177[7:0]) +
	( 16'sd 29463) * $signed(input_fmap_178[7:0]) +
	( 16'sd 29276) * $signed(input_fmap_179[7:0]) +
	( 15'sd 11116) * $signed(input_fmap_180[7:0]) +
	( 16'sd 19541) * $signed(input_fmap_181[7:0]) +
	( 14'sd 6513) * $signed(input_fmap_182[7:0]) +
	( 16'sd 31052) * $signed(input_fmap_183[7:0]) +
	( 14'sd 7323) * $signed(input_fmap_184[7:0]) +
	( 14'sd 5354) * $signed(input_fmap_185[7:0]) +
	( 13'sd 2612) * $signed(input_fmap_186[7:0]) +
	( 14'sd 4318) * $signed(input_fmap_187[7:0]) +
	( 16'sd 32565) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17757) * $signed(input_fmap_189[7:0]) +
	( 14'sd 6886) * $signed(input_fmap_190[7:0]) +
	( 14'sd 5477) * $signed(input_fmap_191[7:0]) +
	( 15'sd 11232) * $signed(input_fmap_192[7:0]) +
	( 16'sd 31887) * $signed(input_fmap_193[7:0]) +
	( 16'sd 28829) * $signed(input_fmap_194[7:0]) +
	( 16'sd 24889) * $signed(input_fmap_195[7:0]) +
	( 15'sd 8755) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25468) * $signed(input_fmap_197[7:0]) +
	( 15'sd 10128) * $signed(input_fmap_198[7:0]) +
	( 14'sd 5498) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13706) * $signed(input_fmap_200[7:0]) +
	( 16'sd 20651) * $signed(input_fmap_201[7:0]) +
	( 16'sd 24639) * $signed(input_fmap_202[7:0]) +
	( 10'sd 448) * $signed(input_fmap_203[7:0]) +
	( 16'sd 19562) * $signed(input_fmap_204[7:0]) +
	( 15'sd 15864) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21789) * $signed(input_fmap_206[7:0]) +
	( 15'sd 13179) * $signed(input_fmap_207[7:0]) +
	( 16'sd 21341) * $signed(input_fmap_208[7:0]) +
	( 16'sd 26428) * $signed(input_fmap_209[7:0]) +
	( 12'sd 1979) * $signed(input_fmap_210[7:0]) +
	( 15'sd 16025) * $signed(input_fmap_211[7:0]) +
	( 16'sd 19571) * $signed(input_fmap_212[7:0]) +
	( 15'sd 13304) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15705) * $signed(input_fmap_214[7:0]) +
	( 10'sd 434) * $signed(input_fmap_215[7:0]) +
	( 15'sd 12429) * $signed(input_fmap_216[7:0]) +
	( 15'sd 10249) * $signed(input_fmap_217[7:0]) +
	( 16'sd 29421) * $signed(input_fmap_218[7:0]) +
	( 16'sd 28464) * $signed(input_fmap_219[7:0]) +
	( 16'sd 24754) * $signed(input_fmap_220[7:0]) +
	( 16'sd 28839) * $signed(input_fmap_221[7:0]) +
	( 11'sd 974) * $signed(input_fmap_222[7:0]) +
	( 14'sd 5242) * $signed(input_fmap_223[7:0]) +
	( 15'sd 14970) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2106) * $signed(input_fmap_225[7:0]) +
	( 15'sd 10481) * $signed(input_fmap_226[7:0]) +
	( 15'sd 13761) * $signed(input_fmap_227[7:0]) +
	( 16'sd 24313) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20749) * $signed(input_fmap_229[7:0]) +
	( 16'sd 31333) * $signed(input_fmap_230[7:0]) +
	( 12'sd 1110) * $signed(input_fmap_231[7:0]) +
	( 12'sd 1502) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21011) * $signed(input_fmap_233[7:0]) +
	( 15'sd 15746) * $signed(input_fmap_234[7:0]) +
	( 14'sd 8057) * $signed(input_fmap_235[7:0]) +
	( 13'sd 3132) * $signed(input_fmap_236[7:0]) +
	( 16'sd 27893) * $signed(input_fmap_237[7:0]) +
	( 13'sd 2448) * $signed(input_fmap_238[7:0]) +
	( 16'sd 16552) * $signed(input_fmap_239[7:0]) +
	( 15'sd 8378) * $signed(input_fmap_240[7:0]) +
	( 15'sd 14308) * $signed(input_fmap_241[7:0]) +
	( 12'sd 1724) * $signed(input_fmap_242[7:0]) +
	( 15'sd 8648) * $signed(input_fmap_243[7:0]) +
	( 16'sd 28592) * $signed(input_fmap_244[7:0]) +
	( 16'sd 30719) * $signed(input_fmap_245[7:0]) +
	( 16'sd 28267) * $signed(input_fmap_246[7:0]) +
	( 16'sd 21130) * $signed(input_fmap_247[7:0]) +
	( 16'sd 28659) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4971) * $signed(input_fmap_249[7:0]) +
	( 15'sd 13489) * $signed(input_fmap_250[7:0]) +
	( 16'sd 23354) * $signed(input_fmap_251[7:0]) +
	( 14'sd 5307) * $signed(input_fmap_252[7:0]) +
	( 16'sd 28666) * $signed(input_fmap_253[7:0]) +
	( 13'sd 4000) * $signed(input_fmap_254[7:0]) +
	( 16'sd 27496) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_248;
assign conv_mac_248 = 
	( 16'sd 19460) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32698) * $signed(input_fmap_1[7:0]) +
	( 16'sd 21661) * $signed(input_fmap_2[7:0]) +
	( 16'sd 29840) * $signed(input_fmap_3[7:0]) +
	( 14'sd 7331) * $signed(input_fmap_4[7:0]) +
	( 16'sd 27058) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10493) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29461) * $signed(input_fmap_7[7:0]) +
	( 15'sd 12444) * $signed(input_fmap_8[7:0]) +
	( 16'sd 26207) * $signed(input_fmap_9[7:0]) +
	( 14'sd 7759) * $signed(input_fmap_10[7:0]) +
	( 15'sd 10644) * $signed(input_fmap_11[7:0]) +
	( 16'sd 22304) * $signed(input_fmap_12[7:0]) +
	( 16'sd 25562) * $signed(input_fmap_13[7:0]) +
	( 14'sd 5045) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14577) * $signed(input_fmap_15[7:0]) +
	( 15'sd 8956) * $signed(input_fmap_16[7:0]) +
	( 14'sd 6201) * $signed(input_fmap_17[7:0]) +
	( 16'sd 19313) * $signed(input_fmap_18[7:0]) +
	( 13'sd 2240) * $signed(input_fmap_19[7:0]) +
	( 15'sd 12245) * $signed(input_fmap_20[7:0]) +
	( 16'sd 18766) * $signed(input_fmap_21[7:0]) +
	( 14'sd 7884) * $signed(input_fmap_22[7:0]) +
	( 16'sd 30853) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27151) * $signed(input_fmap_24[7:0]) +
	( 15'sd 15450) * $signed(input_fmap_25[7:0]) +
	( 16'sd 21132) * $signed(input_fmap_26[7:0]) +
	( 13'sd 3254) * $signed(input_fmap_27[7:0]) +
	( 15'sd 11668) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18348) * $signed(input_fmap_29[7:0]) +
	( 15'sd 10933) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5024) * $signed(input_fmap_31[7:0]) +
	( 15'sd 9590) * $signed(input_fmap_32[7:0]) +
	( 16'sd 28132) * $signed(input_fmap_33[7:0]) +
	( 14'sd 6642) * $signed(input_fmap_34[7:0]) +
	( 16'sd 26080) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20248) * $signed(input_fmap_36[7:0]) +
	( 14'sd 6868) * $signed(input_fmap_37[7:0]) +
	( 10'sd 495) * $signed(input_fmap_38[7:0]) +
	( 14'sd 7335) * $signed(input_fmap_39[7:0]) +
	( 16'sd 20274) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28012) * $signed(input_fmap_41[7:0]) +
	( 12'sd 1841) * $signed(input_fmap_42[7:0]) +
	( 16'sd 23551) * $signed(input_fmap_43[7:0]) +
	( 16'sd 19956) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23744) * $signed(input_fmap_45[7:0]) +
	( 13'sd 2600) * $signed(input_fmap_46[7:0]) +
	( 16'sd 16753) * $signed(input_fmap_47[7:0]) +
	( 16'sd 25682) * $signed(input_fmap_48[7:0]) +
	( 14'sd 6870) * $signed(input_fmap_49[7:0]) +
	( 16'sd 19284) * $signed(input_fmap_50[7:0]) +
	( 16'sd 30852) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12362) * $signed(input_fmap_52[7:0]) +
	( 16'sd 17697) * $signed(input_fmap_53[7:0]) +
	( 14'sd 4952) * $signed(input_fmap_54[7:0]) +
	( 16'sd 27778) * $signed(input_fmap_55[7:0]) +
	( 16'sd 26915) * $signed(input_fmap_56[7:0]) +
	( 15'sd 8526) * $signed(input_fmap_57[7:0]) +
	( 16'sd 16656) * $signed(input_fmap_58[7:0]) +
	( 15'sd 11377) * $signed(input_fmap_59[7:0]) +
	( 11'sd 779) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27842) * $signed(input_fmap_61[7:0]) +
	( 13'sd 3457) * $signed(input_fmap_62[7:0]) +
	( 16'sd 18199) * $signed(input_fmap_63[7:0]) +
	( 16'sd 27280) * $signed(input_fmap_64[7:0]) +
	( 16'sd 20718) * $signed(input_fmap_65[7:0]) +
	( 15'sd 9839) * $signed(input_fmap_66[7:0]) +
	( 16'sd 25446) * $signed(input_fmap_67[7:0]) +
	( 16'sd 24017) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26456) * $signed(input_fmap_69[7:0]) +
	( 16'sd 27535) * $signed(input_fmap_70[7:0]) +
	( 16'sd 20708) * $signed(input_fmap_71[7:0]) +
	( 16'sd 28598) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29368) * $signed(input_fmap_73[7:0]) +
	( 16'sd 16670) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7845) * $signed(input_fmap_75[7:0]) +
	( 16'sd 17699) * $signed(input_fmap_76[7:0]) +
	( 15'sd 11754) * $signed(input_fmap_77[7:0]) +
	( 14'sd 4642) * $signed(input_fmap_78[7:0]) +
	( 15'sd 14474) * $signed(input_fmap_79[7:0]) +
	( 16'sd 30495) * $signed(input_fmap_80[7:0]) +
	( 14'sd 6507) * $signed(input_fmap_81[7:0]) +
	( 10'sd 334) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18773) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_84[7:0]) +
	( 15'sd 16357) * $signed(input_fmap_85[7:0]) +
	( 16'sd 22937) * $signed(input_fmap_86[7:0]) +
	( 16'sd 29003) * $signed(input_fmap_87[7:0]) +
	( 14'sd 6029) * $signed(input_fmap_88[7:0]) +
	( 16'sd 18047) * $signed(input_fmap_89[7:0]) +
	( 16'sd 28197) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27500) * $signed(input_fmap_91[7:0]) +
	( 16'sd 16524) * $signed(input_fmap_92[7:0]) +
	( 12'sd 1750) * $signed(input_fmap_93[7:0]) +
	( 16'sd 21285) * $signed(input_fmap_94[7:0]) +
	( 14'sd 7867) * $signed(input_fmap_95[7:0]) +
	( 12'sd 1519) * $signed(input_fmap_96[7:0]) +
	( 16'sd 27485) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22693) * $signed(input_fmap_98[7:0]) +
	( 16'sd 32195) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4164) * $signed(input_fmap_100[7:0]) +
	( 16'sd 28133) * $signed(input_fmap_101[7:0]) +
	( 16'sd 32435) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11817) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_104[7:0]) +
	( 16'sd 21116) * $signed(input_fmap_105[7:0]) +
	( 15'sd 9659) * $signed(input_fmap_106[7:0]) +
	( 15'sd 11858) * $signed(input_fmap_107[7:0]) +
	( 14'sd 4639) * $signed(input_fmap_108[7:0]) +
	( 16'sd 28900) * $signed(input_fmap_109[7:0]) +
	( 15'sd 13159) * $signed(input_fmap_110[7:0]) +
	( 16'sd 19130) * $signed(input_fmap_111[7:0]) +
	( 15'sd 13549) * $signed(input_fmap_112[7:0]) +
	( 15'sd 12672) * $signed(input_fmap_113[7:0]) +
	( 15'sd 11949) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2687) * $signed(input_fmap_115[7:0]) +
	( 16'sd 19912) * $signed(input_fmap_116[7:0]) +
	( 9'sd 241) * $signed(input_fmap_117[7:0]) +
	( 15'sd 14943) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17923) * $signed(input_fmap_119[7:0]) +
	( 16'sd 21865) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14701) * $signed(input_fmap_121[7:0]) +
	( 14'sd 4462) * $signed(input_fmap_122[7:0]) +
	( 14'sd 6765) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17295) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2646) * $signed(input_fmap_125[7:0]) +
	( 16'sd 18847) * $signed(input_fmap_126[7:0]) +
	( 15'sd 12168) * $signed(input_fmap_127[7:0]) +
	( 15'sd 10035) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31137) * $signed(input_fmap_129[7:0]) +
	( 15'sd 16336) * $signed(input_fmap_130[7:0]) +
	( 12'sd 1777) * $signed(input_fmap_131[7:0]) +
	( 15'sd 8903) * $signed(input_fmap_132[7:0]) +
	( 16'sd 19314) * $signed(input_fmap_133[7:0]) +
	( 15'sd 9047) * $signed(input_fmap_134[7:0]) +
	( 16'sd 25679) * $signed(input_fmap_135[7:0]) +
	( 13'sd 3221) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24737) * $signed(input_fmap_137[7:0]) +
	( 14'sd 5814) * $signed(input_fmap_138[7:0]) +
	( 15'sd 16269) * $signed(input_fmap_139[7:0]) +
	( 12'sd 1569) * $signed(input_fmap_140[7:0]) +
	( 15'sd 10905) * $signed(input_fmap_141[7:0]) +
	( 16'sd 23548) * $signed(input_fmap_142[7:0]) +
	( 16'sd 31729) * $signed(input_fmap_143[7:0]) +
	( 11'sd 902) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17526) * $signed(input_fmap_145[7:0]) +
	( 16'sd 25514) * $signed(input_fmap_146[7:0]) +
	( 15'sd 11268) * $signed(input_fmap_147[7:0]) +
	( 16'sd 31013) * $signed(input_fmap_148[7:0]) +
	( 14'sd 6720) * $signed(input_fmap_149[7:0]) +
	( 16'sd 26338) * $signed(input_fmap_150[7:0]) +
	( 16'sd 30810) * $signed(input_fmap_151[7:0]) +
	( 14'sd 7977) * $signed(input_fmap_152[7:0]) +
	( 16'sd 30686) * $signed(input_fmap_153[7:0]) +
	( 15'sd 12343) * $signed(input_fmap_154[7:0]) +
	( 15'sd 14250) * $signed(input_fmap_155[7:0]) +
	( 15'sd 8884) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30554) * $signed(input_fmap_157[7:0]) +
	( 16'sd 27981) * $signed(input_fmap_158[7:0]) +
	( 14'sd 4255) * $signed(input_fmap_159[7:0]) +
	( 15'sd 10502) * $signed(input_fmap_160[7:0]) +
	( 16'sd 22020) * $signed(input_fmap_161[7:0]) +
	( 16'sd 19149) * $signed(input_fmap_162[7:0]) +
	( 13'sd 3770) * $signed(input_fmap_163[7:0]) +
	( 14'sd 4818) * $signed(input_fmap_164[7:0]) +
	( 16'sd 31585) * $signed(input_fmap_165[7:0]) +
	( 13'sd 2455) * $signed(input_fmap_166[7:0]) +
	( 12'sd 1954) * $signed(input_fmap_167[7:0]) +
	( 15'sd 12819) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11528) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9575) * $signed(input_fmap_170[7:0]) +
	( 16'sd 21492) * $signed(input_fmap_171[7:0]) +
	( 16'sd 17825) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23357) * $signed(input_fmap_173[7:0]) +
	( 10'sd 480) * $signed(input_fmap_174[7:0]) +
	( 15'sd 14922) * $signed(input_fmap_175[7:0]) +
	( 15'sd 11011) * $signed(input_fmap_176[7:0]) +
	( 14'sd 8024) * $signed(input_fmap_177[7:0]) +
	( 11'sd 945) * $signed(input_fmap_178[7:0]) +
	( 16'sd 23146) * $signed(input_fmap_179[7:0]) +
	( 16'sd 30141) * $signed(input_fmap_180[7:0]) +
	( 16'sd 31270) * $signed(input_fmap_181[7:0]) +
	( 16'sd 30711) * $signed(input_fmap_182[7:0]) +
	( 12'sd 1047) * $signed(input_fmap_183[7:0]) +
	( 16'sd 27100) * $signed(input_fmap_184[7:0]) +
	( 15'sd 16015) * $signed(input_fmap_185[7:0]) +
	( 16'sd 21531) * $signed(input_fmap_186[7:0]) +
	( 16'sd 22086) * $signed(input_fmap_187[7:0]) +
	( 16'sd 19982) * $signed(input_fmap_188[7:0]) +
	( 16'sd 28437) * $signed(input_fmap_189[7:0]) +
	( 15'sd 12543) * $signed(input_fmap_190[7:0]) +
	( 14'sd 6331) * $signed(input_fmap_191[7:0]) +
	( 16'sd 30804) * $signed(input_fmap_192[7:0]) +
	( 15'sd 14781) * $signed(input_fmap_193[7:0]) +
	( 12'sd 1531) * $signed(input_fmap_194[7:0]) +
	( 14'sd 6376) * $signed(input_fmap_195[7:0]) +
	( 15'sd 14384) * $signed(input_fmap_196[7:0]) +
	( 15'sd 14089) * $signed(input_fmap_197[7:0]) +
	( 15'sd 13829) * $signed(input_fmap_198[7:0]) +
	( 15'sd 10222) * $signed(input_fmap_199[7:0]) +
	( 13'sd 3127) * $signed(input_fmap_200[7:0]) +
	( 16'sd 18435) * $signed(input_fmap_201[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_202[7:0]) +
	( 16'sd 30467) * $signed(input_fmap_203[7:0]) +
	( 16'sd 17027) * $signed(input_fmap_204[7:0]) +
	( 11'sd 668) * $signed(input_fmap_205[7:0]) +
	( 14'sd 7244) * $signed(input_fmap_206[7:0]) +
	( 16'sd 20707) * $signed(input_fmap_207[7:0]) +
	( 15'sd 13706) * $signed(input_fmap_208[7:0]) +
	( 16'sd 25135) * $signed(input_fmap_209[7:0]) +
	( 15'sd 15630) * $signed(input_fmap_210[7:0]) +
	( 16'sd 26455) * $signed(input_fmap_211[7:0]) +
	( 14'sd 4721) * $signed(input_fmap_212[7:0]) +
	( 13'sd 2601) * $signed(input_fmap_213[7:0]) +
	( 15'sd 9461) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11382) * $signed(input_fmap_215[7:0]) +
	( 12'sd 1643) * $signed(input_fmap_216[7:0]) +
	( 15'sd 12521) * $signed(input_fmap_217[7:0]) +
	( 13'sd 3538) * $signed(input_fmap_218[7:0]) +
	( 14'sd 5291) * $signed(input_fmap_219[7:0]) +
	( 16'sd 17058) * $signed(input_fmap_220[7:0]) +
	( 15'sd 10312) * $signed(input_fmap_221[7:0]) +
	( 16'sd 23621) * $signed(input_fmap_222[7:0]) +
	( 16'sd 21896) * $signed(input_fmap_223[7:0]) +
	( 16'sd 20852) * $signed(input_fmap_224[7:0]) +
	( 13'sd 2065) * $signed(input_fmap_225[7:0]) +
	( 12'sd 1464) * $signed(input_fmap_226[7:0]) +
	( 16'sd 30877) * $signed(input_fmap_227[7:0]) +
	( 15'sd 16247) * $signed(input_fmap_228[7:0]) +
	( 16'sd 18664) * $signed(input_fmap_229[7:0]) +
	( 16'sd 28846) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25770) * $signed(input_fmap_231[7:0]) +
	( 15'sd 8726) * $signed(input_fmap_232[7:0]) +
	( 10'sd 311) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4441) * $signed(input_fmap_234[7:0]) +
	( 14'sd 7518) * $signed(input_fmap_235[7:0]) +
	( 14'sd 7050) * $signed(input_fmap_236[7:0]) +
	( 16'sd 19836) * $signed(input_fmap_237[7:0]) +
	( 15'sd 15909) * $signed(input_fmap_238[7:0]) +
	( 16'sd 18570) * $signed(input_fmap_239[7:0]) +
	( 16'sd 26996) * $signed(input_fmap_240[7:0]) +
	( 15'sd 12216) * $signed(input_fmap_241[7:0]) +
	( 14'sd 5376) * $signed(input_fmap_242[7:0]) +
	( 16'sd 21369) * $signed(input_fmap_243[7:0]) +
	( 16'sd 29591) * $signed(input_fmap_244[7:0]) +
	( 16'sd 19122) * $signed(input_fmap_245[7:0]) +
	( 15'sd 14109) * $signed(input_fmap_246[7:0]) +
	( 16'sd 18038) * $signed(input_fmap_247[7:0]) +
	( 15'sd 15020) * $signed(input_fmap_248[7:0]) +
	( 16'sd 20571) * $signed(input_fmap_249[7:0]) +
	( 16'sd 31053) * $signed(input_fmap_250[7:0]) +
	( 15'sd 14244) * $signed(input_fmap_251[7:0]) +
	( 16'sd 18808) * $signed(input_fmap_252[7:0]) +
	( 16'sd 26100) * $signed(input_fmap_253[7:0]) +
	( 12'sd 1250) * $signed(input_fmap_254[7:0]) +
	( 16'sd 32498) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_249;
assign conv_mac_249 = 
	( 16'sd 28742) * $signed(input_fmap_0[7:0]) +
	( 16'sd 22486) * $signed(input_fmap_1[7:0]) +
	( 16'sd 30898) * $signed(input_fmap_2[7:0]) +
	( 14'sd 5836) * $signed(input_fmap_3[7:0]) +
	( 9'sd 200) * $signed(input_fmap_4[7:0]) +
	( 15'sd 14042) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4966) * $signed(input_fmap_6[7:0]) +
	( 16'sd 16612) * $signed(input_fmap_7[7:0]) +
	( 16'sd 16986) * $signed(input_fmap_8[7:0]) +
	( 14'sd 5952) * $signed(input_fmap_9[7:0]) +
	( 12'sd 1979) * $signed(input_fmap_10[7:0]) +
	( 15'sd 14094) * $signed(input_fmap_11[7:0]) +
	( 13'sd 3782) * $signed(input_fmap_12[7:0]) +
	( 15'sd 9914) * $signed(input_fmap_13[7:0]) +
	( 15'sd 10010) * $signed(input_fmap_14[7:0]) +
	( 15'sd 14527) * $signed(input_fmap_15[7:0]) +
	( 13'sd 2360) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26217) * $signed(input_fmap_17[7:0]) +
	( 14'sd 4778) * $signed(input_fmap_18[7:0]) +
	( 16'sd 17463) * $signed(input_fmap_19[7:0]) +
	( 16'sd 18101) * $signed(input_fmap_20[7:0]) +
	( 15'sd 16161) * $signed(input_fmap_21[7:0]) +
	( 16'sd 21830) * $signed(input_fmap_22[7:0]) +
	( 16'sd 29105) * $signed(input_fmap_23[7:0]) +
	( 14'sd 7030) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20163) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22254) * $signed(input_fmap_26[7:0]) +
	( 15'sd 13517) * $signed(input_fmap_27[7:0]) +
	( 12'sd 1981) * $signed(input_fmap_28[7:0]) +
	( 16'sd 23270) * $signed(input_fmap_29[7:0]) +
	( 14'sd 5157) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1681) * $signed(input_fmap_31[7:0]) +
	( 16'sd 16478) * $signed(input_fmap_32[7:0]) +
	( 15'sd 8948) * $signed(input_fmap_33[7:0]) +
	( 16'sd 24142) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11260) * $signed(input_fmap_35[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_36[7:0]) +
	( 15'sd 13283) * $signed(input_fmap_37[7:0]) +
	( 14'sd 4282) * $signed(input_fmap_38[7:0]) +
	( 16'sd 20556) * $signed(input_fmap_39[7:0]) +
	( 16'sd 18900) * $signed(input_fmap_40[7:0]) +
	( 16'sd 17007) * $signed(input_fmap_41[7:0]) +
	( 15'sd 9227) * $signed(input_fmap_42[7:0]) +
	( 16'sd 20357) * $signed(input_fmap_43[7:0]) +
	( 16'sd 22577) * $signed(input_fmap_44[7:0]) +
	( 9'sd 202) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22499) * $signed(input_fmap_46[7:0]) +
	( 14'sd 5014) * $signed(input_fmap_47[7:0]) +
	( 11'sd 617) * $signed(input_fmap_48[7:0]) +
	( 16'sd 18898) * $signed(input_fmap_49[7:0]) +
	( 15'sd 11161) * $signed(input_fmap_50[7:0]) +
	( 8'sd 126) * $signed(input_fmap_51[7:0]) +
	( 15'sd 15128) * $signed(input_fmap_52[7:0]) +
	( 16'sd 16573) * $signed(input_fmap_53[7:0]) +
	( 15'sd 9785) * $signed(input_fmap_54[7:0]) +
	( 15'sd 12259) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20373) * $signed(input_fmap_56[7:0]) +
	( 15'sd 13014) * $signed(input_fmap_57[7:0]) +
	( 16'sd 19114) * $signed(input_fmap_58[7:0]) +
	( 16'sd 31762) * $signed(input_fmap_59[7:0]) +
	( 16'sd 19518) * $signed(input_fmap_60[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8878) * $signed(input_fmap_62[7:0]) +
	( 15'sd 13232) * $signed(input_fmap_63[7:0]) +
	( 16'sd 24654) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4452) * $signed(input_fmap_65[7:0]) +
	( 16'sd 23290) * $signed(input_fmap_66[7:0]) +
	( 16'sd 31886) * $signed(input_fmap_67[7:0]) +
	( 14'sd 7841) * $signed(input_fmap_68[7:0]) +
	( 16'sd 26152) * $signed(input_fmap_69[7:0]) +
	( 15'sd 14375) * $signed(input_fmap_70[7:0]) +
	( 15'sd 14254) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18133) * $signed(input_fmap_72[7:0]) +
	( 16'sd 20393) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9401) * $signed(input_fmap_74[7:0]) +
	( 16'sd 29927) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29218) * $signed(input_fmap_76[7:0]) +
	( 13'sd 2328) * $signed(input_fmap_77[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_78[7:0]) +
	( 16'sd 31960) * $signed(input_fmap_79[7:0]) +
	( 16'sd 16684) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13116) * $signed(input_fmap_81[7:0]) +
	( 15'sd 9231) * $signed(input_fmap_82[7:0]) +
	( 16'sd 17485) * $signed(input_fmap_83[7:0]) +
	( 12'sd 1373) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2193) * $signed(input_fmap_85[7:0]) +
	( 15'sd 15329) * $signed(input_fmap_86[7:0]) +
	( 16'sd 25361) * $signed(input_fmap_87[7:0]) +
	( 12'sd 1272) * $signed(input_fmap_88[7:0]) +
	( 16'sd 31337) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29031) * $signed(input_fmap_90[7:0]) +
	( 16'sd 28043) * $signed(input_fmap_91[7:0]) +
	( 16'sd 24664) * $signed(input_fmap_92[7:0]) +
	( 16'sd 22974) * $signed(input_fmap_93[7:0]) +
	( 14'sd 5467) * $signed(input_fmap_94[7:0]) +
	( 15'sd 8883) * $signed(input_fmap_95[7:0]) +
	( 16'sd 25257) * $signed(input_fmap_96[7:0]) +
	( 14'sd 7059) * $signed(input_fmap_97[7:0]) +
	( 12'sd 1784) * $signed(input_fmap_98[7:0]) +
	( 16'sd 27176) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15600) * $signed(input_fmap_100[7:0]) +
	( 16'sd 19963) * $signed(input_fmap_101[7:0]) +
	( 16'sd 28417) * $signed(input_fmap_102[7:0]) +
	( 16'sd 16886) * $signed(input_fmap_103[7:0]) +
	( 16'sd 21514) * $signed(input_fmap_104[7:0]) +
	( 15'sd 10560) * $signed(input_fmap_105[7:0]) +
	( 15'sd 15389) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_107[7:0]) +
	( 16'sd 30627) * $signed(input_fmap_108[7:0]) +
	( 15'sd 11363) * $signed(input_fmap_109[7:0]) +
	( 16'sd 22157) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22760) * $signed(input_fmap_111[7:0]) +
	( 16'sd 24386) * $signed(input_fmap_112[7:0]) +
	( 15'sd 8192) * $signed(input_fmap_113[7:0]) +
	( 14'sd 6084) * $signed(input_fmap_114[7:0]) +
	( 14'sd 5578) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29530) * $signed(input_fmap_116[7:0]) +
	( 16'sd 24804) * $signed(input_fmap_117[7:0]) +
	( 14'sd 7956) * $signed(input_fmap_118[7:0]) +
	( 16'sd 31848) * $signed(input_fmap_119[7:0]) +
	( 16'sd 22072) * $signed(input_fmap_120[7:0]) +
	( 16'sd 22229) * $signed(input_fmap_121[7:0]) +
	( 16'sd 27984) * $signed(input_fmap_122[7:0]) +
	( 15'sd 15874) * $signed(input_fmap_123[7:0]) +
	( 16'sd 17688) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1624) * $signed(input_fmap_125[7:0]) +
	( 16'sd 30136) * $signed(input_fmap_126[7:0]) +
	( 14'sd 6974) * $signed(input_fmap_127[7:0]) +
	( 15'sd 9257) * $signed(input_fmap_128[7:0]) +
	( 16'sd 17342) * $signed(input_fmap_129[7:0]) +
	( 15'sd 12044) * $signed(input_fmap_130[7:0]) +
	( 16'sd 17279) * $signed(input_fmap_131[7:0]) +
	( 15'sd 14046) * $signed(input_fmap_132[7:0]) +
	( 16'sd 22816) * $signed(input_fmap_133[7:0]) +
	( 16'sd 19205) * $signed(input_fmap_134[7:0]) +
	( 16'sd 32403) * $signed(input_fmap_135[7:0]) +
	( 13'sd 2254) * $signed(input_fmap_136[7:0]) +
	( 15'sd 12666) * $signed(input_fmap_137[7:0]) +
	( 11'sd 752) * $signed(input_fmap_138[7:0]) +
	( 15'sd 11633) * $signed(input_fmap_139[7:0]) +
	( 16'sd 31031) * $signed(input_fmap_140[7:0]) +
	( 16'sd 29888) * $signed(input_fmap_141[7:0]) +
	( 15'sd 12066) * $signed(input_fmap_142[7:0]) +
	( 16'sd 23391) * $signed(input_fmap_143[7:0]) +
	( 16'sd 30535) * $signed(input_fmap_144[7:0]) +
	( 16'sd 28928) * $signed(input_fmap_145[7:0]) +
	( 16'sd 21046) * $signed(input_fmap_146[7:0]) +
	( 16'sd 19955) * $signed(input_fmap_147[7:0]) +
	( 16'sd 29129) * $signed(input_fmap_148[7:0]) +
	( 15'sd 11430) * $signed(input_fmap_149[7:0]) +
	( 15'sd 14884) * $signed(input_fmap_150[7:0]) +
	( 16'sd 23386) * $signed(input_fmap_151[7:0]) +
	( 16'sd 18573) * $signed(input_fmap_152[7:0]) +
	( 14'sd 4983) * $signed(input_fmap_153[7:0]) +
	( 16'sd 28295) * $signed(input_fmap_154[7:0]) +
	( 16'sd 30646) * $signed(input_fmap_155[7:0]) +
	( 11'sd 911) * $signed(input_fmap_156[7:0]) +
	( 16'sd 23111) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20197) * $signed(input_fmap_158[7:0]) +
	( 16'sd 20220) * $signed(input_fmap_159[7:0]) +
	( 16'sd 29745) * $signed(input_fmap_160[7:0]) +
	( 16'sd 19918) * $signed(input_fmap_161[7:0]) +
	( 16'sd 18616) * $signed(input_fmap_162[7:0]) +
	( 16'sd 19118) * $signed(input_fmap_163[7:0]) +
	( 16'sd 18156) * $signed(input_fmap_164[7:0]) +
	( 16'sd 23946) * $signed(input_fmap_165[7:0]) +
	( 15'sd 16125) * $signed(input_fmap_166[7:0]) +
	( 15'sd 9691) * $signed(input_fmap_167[7:0]) +
	( 15'sd 8938) * $signed(input_fmap_168[7:0]) +
	( 16'sd 28663) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5908) * $signed(input_fmap_170[7:0]) +
	( 16'sd 18270) * $signed(input_fmap_171[7:0]) +
	( 16'sd 27877) * $signed(input_fmap_172[7:0]) +
	( 16'sd 32237) * $signed(input_fmap_173[7:0]) +
	( 16'sd 31826) * $signed(input_fmap_174[7:0]) +
	( 16'sd 25768) * $signed(input_fmap_175[7:0]) +
	( 14'sd 7867) * $signed(input_fmap_176[7:0]) +
	( 16'sd 18196) * $signed(input_fmap_177[7:0]) +
	( 16'sd 32068) * $signed(input_fmap_178[7:0]) +
	( 16'sd 28278) * $signed(input_fmap_179[7:0]) +
	( 15'sd 12960) * $signed(input_fmap_180[7:0]) +
	( 16'sd 28063) * $signed(input_fmap_181[7:0]) +
	( 16'sd 18418) * $signed(input_fmap_182[7:0]) +
	( 16'sd 28094) * $signed(input_fmap_183[7:0]) +
	( 10'sd 260) * $signed(input_fmap_184[7:0]) +
	( 15'sd 13631) * $signed(input_fmap_185[7:0]) +
	( 16'sd 23019) * $signed(input_fmap_186[7:0]) +
	( 16'sd 25459) * $signed(input_fmap_187[7:0]) +
	( 16'sd 31389) * $signed(input_fmap_188[7:0]) +
	( 10'sd 423) * $signed(input_fmap_189[7:0]) +
	( 14'sd 4847) * $signed(input_fmap_190[7:0]) +
	( 16'sd 28745) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15419) * $signed(input_fmap_192[7:0]) +
	( 14'sd 4501) * $signed(input_fmap_193[7:0]) +
	( 14'sd 5574) * $signed(input_fmap_194[7:0]) +
	( 16'sd 26475) * $signed(input_fmap_195[7:0]) +
	( 16'sd 31846) * $signed(input_fmap_196[7:0]) +
	( 13'sd 3091) * $signed(input_fmap_197[7:0]) +
	( 13'sd 2457) * $signed(input_fmap_198[7:0]) +
	( 16'sd 22610) * $signed(input_fmap_199[7:0]) +
	( 15'sd 13399) * $signed(input_fmap_200[7:0]) +
	( 16'sd 26852) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2844) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2380) * $signed(input_fmap_203[7:0]) +
	( 12'sd 1682) * $signed(input_fmap_204[7:0]) +
	( 13'sd 3774) * $signed(input_fmap_205[7:0]) +
	( 15'sd 14058) * $signed(input_fmap_206[7:0]) +
	( 16'sd 19116) * $signed(input_fmap_207[7:0]) +
	( 16'sd 16939) * $signed(input_fmap_208[7:0]) +
	( 15'sd 13689) * $signed(input_fmap_209[7:0]) +
	( 13'sd 2584) * $signed(input_fmap_210[7:0]) +
	( 16'sd 20082) * $signed(input_fmap_211[7:0]) +
	( 15'sd 11034) * $signed(input_fmap_212[7:0]) +
	( 9'sd 213) * $signed(input_fmap_213[7:0]) +
	( 15'sd 15350) * $signed(input_fmap_214[7:0]) +
	( 16'sd 17472) * $signed(input_fmap_215[7:0]) +
	( 16'sd 24421) * $signed(input_fmap_216[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22161) * $signed(input_fmap_218[7:0]) +
	( 16'sd 30207) * $signed(input_fmap_219[7:0]) +
	( 16'sd 19873) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1223) * $signed(input_fmap_221[7:0]) +
	( 13'sd 3837) * $signed(input_fmap_222[7:0]) +
	( 13'sd 2336) * $signed(input_fmap_223[7:0]) +
	( 16'sd 32079) * $signed(input_fmap_224[7:0]) +
	( 16'sd 16696) * $signed(input_fmap_225[7:0]) +
	( 16'sd 27038) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27527) * $signed(input_fmap_227[7:0]) +
	( 16'sd 23342) * $signed(input_fmap_228[7:0]) +
	( 15'sd 16071) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29655) * $signed(input_fmap_230[7:0]) +
	( 16'sd 26351) * $signed(input_fmap_231[7:0]) +
	( 15'sd 12372) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3775) * $signed(input_fmap_233[7:0]) +
	( 14'sd 6294) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3599) * $signed(input_fmap_235[7:0]) +
	( 12'sd 1610) * $signed(input_fmap_236[7:0]) +
	( 15'sd 10122) * $signed(input_fmap_237[7:0]) +
	( 16'sd 30102) * $signed(input_fmap_238[7:0]) +
	( 16'sd 20455) * $signed(input_fmap_239[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_240[7:0]) +
	( 16'sd 18009) * $signed(input_fmap_241[7:0]) +
	( 16'sd 17563) * $signed(input_fmap_242[7:0]) +
	( 14'sd 7406) * $signed(input_fmap_243[7:0]) +
	( 15'sd 13872) * $signed(input_fmap_244[7:0]) +
	( 11'sd 545) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22826) * $signed(input_fmap_246[7:0]) +
	( 14'sd 4490) * $signed(input_fmap_247[7:0]) +
	( 16'sd 18134) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28650) * $signed(input_fmap_249[7:0]) +
	( 16'sd 31248) * $signed(input_fmap_250[7:0]) +
	( 14'sd 6743) * $signed(input_fmap_251[7:0]) +
	( 15'sd 13857) * $signed(input_fmap_252[7:0]) +
	( 16'sd 27794) * $signed(input_fmap_253[7:0]) +
	( 10'sd 451) * $signed(input_fmap_254[7:0]) +
	( 16'sd 16869) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_250;
assign conv_mac_250 = 
	( 14'sd 6715) * $signed(input_fmap_0[7:0]) +
	( 11'sd 948) * $signed(input_fmap_1[7:0]) +
	( 13'sd 2272) * $signed(input_fmap_2[7:0]) +
	( 11'sd 869) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5192) * $signed(input_fmap_4[7:0]) +
	( 16'sd 26626) * $signed(input_fmap_5[7:0]) +
	( 13'sd 3204) * $signed(input_fmap_6[7:0]) +
	( 15'sd 13119) * $signed(input_fmap_7[7:0]) +
	( 11'sd 692) * $signed(input_fmap_8[7:0]) +
	( 16'sd 16479) * $signed(input_fmap_9[7:0]) +
	( 16'sd 32761) * $signed(input_fmap_10[7:0]) +
	( 16'sd 17827) * $signed(input_fmap_11[7:0]) +
	( 10'sd 383) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1166) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27378) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29648) * $signed(input_fmap_15[7:0]) +
	( 16'sd 31509) * $signed(input_fmap_16[7:0]) +
	( 16'sd 26607) * $signed(input_fmap_17[7:0]) +
	( 16'sd 20354) * $signed(input_fmap_18[7:0]) +
	( 14'sd 4513) * $signed(input_fmap_19[7:0]) +
	( 16'sd 16911) * $signed(input_fmap_20[7:0]) +
	( 15'sd 11993) * $signed(input_fmap_21[7:0]) +
	( 16'sd 24905) * $signed(input_fmap_22[7:0]) +
	( 16'sd 17390) * $signed(input_fmap_23[7:0]) +
	( 15'sd 10205) * $signed(input_fmap_24[7:0]) +
	( 16'sd 24198) * $signed(input_fmap_25[7:0]) +
	( 15'sd 16137) * $signed(input_fmap_26[7:0]) +
	( 16'sd 29210) * $signed(input_fmap_27[7:0]) +
	( 15'sd 13032) * $signed(input_fmap_28[7:0]) +
	( 13'sd 3268) * $signed(input_fmap_29[7:0]) +
	( 16'sd 32636) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12126) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2586) * $signed(input_fmap_32[7:0]) +
	( 15'sd 16280) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11690) * $signed(input_fmap_34[7:0]) +
	( 15'sd 14782) * $signed(input_fmap_35[7:0]) +
	( 16'sd 30505) * $signed(input_fmap_36[7:0]) +
	( 13'sd 3160) * $signed(input_fmap_37[7:0]) +
	( 15'sd 15423) * $signed(input_fmap_38[7:0]) +
	( 16'sd 23397) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11849) * $signed(input_fmap_40[7:0]) +
	( 12'sd 1644) * $signed(input_fmap_41[7:0]) +
	( 16'sd 23101) * $signed(input_fmap_42[7:0]) +
	( 15'sd 15315) * $signed(input_fmap_43[7:0]) +
	( 15'sd 15025) * $signed(input_fmap_44[7:0]) +
	( 16'sd 22995) * $signed(input_fmap_45[7:0]) +
	( 15'sd 14789) * $signed(input_fmap_46[7:0]) +
	( 16'sd 28768) * $signed(input_fmap_47[7:0]) +
	( 16'sd 28240) * $signed(input_fmap_48[7:0]) +
	( 15'sd 15630) * $signed(input_fmap_49[7:0]) +
	( 15'sd 12009) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7580) * $signed(input_fmap_51[7:0]) +
	( 15'sd 12685) * $signed(input_fmap_52[7:0]) +
	( 15'sd 13932) * $signed(input_fmap_53[7:0]) +
	( 16'sd 25766) * $signed(input_fmap_54[7:0]) +
	( 16'sd 21241) * $signed(input_fmap_55[7:0]) +
	( 16'sd 32412) * $signed(input_fmap_56[7:0]) +
	( 15'sd 14918) * $signed(input_fmap_57[7:0]) +
	( 16'sd 29787) * $signed(input_fmap_58[7:0]) +
	( 16'sd 23073) * $signed(input_fmap_59[7:0]) +
	( 15'sd 11868) * $signed(input_fmap_60[7:0]) +
	( 16'sd 17715) * $signed(input_fmap_61[7:0]) +
	( 10'sd 406) * $signed(input_fmap_62[7:0]) +
	( 13'sd 4030) * $signed(input_fmap_63[7:0]) +
	( 14'sd 5680) * $signed(input_fmap_64[7:0]) +
	( 16'sd 30732) * $signed(input_fmap_65[7:0]) +
	( 15'sd 11473) * $signed(input_fmap_66[7:0]) +
	( 15'sd 14734) * $signed(input_fmap_67[7:0]) +
	( 16'sd 29724) * $signed(input_fmap_68[7:0]) +
	( 14'sd 5797) * $signed(input_fmap_69[7:0]) +
	( 14'sd 5350) * $signed(input_fmap_70[7:0]) +
	( 16'sd 30564) * $signed(input_fmap_71[7:0]) +
	( 16'sd 18269) * $signed(input_fmap_72[7:0]) +
	( 16'sd 24815) * $signed(input_fmap_73[7:0]) +
	( 15'sd 9342) * $signed(input_fmap_74[7:0]) +
	( 14'sd 6957) * $signed(input_fmap_75[7:0]) +
	( 15'sd 13838) * $signed(input_fmap_76[7:0]) +
	( 16'sd 25002) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9890) * $signed(input_fmap_78[7:0]) +
	( 13'sd 3237) * $signed(input_fmap_79[7:0]) +
	( 16'sd 20968) * $signed(input_fmap_80[7:0]) +
	( 15'sd 13875) * $signed(input_fmap_81[7:0]) +
	( 12'sd 1338) * $signed(input_fmap_82[7:0]) +
	( 15'sd 14542) * $signed(input_fmap_83[7:0]) +
	( 15'sd 11723) * $signed(input_fmap_84[7:0]) +
	( 13'sd 2650) * $signed(input_fmap_85[7:0]) +
	( 16'sd 28531) * $signed(input_fmap_86[7:0]) +
	( 16'sd 17422) * $signed(input_fmap_87[7:0]) +
	( 14'sd 7405) * $signed(input_fmap_88[7:0]) +
	( 13'sd 2338) * $signed(input_fmap_89[7:0]) +
	( 12'sd 2046) * $signed(input_fmap_90[7:0]) +
	( 16'sd 17936) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3215) * $signed(input_fmap_92[7:0]) +
	( 16'sd 32595) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12852) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30880) * $signed(input_fmap_95[7:0]) +
	( 16'sd 21509) * $signed(input_fmap_96[7:0]) +
	( 12'sd 1777) * $signed(input_fmap_97[7:0]) +
	( 16'sd 22280) * $signed(input_fmap_98[7:0]) +
	( 11'sd 855) * $signed(input_fmap_99[7:0]) +
	( 14'sd 4661) * $signed(input_fmap_100[7:0]) +
	( 15'sd 12053) * $signed(input_fmap_101[7:0]) +
	( 14'sd 4786) * $signed(input_fmap_102[7:0]) +
	( 15'sd 13299) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30028) * $signed(input_fmap_104[7:0]) +
	( 16'sd 30472) * $signed(input_fmap_105[7:0]) +
	( 16'sd 22694) * $signed(input_fmap_106[7:0]) +
	( 14'sd 4776) * $signed(input_fmap_107[7:0]) +
	( 15'sd 14073) * $signed(input_fmap_108[7:0]) +
	( 16'sd 26283) * $signed(input_fmap_109[7:0]) +
	( 13'sd 2567) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26309) * $signed(input_fmap_111[7:0]) +
	( 11'sd 789) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5841) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17540) * $signed(input_fmap_114[7:0]) +
	( 16'sd 31879) * $signed(input_fmap_115[7:0]) +
	( 15'sd 14468) * $signed(input_fmap_116[7:0]) +
	( 16'sd 32501) * $signed(input_fmap_117[7:0]) +
	( 14'sd 4098) * $signed(input_fmap_118[7:0]) +
	( 16'sd 22084) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11421) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14735) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15663) * $signed(input_fmap_122[7:0]) +
	( 16'sd 26901) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27819) * $signed(input_fmap_124[7:0]) +
	( 12'sd 1767) * $signed(input_fmap_125[7:0]) +
	( 15'sd 14374) * $signed(input_fmap_126[7:0]) +
	( 16'sd 22477) * $signed(input_fmap_127[7:0]) +
	( 15'sd 15024) * $signed(input_fmap_128[7:0]) +
	( 16'sd 28380) * $signed(input_fmap_129[7:0]) +
	( 16'sd 19993) * $signed(input_fmap_130[7:0]) +
	( 16'sd 26035) * $signed(input_fmap_131[7:0]) +
	( 14'sd 5226) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12473) * $signed(input_fmap_133[7:0]) +
	( 16'sd 26312) * $signed(input_fmap_134[7:0]) +
	( 16'sd 17932) * $signed(input_fmap_135[7:0]) +
	( 16'sd 16973) * $signed(input_fmap_136[7:0]) +
	( 7'sd 42) * $signed(input_fmap_137[7:0]) +
	( 14'sd 7738) * $signed(input_fmap_138[7:0]) +
	( 15'sd 15221) * $signed(input_fmap_139[7:0]) +
	( 16'sd 17394) * $signed(input_fmap_140[7:0]) +
	( 16'sd 26554) * $signed(input_fmap_141[7:0]) +
	( 16'sd 23308) * $signed(input_fmap_142[7:0]) +
	( 15'sd 12458) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5679) * $signed(input_fmap_144[7:0]) +
	( 15'sd 10188) * $signed(input_fmap_145[7:0]) +
	( 16'sd 32230) * $signed(input_fmap_146[7:0]) +
	( 16'sd 26498) * $signed(input_fmap_147[7:0]) +
	( 14'sd 7173) * $signed(input_fmap_148[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_149[7:0]) +
	( 13'sd 2851) * $signed(input_fmap_150[7:0]) +
	( 16'sd 22395) * $signed(input_fmap_151[7:0]) +
	( 15'sd 9499) * $signed(input_fmap_152[7:0]) +
	( 15'sd 14519) * $signed(input_fmap_153[7:0]) +
	( 16'sd 30608) * $signed(input_fmap_154[7:0]) +
	( 16'sd 25437) * $signed(input_fmap_155[7:0]) +
	( 10'sd 461) * $signed(input_fmap_156[7:0]) +
	( 16'sd 21268) * $signed(input_fmap_157[7:0]) +
	( 15'sd 13708) * $signed(input_fmap_158[7:0]) +
	( 13'sd 3793) * $signed(input_fmap_159[7:0]) +
	( 15'sd 13300) * $signed(input_fmap_160[7:0]) +
	( 14'sd 5438) * $signed(input_fmap_161[7:0]) +
	( 16'sd 18236) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27871) * $signed(input_fmap_163[7:0]) +
	( 14'sd 4409) * $signed(input_fmap_164[7:0]) +
	( 16'sd 20249) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30774) * $signed(input_fmap_166[7:0]) +
	( 14'sd 8077) * $signed(input_fmap_167[7:0]) +
	( 16'sd 28211) * $signed(input_fmap_168[7:0]) +
	( 15'sd 14428) * $signed(input_fmap_169[7:0]) +
	( 16'sd 31672) * $signed(input_fmap_170[7:0]) +
	( 14'sd 7520) * $signed(input_fmap_171[7:0]) +
	( 16'sd 23498) * $signed(input_fmap_172[7:0]) +
	( 16'sd 19166) * $signed(input_fmap_173[7:0]) +
	( 14'sd 7980) * $signed(input_fmap_174[7:0]) +
	( 15'sd 9439) * $signed(input_fmap_175[7:0]) +
	( 16'sd 18528) * $signed(input_fmap_176[7:0]) +
	( 15'sd 11359) * $signed(input_fmap_177[7:0]) +
	( 14'sd 6401) * $signed(input_fmap_178[7:0]) +
	( 16'sd 21697) * $signed(input_fmap_179[7:0]) +
	( 16'sd 19726) * $signed(input_fmap_180[7:0]) +
	( 16'sd 25353) * $signed(input_fmap_181[7:0]) +
	( 16'sd 32149) * $signed(input_fmap_182[7:0]) +
	( 16'sd 26624) * $signed(input_fmap_183[7:0]) +
	( 12'sd 1779) * $signed(input_fmap_184[7:0]) +
	( 16'sd 32581) * $signed(input_fmap_185[7:0]) +
	( 16'sd 32180) * $signed(input_fmap_186[7:0]) +
	( 16'sd 26968) * $signed(input_fmap_187[7:0]) +
	( 16'sd 23256) * $signed(input_fmap_188[7:0]) +
	( 15'sd 14566) * $signed(input_fmap_189[7:0]) +
	( 16'sd 22849) * $signed(input_fmap_190[7:0]) +
	( 15'sd 12886) * $signed(input_fmap_191[7:0]) +
	( 15'sd 15252) * $signed(input_fmap_192[7:0]) +
	( 16'sd 30716) * $signed(input_fmap_193[7:0]) +
	( 16'sd 31557) * $signed(input_fmap_194[7:0]) +
	( 14'sd 7466) * $signed(input_fmap_195[7:0]) +
	( 14'sd 7531) * $signed(input_fmap_196[7:0]) +
	( 16'sd 26077) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5923) * $signed(input_fmap_198[7:0]) +
	( 16'sd 31364) * $signed(input_fmap_199[7:0]) +
	( 15'sd 12461) * $signed(input_fmap_200[7:0]) +
	( 16'sd 31525) * $signed(input_fmap_201[7:0]) +
	( 16'sd 19613) * $signed(input_fmap_202[7:0]) +
	( 16'sd 26501) * $signed(input_fmap_203[7:0]) +
	( 11'sd 651) * $signed(input_fmap_204[7:0]) +
	( 16'sd 24471) * $signed(input_fmap_205[7:0]) +
	( 16'sd 25817) * $signed(input_fmap_206[7:0]) +
	( 16'sd 28670) * $signed(input_fmap_207[7:0]) +
	( 16'sd 25210) * $signed(input_fmap_208[7:0]) +
	( 16'sd 20803) * $signed(input_fmap_209[7:0]) +
	( 14'sd 5685) * $signed(input_fmap_210[7:0]) +
	( 15'sd 15051) * $signed(input_fmap_211[7:0]) +
	( 16'sd 16483) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3403) * $signed(input_fmap_213[7:0]) +
	( 16'sd 30209) * $signed(input_fmap_214[7:0]) +
	( 16'sd 22773) * $signed(input_fmap_215[7:0]) +
	( 14'sd 4895) * $signed(input_fmap_216[7:0]) +
	( 13'sd 3304) * $signed(input_fmap_217[7:0]) +
	( 16'sd 22220) * $signed(input_fmap_218[7:0]) +
	( 16'sd 29962) * $signed(input_fmap_219[7:0]) +
	( 16'sd 29648) * $signed(input_fmap_220[7:0]) +
	( 16'sd 27500) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5198) * $signed(input_fmap_222[7:0]) +
	( 16'sd 22176) * $signed(input_fmap_223[7:0]) +
	( 15'sd 8352) * $signed(input_fmap_224[7:0]) +
	( 15'sd 9499) * $signed(input_fmap_225[7:0]) +
	( 13'sd 3472) * $signed(input_fmap_226[7:0]) +
	( 16'sd 20488) * $signed(input_fmap_227[7:0]) +
	( 12'sd 1646) * $signed(input_fmap_228[7:0]) +
	( 16'sd 25231) * $signed(input_fmap_229[7:0]) +
	( 16'sd 25209) * $signed(input_fmap_230[7:0]) +
	( 16'sd 24887) * $signed(input_fmap_231[7:0]) +
	( 16'sd 28730) * $signed(input_fmap_232[7:0]) +
	( 16'sd 18462) * $signed(input_fmap_233[7:0]) +
	( 14'sd 4784) * $signed(input_fmap_234[7:0]) +
	( 13'sd 3228) * $signed(input_fmap_235[7:0]) +
	( 16'sd 25338) * $signed(input_fmap_236[7:0]) +
	( 13'sd 4053) * $signed(input_fmap_237[7:0]) +
	( 16'sd 31867) * $signed(input_fmap_238[7:0]) +
	( 15'sd 14149) * $signed(input_fmap_239[7:0]) +
	( 15'sd 9969) * $signed(input_fmap_240[7:0]) +
	( 15'sd 9627) * $signed(input_fmap_241[7:0]) +
	( 13'sd 4091) * $signed(input_fmap_242[7:0]) +
	( 14'sd 6289) * $signed(input_fmap_243[7:0]) +
	( 14'sd 5161) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24410) * $signed(input_fmap_245[7:0]) +
	( 15'sd 11780) * $signed(input_fmap_246[7:0]) +
	( 14'sd 6373) * $signed(input_fmap_247[7:0]) +
	( 15'sd 14306) * $signed(input_fmap_248[7:0]) +
	( 14'sd 6817) * $signed(input_fmap_249[7:0]) +
	( 16'sd 29242) * $signed(input_fmap_250[7:0]) +
	( 15'sd 16255) * $signed(input_fmap_251[7:0]) +
	( 16'sd 27516) * $signed(input_fmap_252[7:0]) +
	( 16'sd 21781) * $signed(input_fmap_253[7:0]) +
	( 13'sd 2351) * $signed(input_fmap_254[7:0]) +
	( 16'sd 20102) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_251;
assign conv_mac_251 = 
	( 16'sd 27756) * $signed(input_fmap_0[7:0]) +
	( 13'sd 3955) * $signed(input_fmap_1[7:0]) +
	( 16'sd 31383) * $signed(input_fmap_2[7:0]) +
	( 16'sd 27736) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32150) * $signed(input_fmap_4[7:0]) +
	( 15'sd 15207) * $signed(input_fmap_5[7:0]) +
	( 11'sd 876) * $signed(input_fmap_6[7:0]) +
	( 16'sd 19087) * $signed(input_fmap_7[7:0]) +
	( 16'sd 18485) * $signed(input_fmap_8[7:0]) +
	( 16'sd 27461) * $signed(input_fmap_9[7:0]) +
	( 16'sd 17339) * $signed(input_fmap_10[7:0]) +
	( 16'sd 19412) * $signed(input_fmap_11[7:0]) +
	( 16'sd 23228) * $signed(input_fmap_12[7:0]) +
	( 16'sd 28564) * $signed(input_fmap_13[7:0]) +
	( 14'sd 4574) * $signed(input_fmap_14[7:0]) +
	( 16'sd 29537) * $signed(input_fmap_15[7:0]) +
	( 13'sd 4010) * $signed(input_fmap_16[7:0]) +
	( 15'sd 11655) * $signed(input_fmap_17[7:0]) +
	( 16'sd 17280) * $signed(input_fmap_18[7:0]) +
	( 14'sd 6305) * $signed(input_fmap_19[7:0]) +
	( 16'sd 20288) * $signed(input_fmap_20[7:0]) +
	( 12'sd 1258) * $signed(input_fmap_21[7:0]) +
	( 15'sd 11252) * $signed(input_fmap_22[7:0]) +
	( 16'sd 23646) * $signed(input_fmap_23[7:0]) +
	( 16'sd 20350) * $signed(input_fmap_24[7:0]) +
	( 16'sd 32277) * $signed(input_fmap_25[7:0]) +
	( 16'sd 28026) * $signed(input_fmap_26[7:0]) +
	( 16'sd 21976) * $signed(input_fmap_27[7:0]) +
	( 16'sd 30720) * $signed(input_fmap_28[7:0]) +
	( 16'sd 21594) * $signed(input_fmap_29[7:0]) +
	( 16'sd 19088) * $signed(input_fmap_30[7:0]) +
	( 15'sd 12362) * $signed(input_fmap_31[7:0]) +
	( 15'sd 15822) * $signed(input_fmap_32[7:0]) +
	( 8'sd 78) * $signed(input_fmap_33[7:0]) +
	( 16'sd 31124) * $signed(input_fmap_34[7:0]) +
	( 16'sd 21180) * $signed(input_fmap_35[7:0]) +
	( 14'sd 7945) * $signed(input_fmap_36[7:0]) +
	( 15'sd 9283) * $signed(input_fmap_37[7:0]) +
	( 15'sd 8246) * $signed(input_fmap_38[7:0]) +
	( 16'sd 24332) * $signed(input_fmap_39[7:0]) +
	( 15'sd 11720) * $signed(input_fmap_40[7:0]) +
	( 16'sd 30649) * $signed(input_fmap_41[7:0]) +
	( 15'sd 14005) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26552) * $signed(input_fmap_43[7:0]) +
	( 13'sd 4089) * $signed(input_fmap_44[7:0]) +
	( 16'sd 21726) * $signed(input_fmap_45[7:0]) +
	( 15'sd 16285) * $signed(input_fmap_46[7:0]) +
	( 13'sd 3769) * $signed(input_fmap_47[7:0]) +
	( 16'sd 19708) * $signed(input_fmap_48[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_49[7:0]) +
	( 15'sd 10197) * $signed(input_fmap_50[7:0]) +
	( 15'sd 14290) * $signed(input_fmap_51[7:0]) +
	( 16'sd 32618) * $signed(input_fmap_52[7:0]) +
	( 16'sd 24162) * $signed(input_fmap_53[7:0]) +
	( 15'sd 11786) * $signed(input_fmap_54[7:0]) +
	( 11'sd 620) * $signed(input_fmap_55[7:0]) +
	( 16'sd 17177) * $signed(input_fmap_56[7:0]) +
	( 11'sd 832) * $signed(input_fmap_57[7:0]) +
	( 15'sd 10047) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21600) * $signed(input_fmap_59[7:0]) +
	( 14'sd 6804) * $signed(input_fmap_60[7:0]) +
	( 15'sd 12656) * $signed(input_fmap_61[7:0]) +
	( 15'sd 8941) * $signed(input_fmap_62[7:0]) +
	( 16'sd 25181) * $signed(input_fmap_63[7:0]) +
	( 15'sd 11145) * $signed(input_fmap_64[7:0]) +
	( 13'sd 4068) * $signed(input_fmap_65[7:0]) +
	( 15'sd 14356) * $signed(input_fmap_66[7:0]) +
	( 16'sd 22446) * $signed(input_fmap_67[7:0]) +
	( 16'sd 25039) * $signed(input_fmap_68[7:0]) +
	( 16'sd 31564) * $signed(input_fmap_69[7:0]) +
	( 14'sd 7011) * $signed(input_fmap_70[7:0]) +
	( 16'sd 17526) * $signed(input_fmap_71[7:0]) +
	( 15'sd 13843) * $signed(input_fmap_72[7:0]) +
	( 16'sd 21226) * $signed(input_fmap_73[7:0]) +
	( 16'sd 20133) * $signed(input_fmap_74[7:0]) +
	( 16'sd 24567) * $signed(input_fmap_75[7:0]) +
	( 15'sd 8257) * $signed(input_fmap_76[7:0]) +
	( 16'sd 22522) * $signed(input_fmap_77[7:0]) +
	( 16'sd 21547) * $signed(input_fmap_78[7:0]) +
	( 16'sd 17081) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19042) * $signed(input_fmap_80[7:0]) +
	( 15'sd 12550) * $signed(input_fmap_81[7:0]) +
	( 16'sd 26771) * $signed(input_fmap_82[7:0]) +
	( 16'sd 28690) * $signed(input_fmap_83[7:0]) +
	( 14'sd 8062) * $signed(input_fmap_84[7:0]) +
	( 15'sd 12059) * $signed(input_fmap_85[7:0]) +
	( 16'sd 32047) * $signed(input_fmap_86[7:0]) +
	( 15'sd 15998) * $signed(input_fmap_87[7:0]) +
	( 15'sd 10386) * $signed(input_fmap_88[7:0]) +
	( 16'sd 19614) * $signed(input_fmap_89[7:0]) +
	( 16'sd 29950) * $signed(input_fmap_90[7:0]) +
	( 16'sd 16751) * $signed(input_fmap_91[7:0]) +
	( 16'sd 31613) * $signed(input_fmap_92[7:0]) +
	( 16'sd 20041) * $signed(input_fmap_93[7:0]) +
	( 15'sd 13228) * $signed(input_fmap_94[7:0]) +
	( 16'sd 20694) * $signed(input_fmap_95[7:0]) +
	( 14'sd 6984) * $signed(input_fmap_96[7:0]) +
	( 16'sd 19692) * $signed(input_fmap_97[7:0]) +
	( 16'sd 23415) * $signed(input_fmap_98[7:0]) +
	( 16'sd 21545) * $signed(input_fmap_99[7:0]) +
	( 15'sd 15423) * $signed(input_fmap_100[7:0]) +
	( 16'sd 31356) * $signed(input_fmap_101[7:0]) +
	( 16'sd 27717) * $signed(input_fmap_102[7:0]) +
	( 16'sd 18505) * $signed(input_fmap_103[7:0]) +
	( 16'sd 16453) * $signed(input_fmap_104[7:0]) +
	( 16'sd 28741) * $signed(input_fmap_105[7:0]) +
	( 14'sd 6127) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7687) * $signed(input_fmap_107[7:0]) +
	( 15'sd 9346) * $signed(input_fmap_108[7:0]) +
	( 16'sd 23841) * $signed(input_fmap_109[7:0]) +
	( 16'sd 27081) * $signed(input_fmap_110[7:0]) +
	( 16'sd 22519) * $signed(input_fmap_111[7:0]) +
	( 16'sd 27108) * $signed(input_fmap_112[7:0]) +
	( 14'sd 5488) * $signed(input_fmap_113[7:0]) +
	( 16'sd 16496) * $signed(input_fmap_114[7:0]) +
	( 16'sd 23019) * $signed(input_fmap_115[7:0]) +
	( 16'sd 21095) * $signed(input_fmap_116[7:0]) +
	( 11'sd 721) * $signed(input_fmap_117[7:0]) +
	( 16'sd 32518) * $signed(input_fmap_118[7:0]) +
	( 14'sd 5314) * $signed(input_fmap_119[7:0]) +
	( 15'sd 8991) * $signed(input_fmap_120[7:0]) +
	( 15'sd 15404) * $signed(input_fmap_121[7:0]) +
	( 12'sd 1921) * $signed(input_fmap_122[7:0]) +
	( 16'sd 28181) * $signed(input_fmap_123[7:0]) +
	( 16'sd 23296) * $signed(input_fmap_124[7:0]) +
	( 16'sd 20407) * $signed(input_fmap_125[7:0]) +
	( 14'sd 4294) * $signed(input_fmap_126[7:0]) +
	( 16'sd 21566) * $signed(input_fmap_127[7:0]) +
	( 13'sd 3015) * $signed(input_fmap_128[7:0]) +
	( 15'sd 9940) * $signed(input_fmap_129[7:0]) +
	( 15'sd 15488) * $signed(input_fmap_130[7:0]) +
	( 16'sd 21074) * $signed(input_fmap_131[7:0]) +
	( 13'sd 3209) * $signed(input_fmap_132[7:0]) +
	( 16'sd 29926) * $signed(input_fmap_133[7:0]) +
	( 16'sd 27870) * $signed(input_fmap_134[7:0]) +
	( 16'sd 23700) * $signed(input_fmap_135[7:0]) +
	( 15'sd 9931) * $signed(input_fmap_136[7:0]) +
	( 16'sd 24637) * $signed(input_fmap_137[7:0]) +
	( 15'sd 11009) * $signed(input_fmap_138[7:0]) +
	( 16'sd 17582) * $signed(input_fmap_139[7:0]) +
	( 14'sd 5872) * $signed(input_fmap_140[7:0]) +
	( 14'sd 7070) * $signed(input_fmap_141[7:0]) +
	( 15'sd 8357) * $signed(input_fmap_142[7:0]) +
	( 16'sd 18742) * $signed(input_fmap_143[7:0]) +
	( 15'sd 12286) * $signed(input_fmap_144[7:0]) +
	( 16'sd 20191) * $signed(input_fmap_145[7:0]) +
	( 12'sd 1919) * $signed(input_fmap_146[7:0]) +
	( 16'sd 21085) * $signed(input_fmap_147[7:0]) +
	( 14'sd 5463) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25310) * $signed(input_fmap_149[7:0]) +
	( 16'sd 23086) * $signed(input_fmap_150[7:0]) +
	( 16'sd 19712) * $signed(input_fmap_151[7:0]) +
	( 16'sd 23276) * $signed(input_fmap_152[7:0]) +
	( 15'sd 12731) * $signed(input_fmap_153[7:0]) +
	( 14'sd 7848) * $signed(input_fmap_154[7:0]) +
	( 15'sd 10304) * $signed(input_fmap_155[7:0]) +
	( 16'sd 27148) * $signed(input_fmap_156[7:0]) +
	( 14'sd 7429) * $signed(input_fmap_157[7:0]) +
	( 15'sd 8855) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6735) * $signed(input_fmap_159[7:0]) +
	( 16'sd 26487) * $signed(input_fmap_160[7:0]) +
	( 15'sd 9009) * $signed(input_fmap_161[7:0]) +
	( 14'sd 7408) * $signed(input_fmap_162[7:0]) +
	( 8'sd 86) * $signed(input_fmap_163[7:0]) +
	( 15'sd 10007) * $signed(input_fmap_164[7:0]) +
	( 15'sd 10143) * $signed(input_fmap_165[7:0]) +
	( 16'sd 30394) * $signed(input_fmap_166[7:0]) +
	( 16'sd 28169) * $signed(input_fmap_167[7:0]) +
	( 16'sd 26028) * $signed(input_fmap_168[7:0]) +
	( 16'sd 21578) * $signed(input_fmap_169[7:0]) +
	( 15'sd 9143) * $signed(input_fmap_170[7:0]) +
	( 12'sd 1874) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1487) * $signed(input_fmap_172[7:0]) +
	( 14'sd 6939) * $signed(input_fmap_173[7:0]) +
	( 15'sd 12907) * $signed(input_fmap_174[7:0]) +
	( 14'sd 6002) * $signed(input_fmap_175[7:0]) +
	( 7'sd 45) * $signed(input_fmap_176[7:0]) +
	( 16'sd 17407) * $signed(input_fmap_177[7:0]) +
	( 16'sd 27012) * $signed(input_fmap_178[7:0]) +
	( 16'sd 22511) * $signed(input_fmap_179[7:0]) +
	( 15'sd 15909) * $signed(input_fmap_180[7:0]) +
	( 12'sd 2037) * $signed(input_fmap_181[7:0]) +
	( 11'sd 630) * $signed(input_fmap_182[7:0]) +
	( 16'sd 21887) * $signed(input_fmap_183[7:0]) +
	( 15'sd 14007) * $signed(input_fmap_184[7:0]) +
	( 15'sd 14429) * $signed(input_fmap_185[7:0]) +
	( 15'sd 8510) * $signed(input_fmap_186[7:0]) +
	( 16'sd 21651) * $signed(input_fmap_187[7:0]) +
	( 15'sd 11679) * $signed(input_fmap_188[7:0]) +
	( 16'sd 19527) * $signed(input_fmap_189[7:0]) +
	( 14'sd 7978) * $signed(input_fmap_190[7:0]) +
	( 13'sd 3598) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19665) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22250) * $signed(input_fmap_193[7:0]) +
	( 16'sd 30281) * $signed(input_fmap_194[7:0]) +
	( 11'sd 594) * $signed(input_fmap_195[7:0]) +
	( 12'sd 1969) * $signed(input_fmap_196[7:0]) +
	( 16'sd 29074) * $signed(input_fmap_197[7:0]) +
	( 16'sd 30094) * $signed(input_fmap_198[7:0]) +
	( 15'sd 14394) * $signed(input_fmap_199[7:0]) +
	( 16'sd 25363) * $signed(input_fmap_200[7:0]) +
	( 12'sd 1222) * $signed(input_fmap_201[7:0]) +
	( 16'sd 23054) * $signed(input_fmap_202[7:0]) +
	( 16'sd 23905) * $signed(input_fmap_203[7:0]) +
	( 14'sd 4394) * $signed(input_fmap_204[7:0]) +
	( 16'sd 31981) * $signed(input_fmap_205[7:0]) +
	( 16'sd 24674) * $signed(input_fmap_206[7:0]) +
	( 16'sd 22251) * $signed(input_fmap_207[7:0]) +
	( 14'sd 8104) * $signed(input_fmap_208[7:0]) +
	( 16'sd 24466) * $signed(input_fmap_209[7:0]) +
	( 11'sd 687) * $signed(input_fmap_210[7:0]) +
	( 16'sd 16757) * $signed(input_fmap_211[7:0]) +
	( 16'sd 21007) * $signed(input_fmap_212[7:0]) +
	( 13'sd 3443) * $signed(input_fmap_213[7:0]) +
	( 12'sd 1719) * $signed(input_fmap_214[7:0]) +
	( 15'sd 11793) * $signed(input_fmap_215[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_216[7:0]) +
	( 13'sd 2983) * $signed(input_fmap_217[7:0]) +
	( 16'sd 31872) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15058) * $signed(input_fmap_219[7:0]) +
	( 16'sd 27208) * $signed(input_fmap_220[7:0]) +
	( 15'sd 10873) * $signed(input_fmap_221[7:0]) +
	( 14'sd 5550) * $signed(input_fmap_222[7:0]) +
	( 16'sd 18839) * $signed(input_fmap_223[7:0]) +
	( 16'sd 16456) * $signed(input_fmap_224[7:0]) +
	( 16'sd 20049) * $signed(input_fmap_225[7:0]) +
	( 15'sd 11715) * $signed(input_fmap_226[7:0]) +
	( 16'sd 27561) * $signed(input_fmap_227[7:0]) +
	( 16'sd 26765) * $signed(input_fmap_228[7:0]) +
	( 16'sd 28449) * $signed(input_fmap_229[7:0]) +
	( 16'sd 29970) * $signed(input_fmap_230[7:0]) +
	( 15'sd 13974) * $signed(input_fmap_231[7:0]) +
	( 15'sd 16202) * $signed(input_fmap_232[7:0]) +
	( 16'sd 32568) * $signed(input_fmap_233[7:0]) +
	( 13'sd 2402) * $signed(input_fmap_234[7:0]) +
	( 14'sd 4279) * $signed(input_fmap_235[7:0]) +
	( 16'sd 28129) * $signed(input_fmap_236[7:0]) +
	( 16'sd 26878) * $signed(input_fmap_237[7:0]) +
	( 15'sd 13390) * $signed(input_fmap_238[7:0]) +
	( 16'sd 19346) * $signed(input_fmap_239[7:0]) +
	( 16'sd 20521) * $signed(input_fmap_240[7:0]) +
	( 16'sd 16517) * $signed(input_fmap_241[7:0]) +
	( 15'sd 11910) * $signed(input_fmap_242[7:0]) +
	( 14'sd 5676) * $signed(input_fmap_243[7:0]) +
	( 11'sd 645) * $signed(input_fmap_244[7:0]) +
	( 16'sd 16546) * $signed(input_fmap_245[7:0]) +
	( 15'sd 13679) * $signed(input_fmap_246[7:0]) +
	( 13'sd 3460) * $signed(input_fmap_247[7:0]) +
	( 16'sd 27242) * $signed(input_fmap_248[7:0]) +
	( 14'sd 4658) * $signed(input_fmap_249[7:0]) +
	( 16'sd 22893) * $signed(input_fmap_250[7:0]) +
	( 15'sd 11050) * $signed(input_fmap_251[7:0]) +
	( 15'sd 8769) * $signed(input_fmap_252[7:0]) +
	( 15'sd 9371) * $signed(input_fmap_253[7:0]) +
	( 15'sd 12528) * $signed(input_fmap_254[7:0]) +
	( 16'sd 26642) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_252;
assign conv_mac_252 = 
	( 16'sd 20072) * $signed(input_fmap_0[7:0]) +
	( 16'sd 23448) * $signed(input_fmap_1[7:0]) +
	( 14'sd 4781) * $signed(input_fmap_2[7:0]) +
	( 14'sd 6903) * $signed(input_fmap_3[7:0]) +
	( 14'sd 5946) * $signed(input_fmap_4[7:0]) +
	( 16'sd 17193) * $signed(input_fmap_5[7:0]) +
	( 14'sd 4173) * $signed(input_fmap_6[7:0]) +
	( 15'sd 8691) * $signed(input_fmap_7[7:0]) +
	( 15'sd 11383) * $signed(input_fmap_8[7:0]) +
	( 14'sd 4502) * $signed(input_fmap_9[7:0]) +
	( 15'sd 10020) * $signed(input_fmap_10[7:0]) +
	( 16'sd 25748) * $signed(input_fmap_11[7:0]) +
	( 14'sd 5252) * $signed(input_fmap_12[7:0]) +
	( 15'sd 15891) * $signed(input_fmap_13[7:0]) +
	( 15'sd 15191) * $signed(input_fmap_14[7:0]) +
	( 16'sd 24329) * $signed(input_fmap_15[7:0]) +
	( 15'sd 12989) * $signed(input_fmap_16[7:0]) +
	( 13'sd 2888) * $signed(input_fmap_17[7:0]) +
	( 14'sd 7797) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13492) * $signed(input_fmap_19[7:0]) +
	( 15'sd 11983) * $signed(input_fmap_20[7:0]) +
	( 13'sd 3009) * $signed(input_fmap_21[7:0]) +
	( 15'sd 14896) * $signed(input_fmap_22[7:0]) +
	( 13'sd 2983) * $signed(input_fmap_23[7:0]) +
	( 16'sd 26937) * $signed(input_fmap_24[7:0]) +
	( 16'sd 19607) * $signed(input_fmap_25[7:0]) +
	( 15'sd 15813) * $signed(input_fmap_26[7:0]) +
	( 16'sd 17179) * $signed(input_fmap_27[7:0]) +
	( 16'sd 18470) * $signed(input_fmap_28[7:0]) +
	( 15'sd 15240) * $signed(input_fmap_29[7:0]) +
	( 16'sd 26777) * $signed(input_fmap_30[7:0]) +
	( 14'sd 5002) * $signed(input_fmap_31[7:0]) +
	( 5'sd 13) * $signed(input_fmap_32[7:0]) +
	( 16'sd 26457) * $signed(input_fmap_33[7:0]) +
	( 13'sd 3010) * $signed(input_fmap_34[7:0]) +
	( 15'sd 11541) * $signed(input_fmap_35[7:0]) +
	( 16'sd 20027) * $signed(input_fmap_36[7:0]) +
	( 16'sd 29629) * $signed(input_fmap_37[7:0]) +
	( 16'sd 22745) * $signed(input_fmap_38[7:0]) +
	( 15'sd 13405) * $signed(input_fmap_39[7:0]) +
	( 14'sd 4881) * $signed(input_fmap_40[7:0]) +
	( 15'sd 11680) * $signed(input_fmap_41[7:0]) +
	( 15'sd 15416) * $signed(input_fmap_42[7:0]) +
	( 16'sd 24025) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17707) * $signed(input_fmap_44[7:0]) +
	( 16'sd 23826) * $signed(input_fmap_45[7:0]) +
	( 16'sd 23010) * $signed(input_fmap_46[7:0]) +
	( 15'sd 12865) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14062) * $signed(input_fmap_48[7:0]) +
	( 16'sd 23547) * $signed(input_fmap_49[7:0]) +
	( 16'sd 26401) * $signed(input_fmap_50[7:0]) +
	( 14'sd 7664) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20965) * $signed(input_fmap_52[7:0]) +
	( 15'sd 15661) * $signed(input_fmap_53[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_54[7:0]) +
	( 16'sd 30258) * $signed(input_fmap_55[7:0]) +
	( 16'sd 19300) * $signed(input_fmap_56[7:0]) +
	( 16'sd 18130) * $signed(input_fmap_57[7:0]) +
	( 16'sd 28151) * $signed(input_fmap_58[7:0]) +
	( 16'sd 22817) * $signed(input_fmap_59[7:0]) +
	( 16'sd 28810) * $signed(input_fmap_60[7:0]) +
	( 15'sd 13600) * $signed(input_fmap_61[7:0]) +
	( 15'sd 11055) * $signed(input_fmap_62[7:0]) +
	( 14'sd 6865) * $signed(input_fmap_63[7:0]) +
	( 16'sd 28563) * $signed(input_fmap_64[7:0]) +
	( 15'sd 10835) * $signed(input_fmap_65[7:0]) +
	( 16'sd 32314) * $signed(input_fmap_66[7:0]) +
	( 14'sd 7063) * $signed(input_fmap_67[7:0]) +
	( 16'sd 18117) * $signed(input_fmap_68[7:0]) +
	( 16'sd 19901) * $signed(input_fmap_69[7:0]) +
	( 11'sd 883) * $signed(input_fmap_70[7:0]) +
	( 16'sd 24896) * $signed(input_fmap_71[7:0]) +
	( 16'sd 23058) * $signed(input_fmap_72[7:0]) +
	( 14'sd 7411) * $signed(input_fmap_73[7:0]) +
	( 14'sd 5130) * $signed(input_fmap_74[7:0]) +
	( 14'sd 5886) * $signed(input_fmap_75[7:0]) +
	( 16'sd 31911) * $signed(input_fmap_76[7:0]) +
	( 12'sd 1094) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9202) * $signed(input_fmap_78[7:0]) +
	( 16'sd 16529) * $signed(input_fmap_79[7:0]) +
	( 14'sd 4279) * $signed(input_fmap_80[7:0]) +
	( 16'sd 28330) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22573) * $signed(input_fmap_82[7:0]) +
	( 16'sd 18322) * $signed(input_fmap_83[7:0]) +
	( 16'sd 23220) * $signed(input_fmap_84[7:0]) +
	( 16'sd 22939) * $signed(input_fmap_85[7:0]) +
	( 15'sd 13125) * $signed(input_fmap_86[7:0]) +
	( 15'sd 14861) * $signed(input_fmap_87[7:0]) +
	( 16'sd 22422) * $signed(input_fmap_88[7:0]) +
	( 15'sd 9366) * $signed(input_fmap_89[7:0]) +
	( 15'sd 10172) * $signed(input_fmap_90[7:0]) +
	( 16'sd 26496) * $signed(input_fmap_91[7:0]) +
	( 16'sd 28045) * $signed(input_fmap_92[7:0]) +
	( 16'sd 24421) * $signed(input_fmap_93[7:0]) +
	( 15'sd 12985) * $signed(input_fmap_94[7:0]) +
	( 16'sd 30903) * $signed(input_fmap_95[7:0]) +
	( 16'sd 19848) * $signed(input_fmap_96[7:0]) +
	( 15'sd 12374) * $signed(input_fmap_97[7:0]) +
	( 14'sd 7908) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29991) * $signed(input_fmap_99[7:0]) +
	( 16'sd 30227) * $signed(input_fmap_100[7:0]) +
	( 16'sd 17816) * $signed(input_fmap_101[7:0]) +
	( 16'sd 18016) * $signed(input_fmap_102[7:0]) +
	( 15'sd 10645) * $signed(input_fmap_103[7:0]) +
	( 16'sd 22405) * $signed(input_fmap_104[7:0]) +
	( 16'sd 27399) * $signed(input_fmap_105[7:0]) +
	( 16'sd 17911) * $signed(input_fmap_106[7:0]) +
	( 14'sd 7351) * $signed(input_fmap_107[7:0]) +
	( 16'sd 19386) * $signed(input_fmap_108[7:0]) +
	( 16'sd 21558) * $signed(input_fmap_109[7:0]) +
	( 16'sd 20461) * $signed(input_fmap_110[7:0]) +
	( 16'sd 26869) * $signed(input_fmap_111[7:0]) +
	( 16'sd 29359) * $signed(input_fmap_112[7:0]) +
	( 16'sd 18193) * $signed(input_fmap_113[7:0]) +
	( 15'sd 9007) * $signed(input_fmap_114[7:0]) +
	( 16'sd 27136) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29588) * $signed(input_fmap_116[7:0]) +
	( 16'sd 23508) * $signed(input_fmap_117[7:0]) +
	( 16'sd 17983) * $signed(input_fmap_118[7:0]) +
	( 16'sd 32203) * $signed(input_fmap_119[7:0]) +
	( 15'sd 12128) * $signed(input_fmap_120[7:0]) +
	( 14'sd 7634) * $signed(input_fmap_121[7:0]) +
	( 16'sd 22782) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27256) * $signed(input_fmap_123[7:0]) +
	( 16'sd 18654) * $signed(input_fmap_124[7:0]) +
	( 16'sd 25067) * $signed(input_fmap_125[7:0]) +
	( 15'sd 15758) * $signed(input_fmap_126[7:0]) +
	( 16'sd 26533) * $signed(input_fmap_127[7:0]) +
	( 16'sd 26582) * $signed(input_fmap_128[7:0]) +
	( 16'sd 23917) * $signed(input_fmap_129[7:0]) +
	( 9'sd 167) * $signed(input_fmap_130[7:0]) +
	( 14'sd 7382) * $signed(input_fmap_131[7:0]) +
	( 12'sd 1800) * $signed(input_fmap_132[7:0]) +
	( 15'sd 12683) * $signed(input_fmap_133[7:0]) +
	( 16'sd 18544) * $signed(input_fmap_134[7:0]) +
	( 16'sd 18739) * $signed(input_fmap_135[7:0]) +
	( 16'sd 32406) * $signed(input_fmap_136[7:0]) +
	( 14'sd 7069) * $signed(input_fmap_137[7:0]) +
	( 16'sd 20104) * $signed(input_fmap_138[7:0]) +
	( 15'sd 10481) * $signed(input_fmap_139[7:0]) +
	( 13'sd 4045) * $signed(input_fmap_140[7:0]) +
	( 16'sd 31323) * $signed(input_fmap_141[7:0]) +
	( 14'sd 5228) * $signed(input_fmap_142[7:0]) +
	( 16'sd 29501) * $signed(input_fmap_143[7:0]) +
	( 15'sd 14749) * $signed(input_fmap_144[7:0]) +
	( 16'sd 17251) * $signed(input_fmap_145[7:0]) +
	( 16'sd 31314) * $signed(input_fmap_146[7:0]) +
	( 12'sd 1799) * $signed(input_fmap_147[7:0]) +
	( 15'sd 15614) * $signed(input_fmap_148[7:0]) +
	( 16'sd 24182) * $signed(input_fmap_149[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_150[7:0]) +
	( 16'sd 21447) * $signed(input_fmap_151[7:0]) +
	( 16'sd 25280) * $signed(input_fmap_152[7:0]) +
	( 16'sd 31130) * $signed(input_fmap_153[7:0]) +
	( 15'sd 10731) * $signed(input_fmap_154[7:0]) +
	( 16'sd 21493) * $signed(input_fmap_155[7:0]) +
	( 14'sd 5648) * $signed(input_fmap_156[7:0]) +
	( 13'sd 3553) * $signed(input_fmap_157[7:0]) +
	( 16'sd 20588) * $signed(input_fmap_158[7:0]) +
	( 13'sd 2805) * $signed(input_fmap_159[7:0]) +
	( 14'sd 5310) * $signed(input_fmap_160[7:0]) +
	( 16'sd 29338) * $signed(input_fmap_161[7:0]) +
	( 16'sd 24737) * $signed(input_fmap_162[7:0]) +
	( 13'sd 2725) * $signed(input_fmap_163[7:0]) +
	( 14'sd 5555) * $signed(input_fmap_164[7:0]) +
	( 16'sd 16962) * $signed(input_fmap_165[7:0]) +
	( 5'sd 8) * $signed(input_fmap_166[7:0]) +
	( 16'sd 21343) * $signed(input_fmap_167[7:0]) +
	( 15'sd 14003) * $signed(input_fmap_168[7:0]) +
	( 15'sd 11772) * $signed(input_fmap_169[7:0]) +
	( 14'sd 5497) * $signed(input_fmap_170[7:0]) +
	( 15'sd 9308) * $signed(input_fmap_171[7:0]) +
	( 12'sd 1847) * $signed(input_fmap_172[7:0]) +
	( 15'sd 8762) * $signed(input_fmap_173[7:0]) +
	( 15'sd 15201) * $signed(input_fmap_174[7:0]) +
	( 15'sd 10162) * $signed(input_fmap_175[7:0]) +
	( 13'sd 2295) * $signed(input_fmap_176[7:0]) +
	( 15'sd 9516) * $signed(input_fmap_177[7:0]) +
	( 16'sd 26908) * $signed(input_fmap_178[7:0]) +
	( 11'sd 887) * $signed(input_fmap_179[7:0]) +
	( 16'sd 22715) * $signed(input_fmap_180[7:0]) +
	( 15'sd 10833) * $signed(input_fmap_181[7:0]) +
	( 14'sd 5542) * $signed(input_fmap_182[7:0]) +
	( 16'sd 24920) * $signed(input_fmap_183[7:0]) +
	( 15'sd 11929) * $signed(input_fmap_184[7:0]) +
	( 16'sd 28528) * $signed(input_fmap_185[7:0]) +
	( 16'sd 17303) * $signed(input_fmap_186[7:0]) +
	( 16'sd 32320) * $signed(input_fmap_187[7:0]) +
	( 16'sd 30255) * $signed(input_fmap_188[7:0]) +
	( 13'sd 3769) * $signed(input_fmap_189[7:0]) +
	( 16'sd 22597) * $signed(input_fmap_190[7:0]) +
	( 15'sd 10022) * $signed(input_fmap_191[7:0]) +
	( 15'sd 12000) * $signed(input_fmap_192[7:0]) +
	( 15'sd 13254) * $signed(input_fmap_193[7:0]) +
	( 14'sd 6248) * $signed(input_fmap_194[7:0]) +
	( 15'sd 12024) * $signed(input_fmap_195[7:0]) +
	( 14'sd 6782) * $signed(input_fmap_196[7:0]) +
	( 16'sd 25069) * $signed(input_fmap_197[7:0]) +
	( 16'sd 31564) * $signed(input_fmap_198[7:0]) +
	( 11'sd 886) * $signed(input_fmap_199[7:0]) +
	( 14'sd 6999) * $signed(input_fmap_200[7:0]) +
	( 16'sd 22111) * $signed(input_fmap_201[7:0]) +
	( 16'sd 29860) * $signed(input_fmap_202[7:0]) +
	( 16'sd 19704) * $signed(input_fmap_203[7:0]) +
	( 16'sd 30390) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18979) * $signed(input_fmap_205[7:0]) +
	( 16'sd 29432) * $signed(input_fmap_206[7:0]) +
	( 13'sd 3274) * $signed(input_fmap_207[7:0]) +
	( 10'sd 453) * $signed(input_fmap_208[7:0]) +
	( 16'sd 18022) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23597) * $signed(input_fmap_210[7:0]) +
	( 16'sd 17904) * $signed(input_fmap_211[7:0]) +
	( 16'sd 20905) * $signed(input_fmap_212[7:0]) +
	( 15'sd 12353) * $signed(input_fmap_213[7:0]) +
	( 16'sd 28984) * $signed(input_fmap_214[7:0]) +
	( 15'sd 10738) * $signed(input_fmap_215[7:0]) +
	( 15'sd 14309) * $signed(input_fmap_216[7:0]) +
	( 16'sd 20942) * $signed(input_fmap_217[7:0]) +
	( 14'sd 6431) * $signed(input_fmap_218[7:0]) +
	( 14'sd 6955) * $signed(input_fmap_219[7:0]) +
	( 15'sd 14017) * $signed(input_fmap_220[7:0]) +
	( 12'sd 1428) * $signed(input_fmap_221[7:0]) +
	( 15'sd 9946) * $signed(input_fmap_222[7:0]) +
	( 16'sd 29019) * $signed(input_fmap_223[7:0]) +
	( 12'sd 1139) * $signed(input_fmap_224[7:0]) +
	( 14'sd 6850) * $signed(input_fmap_225[7:0]) +
	( 16'sd 22150) * $signed(input_fmap_226[7:0]) +
	( 15'sd 12178) * $signed(input_fmap_227[7:0]) +
	( 14'sd 6960) * $signed(input_fmap_228[7:0]) +
	( 15'sd 14228) * $signed(input_fmap_229[7:0]) +
	( 15'sd 14490) * $signed(input_fmap_230[7:0]) +
	( 15'sd 14722) * $signed(input_fmap_231[7:0]) +
	( 15'sd 14372) * $signed(input_fmap_232[7:0]) +
	( 16'sd 27100) * $signed(input_fmap_233[7:0]) +
	( 16'sd 16557) * $signed(input_fmap_234[7:0]) +
	( 16'sd 27333) * $signed(input_fmap_235[7:0]) +
	( 16'sd 18945) * $signed(input_fmap_236[7:0]) +
	( 12'sd 1318) * $signed(input_fmap_237[7:0]) +
	( 16'sd 27957) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23803) * $signed(input_fmap_239[7:0]) +
	( 16'sd 22399) * $signed(input_fmap_240[7:0]) +
	( 15'sd 13142) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27508) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25341) * $signed(input_fmap_243[7:0]) +
	( 16'sd 22560) * $signed(input_fmap_244[7:0]) +
	( 16'sd 29585) * $signed(input_fmap_245[7:0]) +
	( 15'sd 8217) * $signed(input_fmap_246[7:0]) +
	( 16'sd 24877) * $signed(input_fmap_247[7:0]) +
	( 9'sd 219) * $signed(input_fmap_248[7:0]) +
	( 15'sd 11413) * $signed(input_fmap_249[7:0]) +
	( 15'sd 8538) * $signed(input_fmap_250[7:0]) +
	( 16'sd 22307) * $signed(input_fmap_251[7:0]) +
	( 14'sd 4540) * $signed(input_fmap_252[7:0]) +
	( 16'sd 25355) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26379) * $signed(input_fmap_254[7:0]) +
	( 16'sd 22296) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_253;
assign conv_mac_253 = 
	( 16'sd 17358) * $signed(input_fmap_0[7:0]) +
	( 16'sd 30427) * $signed(input_fmap_1[7:0]) +
	( 16'sd 25581) * $signed(input_fmap_2[7:0]) +
	( 16'sd 28601) * $signed(input_fmap_3[7:0]) +
	( 14'sd 4884) * $signed(input_fmap_4[7:0]) +
	( 15'sd 11044) * $signed(input_fmap_5[7:0]) +
	( 15'sd 10013) * $signed(input_fmap_6[7:0]) +
	( 14'sd 7421) * $signed(input_fmap_7[7:0]) +
	( 14'sd 7235) * $signed(input_fmap_8[7:0]) +
	( 15'sd 10412) * $signed(input_fmap_9[7:0]) +
	( 16'sd 25664) * $signed(input_fmap_10[7:0]) +
	( 16'sd 31929) * $signed(input_fmap_11[7:0]) +
	( 15'sd 11254) * $signed(input_fmap_12[7:0]) +
	( 12'sd 2009) * $signed(input_fmap_13[7:0]) +
	( 15'sd 9354) * $signed(input_fmap_14[7:0]) +
	( 16'sd 22003) * $signed(input_fmap_15[7:0]) +
	( 15'sd 16191) * $signed(input_fmap_16[7:0]) +
	( 16'sd 23234) * $signed(input_fmap_17[7:0]) +
	( 15'sd 15278) * $signed(input_fmap_18[7:0]) +
	( 14'sd 7194) * $signed(input_fmap_19[7:0]) +
	( 15'sd 16056) * $signed(input_fmap_20[7:0]) +
	( 15'sd 13217) * $signed(input_fmap_21[7:0]) +
	( 16'sd 22839) * $signed(input_fmap_22[7:0]) +
	( 16'sd 24753) * $signed(input_fmap_23[7:0]) +
	( 14'sd 4293) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12558) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20653) * $signed(input_fmap_26[7:0]) +
	( 16'sd 16947) * $signed(input_fmap_27[7:0]) +
	( 16'sd 23658) * $signed(input_fmap_28[7:0]) +
	( 7'sd 42) * $signed(input_fmap_29[7:0]) +
	( 15'sd 9654) * $signed(input_fmap_30[7:0]) +
	( 12'sd 1854) * $signed(input_fmap_31[7:0]) +
	( 13'sd 2181) * $signed(input_fmap_32[7:0]) +
	( 14'sd 4846) * $signed(input_fmap_33[7:0]) +
	( 15'sd 11897) * $signed(input_fmap_34[7:0]) +
	( 15'sd 12154) * $signed(input_fmap_35[7:0]) +
	( 15'sd 10484) * $signed(input_fmap_36[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_37[7:0]) +
	( 16'sd 32377) * $signed(input_fmap_38[7:0]) +
	( 12'sd 1202) * $signed(input_fmap_39[7:0]) +
	( 15'sd 10599) * $signed(input_fmap_40[7:0]) +
	( 16'sd 28586) * $signed(input_fmap_41[7:0]) +
	( 15'sd 12977) * $signed(input_fmap_42[7:0]) +
	( 11'sd 576) * $signed(input_fmap_43[7:0]) +
	( 15'sd 13875) * $signed(input_fmap_44[7:0]) +
	( 15'sd 11066) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22696) * $signed(input_fmap_46[7:0]) +
	( 16'sd 17012) * $signed(input_fmap_47[7:0]) +
	( 15'sd 14978) * $signed(input_fmap_48[7:0]) +
	( 16'sd 30036) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9729) * $signed(input_fmap_50[7:0]) +
	( 16'sd 32641) * $signed(input_fmap_51[7:0]) +
	( 16'sd 24395) * $signed(input_fmap_52[7:0]) +
	( 16'sd 20755) * $signed(input_fmap_53[7:0]) +
	( 16'sd 24174) * $signed(input_fmap_54[7:0]) +
	( 16'sd 19370) * $signed(input_fmap_55[7:0]) +
	( 15'sd 13739) * $signed(input_fmap_56[7:0]) +
	( 16'sd 23151) * $signed(input_fmap_57[7:0]) +
	( 14'sd 6072) * $signed(input_fmap_58[7:0]) +
	( 16'sd 26823) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_60[7:0]) +
	( 16'sd 21289) * $signed(input_fmap_61[7:0]) +
	( 15'sd 13673) * $signed(input_fmap_62[7:0]) +
	( 15'sd 15604) * $signed(input_fmap_63[7:0]) +
	( 16'sd 21194) * $signed(input_fmap_64[7:0]) +
	( 14'sd 4994) * $signed(input_fmap_65[7:0]) +
	( 16'sd 27817) * $signed(input_fmap_66[7:0]) +
	( 16'sd 26665) * $signed(input_fmap_67[7:0]) +
	( 15'sd 9889) * $signed(input_fmap_68[7:0]) +
	( 12'sd 1902) * $signed(input_fmap_69[7:0]) +
	( 16'sd 16778) * $signed(input_fmap_70[7:0]) +
	( 12'sd 1802) * $signed(input_fmap_71[7:0]) +
	( 10'sd 399) * $signed(input_fmap_72[7:0]) +
	( 12'sd 1688) * $signed(input_fmap_73[7:0]) +
	( 13'sd 2950) * $signed(input_fmap_74[7:0]) +
	( 14'sd 7962) * $signed(input_fmap_75[7:0]) +
	( 13'sd 3796) * $signed(input_fmap_76[7:0]) +
	( 16'sd 30240) * $signed(input_fmap_77[7:0]) +
	( 16'sd 28287) * $signed(input_fmap_78[7:0]) +
	( 16'sd 29171) * $signed(input_fmap_79[7:0]) +
	( 14'sd 7526) * $signed(input_fmap_80[7:0]) +
	( 16'sd 17094) * $signed(input_fmap_81[7:0]) +
	( 16'sd 22091) * $signed(input_fmap_82[7:0]) +
	( 16'sd 21327) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5471) * $signed(input_fmap_84[7:0]) +
	( 16'sd 19597) * $signed(input_fmap_85[7:0]) +
	( 15'sd 14177) * $signed(input_fmap_86[7:0]) +
	( 16'sd 32691) * $signed(input_fmap_87[7:0]) +
	( 15'sd 9622) * $signed(input_fmap_88[7:0]) +
	( 14'sd 5957) * $signed(input_fmap_89[7:0]) +
	( 16'sd 17387) * $signed(input_fmap_90[7:0]) +
	( 15'sd 15603) * $signed(input_fmap_91[7:0]) +
	( 13'sd 3324) * $signed(input_fmap_92[7:0]) +
	( 15'sd 16052) * $signed(input_fmap_93[7:0]) +
	( 15'sd 14686) * $signed(input_fmap_94[7:0]) +
	( 16'sd 29013) * $signed(input_fmap_95[7:0]) +
	( 16'sd 28555) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11771) * $signed(input_fmap_97[7:0]) +
	( 16'sd 26371) * $signed(input_fmap_98[7:0]) +
	( 16'sd 30758) * $signed(input_fmap_99[7:0]) +
	( 16'sd 16972) * $signed(input_fmap_100[7:0]) +
	( 16'sd 25473) * $signed(input_fmap_101[7:0]) +
	( 16'sd 23443) * $signed(input_fmap_102[7:0]) +
	( 15'sd 15364) * $signed(input_fmap_103[7:0]) +
	( 16'sd 30572) * $signed(input_fmap_104[7:0]) +
	( 16'sd 24106) * $signed(input_fmap_105[7:0]) +
	( 13'sd 2611) * $signed(input_fmap_106[7:0]) +
	( 15'sd 10000) * $signed(input_fmap_107[7:0]) +
	( 16'sd 28985) * $signed(input_fmap_108[7:0]) +
	( 16'sd 24967) * $signed(input_fmap_109[7:0]) +
	( 10'sd 459) * $signed(input_fmap_110[7:0]) +
	( 16'sd 24816) * $signed(input_fmap_111[7:0]) +
	( 16'sd 23155) * $signed(input_fmap_112[7:0]) +
	( 13'sd 4011) * $signed(input_fmap_113[7:0]) +
	( 16'sd 17043) * $signed(input_fmap_114[7:0]) +
	( 13'sd 2464) * $signed(input_fmap_115[7:0]) +
	( 16'sd 26773) * $signed(input_fmap_116[7:0]) +
	( 13'sd 3245) * $signed(input_fmap_117[7:0]) +
	( 11'sd 866) * $signed(input_fmap_118[7:0]) +
	( 16'sd 19350) * $signed(input_fmap_119[7:0]) +
	( 14'sd 4543) * $signed(input_fmap_120[7:0]) +
	( 16'sd 19211) * $signed(input_fmap_121[7:0]) +
	( 15'sd 15757) * $signed(input_fmap_122[7:0]) +
	( 16'sd 27641) * $signed(input_fmap_123[7:0]) +
	( 15'sd 12196) * $signed(input_fmap_124[7:0]) +
	( 13'sd 2096) * $signed(input_fmap_125[7:0]) +
	( 16'sd 20122) * $signed(input_fmap_126[7:0]) +
	( 14'sd 7196) * $signed(input_fmap_127[7:0]) +
	( 15'sd 13258) * $signed(input_fmap_128[7:0]) +
	( 14'sd 5916) * $signed(input_fmap_129[7:0]) +
	( 15'sd 14830) * $signed(input_fmap_130[7:0]) +
	( 16'sd 17813) * $signed(input_fmap_131[7:0]) +
	( 16'sd 16423) * $signed(input_fmap_132[7:0]) +
	( 14'sd 7704) * $signed(input_fmap_133[7:0]) +
	( 16'sd 32050) * $signed(input_fmap_134[7:0]) +
	( 16'sd 17324) * $signed(input_fmap_135[7:0]) +
	( 15'sd 8496) * $signed(input_fmap_136[7:0]) +
	( 16'sd 27822) * $signed(input_fmap_137[7:0]) +
	( 15'sd 13678) * $signed(input_fmap_138[7:0]) +
	( 14'sd 4329) * $signed(input_fmap_139[7:0]) +
	( 15'sd 9528) * $signed(input_fmap_140[7:0]) +
	( 16'sd 16512) * $signed(input_fmap_141[7:0]) +
	( 16'sd 25698) * $signed(input_fmap_142[7:0]) +
	( 15'sd 9609) * $signed(input_fmap_143[7:0]) +
	( 15'sd 12822) * $signed(input_fmap_144[7:0]) +
	( 16'sd 30217) * $signed(input_fmap_145[7:0]) +
	( 16'sd 29755) * $signed(input_fmap_146[7:0]) +
	( 15'sd 13580) * $signed(input_fmap_147[7:0]) +
	( 15'sd 15797) * $signed(input_fmap_148[7:0]) +
	( 16'sd 26547) * $signed(input_fmap_149[7:0]) +
	( 16'sd 17172) * $signed(input_fmap_150[7:0]) +
	( 16'sd 17381) * $signed(input_fmap_151[7:0]) +
	( 15'sd 8309) * $signed(input_fmap_152[7:0]) +
	( 16'sd 28338) * $signed(input_fmap_153[7:0]) +
	( 14'sd 6736) * $signed(input_fmap_154[7:0]) +
	( 11'sd 922) * $signed(input_fmap_155[7:0]) +
	( 16'sd 20760) * $signed(input_fmap_156[7:0]) +
	( 15'sd 15545) * $signed(input_fmap_157[7:0]) +
	( 14'sd 4145) * $signed(input_fmap_158[7:0]) +
	( 15'sd 8565) * $signed(input_fmap_159[7:0]) +
	( 16'sd 32015) * $signed(input_fmap_160[7:0]) +
	( 15'sd 9479) * $signed(input_fmap_161[7:0]) +
	( 16'sd 21330) * $signed(input_fmap_162[7:0]) +
	( 14'sd 6288) * $signed(input_fmap_163[7:0]) +
	( 15'sd 12205) * $signed(input_fmap_164[7:0]) +
	( 14'sd 5186) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18254) * $signed(input_fmap_166[7:0]) +
	( 16'sd 17932) * $signed(input_fmap_167[7:0]) +
	( 14'sd 7623) * $signed(input_fmap_168[7:0]) +
	( 16'sd 26690) * $signed(input_fmap_169[7:0]) +
	( 16'sd 18271) * $signed(input_fmap_170[7:0]) +
	( 16'sd 23092) * $signed(input_fmap_171[7:0]) +
	( 16'sd 17473) * $signed(input_fmap_172[7:0]) +
	( 15'sd 13491) * $signed(input_fmap_173[7:0]) +
	( 16'sd 16557) * $signed(input_fmap_174[7:0]) +
	( 15'sd 8759) * $signed(input_fmap_175[7:0]) +
	( 16'sd 30688) * $signed(input_fmap_176[7:0]) +
	( 16'sd 30177) * $signed(input_fmap_177[7:0]) +
	( 11'sd 942) * $signed(input_fmap_178[7:0]) +
	( 16'sd 25055) * $signed(input_fmap_179[7:0]) +
	( 15'sd 8297) * $signed(input_fmap_180[7:0]) +
	( 12'sd 1208) * $signed(input_fmap_181[7:0]) +
	( 16'sd 18416) * $signed(input_fmap_182[7:0]) +
	( 13'sd 2441) * $signed(input_fmap_183[7:0]) +
	( 13'sd 2686) * $signed(input_fmap_184[7:0]) +
	( 13'sd 2799) * $signed(input_fmap_185[7:0]) +
	( 14'sd 4392) * $signed(input_fmap_186[7:0]) +
	( 15'sd 13139) * $signed(input_fmap_187[7:0]) +
	( 16'sd 17594) * $signed(input_fmap_188[7:0]) +
	( 14'sd 7199) * $signed(input_fmap_189[7:0]) +
	( 15'sd 15146) * $signed(input_fmap_190[7:0]) +
	( 16'sd 31668) * $signed(input_fmap_191[7:0]) +
	( 12'sd 1300) * $signed(input_fmap_192[7:0]) +
	( 16'sd 17275) * $signed(input_fmap_193[7:0]) +
	( 14'sd 4176) * $signed(input_fmap_194[7:0]) +
	( 16'sd 22385) * $signed(input_fmap_195[7:0]) +
	( 15'sd 12897) * $signed(input_fmap_196[7:0]) +
	( 16'sd 29710) * $signed(input_fmap_197[7:0]) +
	( 15'sd 13212) * $signed(input_fmap_198[7:0]) +
	( 15'sd 15669) * $signed(input_fmap_199[7:0]) +
	( 16'sd 30097) * $signed(input_fmap_200[7:0]) +
	( 16'sd 26492) * $signed(input_fmap_201[7:0]) +
	( 13'sd 2752) * $signed(input_fmap_202[7:0]) +
	( 16'sd 23631) * $signed(input_fmap_203[7:0]) +
	( 16'sd 30290) * $signed(input_fmap_204[7:0]) +
	( 16'sd 29681) * $signed(input_fmap_205[7:0]) +
	( 16'sd 21250) * $signed(input_fmap_206[7:0]) +
	( 12'sd 1808) * $signed(input_fmap_207[7:0]) +
	( 15'sd 14165) * $signed(input_fmap_208[7:0]) +
	( 12'sd 1886) * $signed(input_fmap_209[7:0]) +
	( 16'sd 23461) * $signed(input_fmap_210[7:0]) +
	( 16'sd 30926) * $signed(input_fmap_211[7:0]) +
	( 16'sd 17235) * $signed(input_fmap_212[7:0]) +
	( 14'sd 7533) * $signed(input_fmap_213[7:0]) +
	( 14'sd 7340) * $signed(input_fmap_214[7:0]) +
	( 15'sd 9138) * $signed(input_fmap_215[7:0]) +
	( 14'sd 7293) * $signed(input_fmap_216[7:0]) +
	( 8'sd 76) * $signed(input_fmap_217[7:0]) +
	( 14'sd 4220) * $signed(input_fmap_218[7:0]) +
	( 15'sd 15850) * $signed(input_fmap_219[7:0]) +
	( 14'sd 6488) * $signed(input_fmap_220[7:0]) +
	( 16'sd 19417) * $signed(input_fmap_221[7:0]) +
	( 12'sd 1829) * $signed(input_fmap_222[7:0]) +
	( 14'sd 8046) * $signed(input_fmap_223[7:0]) +
	( 16'sd 16430) * $signed(input_fmap_224[7:0]) +
	( 16'sd 24799) * $signed(input_fmap_225[7:0]) +
	( 14'sd 4246) * $signed(input_fmap_226[7:0]) +
	( 15'sd 11519) * $signed(input_fmap_227[7:0]) +
	( 10'sd 454) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20774) * $signed(input_fmap_229[7:0]) +
	( 15'sd 9994) * $signed(input_fmap_230[7:0]) +
	( 16'sd 25647) * $signed(input_fmap_231[7:0]) +
	( 16'sd 20932) * $signed(input_fmap_232[7:0]) +
	( 16'sd 21014) * $signed(input_fmap_233[7:0]) +
	( 15'sd 14571) * $signed(input_fmap_234[7:0]) +
	( 12'sd 1787) * $signed(input_fmap_235[7:0]) +
	( 15'sd 13007) * $signed(input_fmap_236[7:0]) +
	( 16'sd 28945) * $signed(input_fmap_237[7:0]) +
	( 16'sd 22571) * $signed(input_fmap_238[7:0]) +
	( 16'sd 25402) * $signed(input_fmap_239[7:0]) +
	( 15'sd 8699) * $signed(input_fmap_240[7:0]) +
	( 14'sd 7055) * $signed(input_fmap_241[7:0]) +
	( 16'sd 23579) * $signed(input_fmap_242[7:0]) +
	( 13'sd 2924) * $signed(input_fmap_243[7:0]) +
	( 16'sd 26538) * $signed(input_fmap_244[7:0]) +
	( 16'sd 29741) * $signed(input_fmap_245[7:0]) +
	( 16'sd 22695) * $signed(input_fmap_246[7:0]) +
	( 15'sd 12336) * $signed(input_fmap_247[7:0]) +
	( 15'sd 9410) * $signed(input_fmap_248[7:0]) +
	( 16'sd 31784) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7202) * $signed(input_fmap_250[7:0]) +
	( 15'sd 8908) * $signed(input_fmap_251[7:0]) +
	( 16'sd 24307) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13127) * $signed(input_fmap_253[7:0]) +
	( 16'sd 21868) * $signed(input_fmap_254[7:0]) +
	( 16'sd 29624) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_254;
assign conv_mac_254 = 
	( 16'sd 31923) * $signed(input_fmap_0[7:0]) +
	( 16'sd 32356) * $signed(input_fmap_1[7:0]) +
	( 16'sd 18858) * $signed(input_fmap_2[7:0]) +
	( 16'sd 25957) * $signed(input_fmap_3[7:0]) +
	( 16'sd 32584) * $signed(input_fmap_4[7:0]) +
	( 15'sd 12200) * $signed(input_fmap_5[7:0]) +
	( 16'sd 24513) * $signed(input_fmap_6[7:0]) +
	( 16'sd 22837) * $signed(input_fmap_7[7:0]) +
	( 15'sd 9868) * $signed(input_fmap_8[7:0]) +
	( 14'sd 7801) * $signed(input_fmap_9[7:0]) +
	( 13'sd 3740) * $signed(input_fmap_10[7:0]) +
	( 16'sd 26409) * $signed(input_fmap_11[7:0]) +
	( 15'sd 12227) * $signed(input_fmap_12[7:0]) +
	( 15'sd 11524) * $signed(input_fmap_13[7:0]) +
	( 16'sd 27420) * $signed(input_fmap_14[7:0]) +
	( 11'sd 977) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23705) * $signed(input_fmap_16[7:0]) +
	( 16'sd 19710) * $signed(input_fmap_17[7:0]) +
	( 14'sd 6139) * $signed(input_fmap_18[7:0]) +
	( 15'sd 13954) * $signed(input_fmap_19[7:0]) +
	( 16'sd 22663) * $signed(input_fmap_20[7:0]) +
	( 15'sd 12888) * $signed(input_fmap_21[7:0]) +
	( 16'sd 18360) * $signed(input_fmap_22[7:0]) +
	( 14'sd 4193) * $signed(input_fmap_23[7:0]) +
	( 16'sd 27639) * $signed(input_fmap_24[7:0]) +
	( 16'sd 20858) * $signed(input_fmap_25[7:0]) +
	( 16'sd 22110) * $signed(input_fmap_26[7:0]) +
	( 15'sd 8272) * $signed(input_fmap_27[7:0]) +
	( 16'sd 26096) * $signed(input_fmap_28[7:0]) +
	( 16'sd 18455) * $signed(input_fmap_29[7:0]) +
	( 16'sd 22601) * $signed(input_fmap_30[7:0]) +
	( 14'sd 4663) * $signed(input_fmap_31[7:0]) +
	( 12'sd 1992) * $signed(input_fmap_32[7:0]) +
	( 15'sd 13508) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5705) * $signed(input_fmap_34[7:0]) +
	( 12'sd 1834) * $signed(input_fmap_35[7:0]) +
	( 12'sd 1782) * $signed(input_fmap_36[7:0]) +
	( 16'sd 26170) * $signed(input_fmap_37[7:0]) +
	( 16'sd 25652) * $signed(input_fmap_38[7:0]) +
	( 16'sd 28445) * $signed(input_fmap_39[7:0]) +
	( 16'sd 25355) * $signed(input_fmap_40[7:0]) +
	( 10'sd 473) * $signed(input_fmap_41[7:0]) +
	( 13'sd 3235) * $signed(input_fmap_42[7:0]) +
	( 14'sd 8091) * $signed(input_fmap_43[7:0]) +
	( 14'sd 6793) * $signed(input_fmap_44[7:0]) +
	( 15'sd 16012) * $signed(input_fmap_45[7:0]) +
	( 16'sd 22308) * $signed(input_fmap_46[7:0]) +
	( 16'sd 22020) * $signed(input_fmap_47[7:0]) +
	( 16'sd 24185) * $signed(input_fmap_48[7:0]) +
	( 15'sd 8714) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9470) * $signed(input_fmap_50[7:0]) +
	( 13'sd 2619) * $signed(input_fmap_51[7:0]) +
	( 16'sd 20495) * $signed(input_fmap_52[7:0]) +
	( 15'sd 16103) * $signed(input_fmap_53[7:0]) +
	( 16'sd 27713) * $signed(input_fmap_54[7:0]) +
	( 15'sd 11751) * $signed(input_fmap_55[7:0]) +
	( 15'sd 12508) * $signed(input_fmap_56[7:0]) +
	( 13'sd 2705) * $signed(input_fmap_57[7:0]) +
	( 14'sd 4646) * $signed(input_fmap_58[7:0]) +
	( 16'sd 19374) * $signed(input_fmap_59[7:0]) +
	( 12'sd 1368) * $signed(input_fmap_60[7:0]) +
	( 16'sd 25745) * $signed(input_fmap_61[7:0]) +
	( 16'sd 31718) * $signed(input_fmap_62[7:0]) +
	( 16'sd 21936) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15946) * $signed(input_fmap_64[7:0]) +
	( 12'sd 1427) * $signed(input_fmap_65[7:0]) +
	( 16'sd 17524) * $signed(input_fmap_66[7:0]) +
	( 15'sd 10631) * $signed(input_fmap_67[7:0]) +
	( 15'sd 13686) * $signed(input_fmap_68[7:0]) +
	( 16'sd 30305) * $signed(input_fmap_69[7:0]) +
	( 16'sd 24562) * $signed(input_fmap_70[7:0]) +
	( 14'sd 6486) * $signed(input_fmap_71[7:0]) +
	( 16'sd 31144) * $signed(input_fmap_72[7:0]) +
	( 16'sd 29078) * $signed(input_fmap_73[7:0]) +
	( 15'sd 10758) * $signed(input_fmap_74[7:0]) +
	( 14'sd 4659) * $signed(input_fmap_75[7:0]) +
	( 16'sd 29102) * $signed(input_fmap_76[7:0]) +
	( 15'sd 10498) * $signed(input_fmap_77[7:0]) +
	( 15'sd 9584) * $signed(input_fmap_78[7:0]) +
	( 16'sd 27239) * $signed(input_fmap_79[7:0]) +
	( 16'sd 19225) * $signed(input_fmap_80[7:0]) +
	( 13'sd 2787) * $signed(input_fmap_81[7:0]) +
	( 16'sd 32036) * $signed(input_fmap_82[7:0]) +
	( 14'sd 6626) * $signed(input_fmap_83[7:0]) +
	( 14'sd 5113) * $signed(input_fmap_84[7:0]) +
	( 14'sd 6563) * $signed(input_fmap_85[7:0]) +
	( 13'sd 3027) * $signed(input_fmap_86[7:0]) +
	( 16'sd 31725) * $signed(input_fmap_87[7:0]) +
	( 16'sd 27995) * $signed(input_fmap_88[7:0]) +
	( 16'sd 32463) * $signed(input_fmap_89[7:0]) +
	( 14'sd 8136) * $signed(input_fmap_90[7:0]) +
	( 16'sd 24766) * $signed(input_fmap_91[7:0]) +
	( 14'sd 6109) * $signed(input_fmap_92[7:0]) +
	( 15'sd 11385) * $signed(input_fmap_93[7:0]) +
	( 14'sd 7441) * $signed(input_fmap_94[7:0]) +
	( 14'sd 5337) * $signed(input_fmap_95[7:0]) +
	( 16'sd 24200) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11113) * $signed(input_fmap_97[7:0]) +
	( 15'sd 9566) * $signed(input_fmap_98[7:0]) +
	( 14'sd 7519) * $signed(input_fmap_99[7:0]) +
	( 16'sd 32572) * $signed(input_fmap_100[7:0]) +
	( 16'sd 24128) * $signed(input_fmap_101[7:0]) +
	( 13'sd 3355) * $signed(input_fmap_102[7:0]) +
	( 15'sd 11273) * $signed(input_fmap_103[7:0]) +
	( 16'sd 17740) * $signed(input_fmap_104[7:0]) +
	( 14'sd 6901) * $signed(input_fmap_105[7:0]) +
	( 15'sd 11462) * $signed(input_fmap_106[7:0]) +
	( 16'sd 25552) * $signed(input_fmap_107[7:0]) +
	( 15'sd 8381) * $signed(input_fmap_108[7:0]) +
	( 15'sd 16332) * $signed(input_fmap_109[7:0]) +
	( 15'sd 11979) * $signed(input_fmap_110[7:0]) +
	( 15'sd 15592) * $signed(input_fmap_111[7:0]) +
	( 10'sd 293) * $signed(input_fmap_112[7:0]) +
	( 16'sd 17460) * $signed(input_fmap_113[7:0]) +
	( 15'sd 16298) * $signed(input_fmap_114[7:0]) +
	( 12'sd 1709) * $signed(input_fmap_115[7:0]) +
	( 16'sd 18076) * $signed(input_fmap_116[7:0]) +
	( 16'sd 19273) * $signed(input_fmap_117[7:0]) +
	( 16'sd 18990) * $signed(input_fmap_118[7:0]) +
	( 15'sd 15758) * $signed(input_fmap_119[7:0]) +
	( 14'sd 8168) * $signed(input_fmap_120[7:0]) +
	( 16'sd 17655) * $signed(input_fmap_121[7:0]) +
	( 16'sd 19370) * $signed(input_fmap_122[7:0]) +
	( 3'sd 3) * $signed(input_fmap_123[7:0]) +
	( 16'sd 27460) * $signed(input_fmap_124[7:0]) +
	( 16'sd 30646) * $signed(input_fmap_125[7:0]) +
	( 16'sd 27430) * $signed(input_fmap_126[7:0]) +
	( 15'sd 10400) * $signed(input_fmap_127[7:0]) +
	( 16'sd 27462) * $signed(input_fmap_128[7:0]) +
	( 15'sd 15031) * $signed(input_fmap_129[7:0]) +
	( 15'sd 10564) * $signed(input_fmap_130[7:0]) +
	( 16'sd 32710) * $signed(input_fmap_131[7:0]) +
	( 16'sd 20772) * $signed(input_fmap_132[7:0]) +
	( 14'sd 6719) * $signed(input_fmap_133[7:0]) +
	( 15'sd 11452) * $signed(input_fmap_134[7:0]) +
	( 16'sd 30825) * $signed(input_fmap_135[7:0]) +
	( 16'sd 21051) * $signed(input_fmap_136[7:0]) +
	( 15'sd 11689) * $signed(input_fmap_137[7:0]) +
	( 13'sd 2165) * $signed(input_fmap_138[7:0]) +
	( 15'sd 14527) * $signed(input_fmap_139[7:0]) +
	( 16'sd 24601) * $signed(input_fmap_140[7:0]) +
	( 13'sd 3397) * $signed(input_fmap_141[7:0]) +
	( 10'sd 355) * $signed(input_fmap_142[7:0]) +
	( 16'sd 20689) * $signed(input_fmap_143[7:0]) +
	( 15'sd 9875) * $signed(input_fmap_144[7:0]) +
	( 16'sd 22940) * $signed(input_fmap_145[7:0]) +
	( 14'sd 4153) * $signed(input_fmap_146[7:0]) +
	( 16'sd 28239) * $signed(input_fmap_147[7:0]) +
	( 16'sd 31293) * $signed(input_fmap_148[7:0]) +
	( 16'sd 26274) * $signed(input_fmap_149[7:0]) +
	( 10'sd 493) * $signed(input_fmap_150[7:0]) +
	( 11'sd 583) * $signed(input_fmap_151[7:0]) +
	( 14'sd 5488) * $signed(input_fmap_152[7:0]) +
	( 14'sd 7244) * $signed(input_fmap_153[7:0]) +
	( 16'sd 26658) * $signed(input_fmap_154[7:0]) +
	( 15'sd 11643) * $signed(input_fmap_155[7:0]) +
	( 14'sd 6777) * $signed(input_fmap_156[7:0]) +
	( 16'sd 30899) * $signed(input_fmap_157[7:0]) +
	( 15'sd 10475) * $signed(input_fmap_158[7:0]) +
	( 16'sd 32181) * $signed(input_fmap_159[7:0]) +
	( 16'sd 23465) * $signed(input_fmap_160[7:0]) +
	( 16'sd 26331) * $signed(input_fmap_161[7:0]) +
	( 16'sd 25302) * $signed(input_fmap_162[7:0]) +
	( 16'sd 22365) * $signed(input_fmap_163[7:0]) +
	( 15'sd 9409) * $signed(input_fmap_164[7:0]) +
	( 16'sd 28721) * $signed(input_fmap_165[7:0]) +
	( 16'sd 18702) * $signed(input_fmap_166[7:0]) +
	( 15'sd 13025) * $signed(input_fmap_167[7:0]) +
	( 12'sd 1945) * $signed(input_fmap_168[7:0]) +
	( 16'sd 30674) * $signed(input_fmap_169[7:0]) +
	( 16'sd 29517) * $signed(input_fmap_170[7:0]) +
	( 16'sd 31994) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19987) * $signed(input_fmap_172[7:0]) +
	( 16'sd 29691) * $signed(input_fmap_173[7:0]) +
	( 15'sd 14663) * $signed(input_fmap_174[7:0]) +
	( 16'sd 18650) * $signed(input_fmap_175[7:0]) +
	( 13'sd 2158) * $signed(input_fmap_176[7:0]) +
	( 13'sd 3165) * $signed(input_fmap_177[7:0]) +
	( 15'sd 11429) * $signed(input_fmap_178[7:0]) +
	( 14'sd 6124) * $signed(input_fmap_179[7:0]) +
	( 16'sd 32479) * $signed(input_fmap_180[7:0]) +
	( 16'sd 21667) * $signed(input_fmap_181[7:0]) +
	( 16'sd 26726) * $signed(input_fmap_182[7:0]) +
	( 16'sd 28849) * $signed(input_fmap_183[7:0]) +
	( 16'sd 24925) * $signed(input_fmap_184[7:0]) +
	( 13'sd 3450) * $signed(input_fmap_185[7:0]) +
	( 15'sd 12251) * $signed(input_fmap_186[7:0]) +
	( 15'sd 14433) * $signed(input_fmap_187[7:0]) +
	( 16'sd 25815) * $signed(input_fmap_188[7:0]) +
	( 16'sd 17590) * $signed(input_fmap_189[7:0]) +
	( 16'sd 32713) * $signed(input_fmap_190[7:0]) +
	( 16'sd 20640) * $signed(input_fmap_191[7:0]) +
	( 16'sd 32076) * $signed(input_fmap_192[7:0]) +
	( 16'sd 22323) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3781) * $signed(input_fmap_194[7:0]) +
	( 16'sd 27856) * $signed(input_fmap_195[7:0]) +
	( 16'sd 19613) * $signed(input_fmap_196[7:0]) +
	( 16'sd 30367) * $signed(input_fmap_197[7:0]) +
	( 14'sd 5902) * $signed(input_fmap_198[7:0]) +
	( 16'sd 21779) * $signed(input_fmap_199[7:0]) +
	( 16'sd 21816) * $signed(input_fmap_200[7:0]) +
	( 15'sd 15256) * $signed(input_fmap_201[7:0]) +
	( 16'sd 25988) * $signed(input_fmap_202[7:0]) +
	( 13'sd 2307) * $signed(input_fmap_203[7:0]) +
	( 14'sd 6161) * $signed(input_fmap_204[7:0]) +
	( 16'sd 18535) * $signed(input_fmap_205[7:0]) +
	( 16'sd 17451) * $signed(input_fmap_206[7:0]) +
	( 14'sd 7573) * $signed(input_fmap_207[7:0]) +
	( 16'sd 18461) * $signed(input_fmap_208[7:0]) +
	( 15'sd 12709) * $signed(input_fmap_209[7:0]) +
	( 15'sd 10093) * $signed(input_fmap_210[7:0]) +
	( 16'sd 25420) * $signed(input_fmap_211[7:0]) +
	( 15'sd 9764) * $signed(input_fmap_212[7:0]) +
	( 16'sd 28106) * $signed(input_fmap_213[7:0]) +
	( 15'sd 16326) * $signed(input_fmap_214[7:0]) +
	( 16'sd 28796) * $signed(input_fmap_215[7:0]) +
	( 15'sd 8722) * $signed(input_fmap_216[7:0]) +
	( 15'sd 14602) * $signed(input_fmap_217[7:0]) +
	( 16'sd 18070) * $signed(input_fmap_218[7:0]) +
	( 16'sd 19503) * $signed(input_fmap_219[7:0]) +
	( 15'sd 10577) * $signed(input_fmap_220[7:0]) +
	( 16'sd 25643) * $signed(input_fmap_221[7:0]) +
	( 16'sd 18368) * $signed(input_fmap_222[7:0]) +
	( 11'sd 714) * $signed(input_fmap_223[7:0]) +
	( 16'sd 29000) * $signed(input_fmap_224[7:0]) +
	( 14'sd 7015) * $signed(input_fmap_225[7:0]) +
	( 16'sd 24233) * $signed(input_fmap_226[7:0]) +
	( 10'sd 471) * $signed(input_fmap_227[7:0]) +
	( 15'sd 10447) * $signed(input_fmap_228[7:0]) +
	( 16'sd 20211) * $signed(input_fmap_229[7:0]) +
	( 11'sd 996) * $signed(input_fmap_230[7:0]) +
	( 15'sd 11334) * $signed(input_fmap_231[7:0]) +
	( 16'sd 28106) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3249) * $signed(input_fmap_233[7:0]) +
	( 16'sd 23005) * $signed(input_fmap_234[7:0]) +
	( 16'sd 24311) * $signed(input_fmap_235[7:0]) +
	( 16'sd 26960) * $signed(input_fmap_236[7:0]) +
	( 16'sd 17756) * $signed(input_fmap_237[7:0]) +
	( 11'sd 822) * $signed(input_fmap_238[7:0]) +
	( 14'sd 7549) * $signed(input_fmap_239[7:0]) +
	( 12'sd 1328) * $signed(input_fmap_240[7:0]) +
	( 14'sd 5446) * $signed(input_fmap_241[7:0]) +
	( 16'sd 27752) * $signed(input_fmap_242[7:0]) +
	( 16'sd 25285) * $signed(input_fmap_243[7:0]) +
	( 16'sd 21614) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24074) * $signed(input_fmap_245[7:0]) +
	( 16'sd 17455) * $signed(input_fmap_246[7:0]) +
	( 12'sd 1365) * $signed(input_fmap_247[7:0]) +
	( 16'sd 31970) * $signed(input_fmap_248[7:0]) +
	( 16'sd 28700) * $signed(input_fmap_249[7:0]) +
	( 14'sd 7854) * $signed(input_fmap_250[7:0]) +
	( 14'sd 4109) * $signed(input_fmap_251[7:0]) +
	( 16'sd 32350) * $signed(input_fmap_252[7:0]) +
	( 15'sd 13244) * $signed(input_fmap_253[7:0]) +
	( 16'sd 26620) * $signed(input_fmap_254[7:0]) +
	( 15'sd 12823) * $signed(input_fmap_255[7:0]);

logic signed [31:0] conv_mac_255;
assign conv_mac_255 = 
	( 14'sd 6279) * $signed(input_fmap_0[7:0]) +
	( 16'sd 26201) * $signed(input_fmap_1[7:0]) +
	( 15'sd 12815) * $signed(input_fmap_2[7:0]) +
	( 15'sd 9694) * $signed(input_fmap_3[7:0]) +
	( 13'sd 3489) * $signed(input_fmap_4[7:0]) +
	( 12'sd 1519) * $signed(input_fmap_5[7:0]) +
	( 16'sd 22089) * $signed(input_fmap_6[7:0]) +
	( 16'sd 29437) * $signed(input_fmap_7[7:0]) +
	( 15'sd 13800) * $signed(input_fmap_8[7:0]) +
	( 14'sd 6686) * $signed(input_fmap_9[7:0]) +
	( 15'sd 12980) * $signed(input_fmap_10[7:0]) +
	( 15'sd 11476) * $signed(input_fmap_11[7:0]) +
	( 15'sd 15587) * $signed(input_fmap_12[7:0]) +
	( 12'sd 1609) * $signed(input_fmap_13[7:0]) +
	( 14'sd 7559) * $signed(input_fmap_14[7:0]) +
	( 13'sd 2845) * $signed(input_fmap_15[7:0]) +
	( 16'sd 23229) * $signed(input_fmap_16[7:0]) +
	( 16'sd 20737) * $signed(input_fmap_17[7:0]) +
	( 16'sd 32087) * $signed(input_fmap_18[7:0]) +
	( 14'sd 5967) * $signed(input_fmap_19[7:0]) +
	( 16'sd 31617) * $signed(input_fmap_20[7:0]) +
	( 14'sd 5549) * $signed(input_fmap_21[7:0]) +
	( 15'sd 9465) * $signed(input_fmap_22[7:0]) +
	( 16'sd 21323) * $signed(input_fmap_23[7:0]) +
	( 15'sd 14342) * $signed(input_fmap_24[7:0]) +
	( 15'sd 12690) * $signed(input_fmap_25[7:0]) +
	( 16'sd 20437) * $signed(input_fmap_26[7:0]) +
	( 15'sd 9813) * $signed(input_fmap_27[7:0]) +
	( 15'sd 14929) * $signed(input_fmap_28[7:0]) +
	( 16'sd 19362) * $signed(input_fmap_29[7:0]) +
	( 13'sd 2669) * $signed(input_fmap_30[7:0]) +
	( 16'sd 18119) * $signed(input_fmap_31[7:0]) +
	( 16'sd 18177) * $signed(input_fmap_32[7:0]) +
	( 13'sd 2541) * $signed(input_fmap_33[7:0]) +
	( 14'sd 5323) * $signed(input_fmap_34[7:0]) +
	( 16'sd 20922) * $signed(input_fmap_35[7:0]) +
	( 13'sd 4015) * $signed(input_fmap_36[7:0]) +
	( 16'sd 24990) * $signed(input_fmap_37[7:0]) +
	( 15'sd 11975) * $signed(input_fmap_38[7:0]) +
	( 15'sd 8975) * $signed(input_fmap_39[7:0]) +
	( 15'sd 8907) * $signed(input_fmap_40[7:0]) +
	( 16'sd 25842) * $signed(input_fmap_41[7:0]) +
	( 16'sd 16592) * $signed(input_fmap_42[7:0]) +
	( 16'sd 26769) * $signed(input_fmap_43[7:0]) +
	( 16'sd 17646) * $signed(input_fmap_44[7:0]) +
	( 16'sd 29153) * $signed(input_fmap_45[7:0]) +
	( 14'sd 7612) * $signed(input_fmap_46[7:0]) +
	( 14'sd 8096) * $signed(input_fmap_47[7:0]) +
	( 15'sd 8919) * $signed(input_fmap_48[7:0]) +
	( 12'sd 2038) * $signed(input_fmap_49[7:0]) +
	( 15'sd 9652) * $signed(input_fmap_50[7:0]) +
	( 16'sd 23302) * $signed(input_fmap_51[7:0]) +
	( 11'sd 528) * $signed(input_fmap_52[7:0]) +
	( 14'sd 5696) * $signed(input_fmap_53[7:0]) +
	( 16'sd 16418) * $signed(input_fmap_54[7:0]) +
	( 14'sd 4702) * $signed(input_fmap_55[7:0]) +
	( 16'sd 20092) * $signed(input_fmap_56[7:0]) +
	( 15'sd 10560) * $signed(input_fmap_57[7:0]) +
	( 16'sd 17536) * $signed(input_fmap_58[7:0]) +
	( 16'sd 21986) * $signed(input_fmap_59[7:0]) +
	( 14'sd 5548) * $signed(input_fmap_60[7:0]) +
	( 14'sd 4991) * $signed(input_fmap_61[7:0]) +
	( 16'sd 16504) * $signed(input_fmap_62[7:0]) +
	( 16'sd 23336) * $signed(input_fmap_63[7:0]) +
	( 15'sd 15633) * $signed(input_fmap_64[7:0]) +
	( 13'sd 2618) * $signed(input_fmap_65[7:0]) +
	( 16'sd 30396) * $signed(input_fmap_66[7:0]) +
	( 15'sd 13818) * $signed(input_fmap_67[7:0]) +
	( 14'sd 5669) * $signed(input_fmap_68[7:0]) +
	( 15'sd 14804) * $signed(input_fmap_69[7:0]) +
	( 16'sd 20944) * $signed(input_fmap_70[7:0]) +
	( 11'sd 680) * $signed(input_fmap_71[7:0]) +
	( 16'sd 20289) * $signed(input_fmap_72[7:0]) +
	( 15'sd 11089) * $signed(input_fmap_73[7:0]) +
	( 15'sd 8572) * $signed(input_fmap_74[7:0]) +
	( 16'sd 32448) * $signed(input_fmap_75[7:0]) +
	( 15'sd 9625) * $signed(input_fmap_76[7:0]) +
	( 16'sd 17682) * $signed(input_fmap_77[7:0]) +
	( 16'sd 29114) * $signed(input_fmap_78[7:0]) +
	( 15'sd 10863) * $signed(input_fmap_79[7:0]) +
	( 15'sd 15609) * $signed(input_fmap_80[7:0]) +
	( 15'sd 10274) * $signed(input_fmap_81[7:0]) +
	( 16'sd 27084) * $signed(input_fmap_82[7:0]) +
	( 15'sd 8825) * $signed(input_fmap_83[7:0]) +
	( 15'sd 15093) * $signed(input_fmap_84[7:0]) +
	( 16'sd 21581) * $signed(input_fmap_85[7:0]) +
	( 16'sd 20336) * $signed(input_fmap_86[7:0]) +
	( 16'sd 16442) * $signed(input_fmap_87[7:0]) +
	( 14'sd 5558) * $signed(input_fmap_88[7:0]) +
	( 16'sd 27359) * $signed(input_fmap_89[7:0]) +
	( 13'sd 4081) * $signed(input_fmap_90[7:0]) +
	( 16'sd 27114) * $signed(input_fmap_91[7:0]) +
	( 14'sd 5934) * $signed(input_fmap_92[7:0]) +
	( 13'sd 3429) * $signed(input_fmap_93[7:0]) +
	( 16'sd 28629) * $signed(input_fmap_94[7:0]) +
	( 16'sd 24927) * $signed(input_fmap_95[7:0]) +
	( 15'sd 10718) * $signed(input_fmap_96[7:0]) +
	( 15'sd 11063) * $signed(input_fmap_97[7:0]) +
	( 16'sd 17220) * $signed(input_fmap_98[7:0]) +
	( 16'sd 29555) * $signed(input_fmap_99[7:0]) +
	( 15'sd 11695) * $signed(input_fmap_100[7:0]) +
	( 16'sd 16421) * $signed(input_fmap_101[7:0]) +
	( 16'sd 20127) * $signed(input_fmap_102[7:0]) +
	( 16'sd 19267) * $signed(input_fmap_103[7:0]) +
	( 16'sd 27390) * $signed(input_fmap_104[7:0]) +
	( 15'sd 15696) * $signed(input_fmap_105[7:0]) +
	( 12'sd 1798) * $signed(input_fmap_106[7:0]) +
	( 16'sd 26320) * $signed(input_fmap_107[7:0]) +
	( 13'sd 2521) * $signed(input_fmap_108[7:0]) +
	( 14'sd 6699) * $signed(input_fmap_109[7:0]) +
	( 14'sd 7438) * $signed(input_fmap_110[7:0]) +
	( 15'sd 16057) * $signed(input_fmap_111[7:0]) +
	( 16'sd 30347) * $signed(input_fmap_112[7:0]) +
	( 14'sd 4357) * $signed(input_fmap_113[7:0]) +
	( 16'sd 26138) * $signed(input_fmap_114[7:0]) +
	( 11'sd 862) * $signed(input_fmap_115[7:0]) +
	( 16'sd 29408) * $signed(input_fmap_116[7:0]) +
	( 16'sd 22299) * $signed(input_fmap_117[7:0]) +
	( 16'sd 27242) * $signed(input_fmap_118[7:0]) +
	( 16'sd 17561) * $signed(input_fmap_119[7:0]) +
	( 15'sd 11981) * $signed(input_fmap_120[7:0]) +
	( 15'sd 14784) * $signed(input_fmap_121[7:0]) +
	( 15'sd 12451) * $signed(input_fmap_122[7:0]) +
	( 16'sd 20255) * $signed(input_fmap_123[7:0]) +
	( 16'sd 28687) * $signed(input_fmap_124[7:0]) +
	( 16'sd 26260) * $signed(input_fmap_125[7:0]) +
	( 16'sd 17217) * $signed(input_fmap_126[7:0]) +
	( 13'sd 2150) * $signed(input_fmap_127[7:0]) +
	( 16'sd 17628) * $signed(input_fmap_128[7:0]) +
	( 16'sd 31909) * $signed(input_fmap_129[7:0]) +
	( 16'sd 29084) * $signed(input_fmap_130[7:0]) +
	( 15'sd 15929) * $signed(input_fmap_131[7:0]) +
	( 14'sd 4393) * $signed(input_fmap_132[7:0]) +
	( 16'sd 25695) * $signed(input_fmap_133[7:0]) +
	( 16'sd 17649) * $signed(input_fmap_134[7:0]) +
	( 16'sd 17312) * $signed(input_fmap_135[7:0]) +
	( 10'sd 275) * $signed(input_fmap_136[7:0]) +
	( 16'sd 22340) * $signed(input_fmap_137[7:0]) +
	( 16'sd 31091) * $signed(input_fmap_138[7:0]) +
	( 16'sd 21997) * $signed(input_fmap_139[7:0]) +
	( 14'sd 8097) * $signed(input_fmap_140[7:0]) +
	( 13'sd 2908) * $signed(input_fmap_141[7:0]) +
	( 16'sd 19577) * $signed(input_fmap_142[7:0]) +
	( 16'sd 28372) * $signed(input_fmap_143[7:0]) +
	( 14'sd 5541) * $signed(input_fmap_144[7:0]) +
	( 16'sd 29568) * $signed(input_fmap_145[7:0]) +
	( 14'sd 6147) * $signed(input_fmap_146[7:0]) +
	( 16'sd 16946) * $signed(input_fmap_147[7:0]) +
	( 14'sd 7877) * $signed(input_fmap_148[7:0]) +
	( 16'sd 25207) * $signed(input_fmap_149[7:0]) +
	( 14'sd 7770) * $signed(input_fmap_150[7:0]) +
	( 16'sd 24591) * $signed(input_fmap_151[7:0]) +
	( 16'sd 32229) * $signed(input_fmap_152[7:0]) +
	( 16'sd 32731) * $signed(input_fmap_153[7:0]) +
	( 16'sd 31287) * $signed(input_fmap_154[7:0]) +
	( 15'sd 12195) * $signed(input_fmap_155[7:0]) +
	( 16'sd 22268) * $signed(input_fmap_156[7:0]) +
	( 16'sd 28467) * $signed(input_fmap_157[7:0]) +
	( 16'sd 23055) * $signed(input_fmap_158[7:0]) +
	( 14'sd 6551) * $signed(input_fmap_159[7:0]) +
	( 16'sd 27090) * $signed(input_fmap_160[7:0]) +
	( 16'sd 17451) * $signed(input_fmap_161[7:0]) +
	( 16'sd 19157) * $signed(input_fmap_162[7:0]) +
	( 16'sd 27549) * $signed(input_fmap_163[7:0]) +
	( 13'sd 3273) * $signed(input_fmap_164[7:0]) +
	( 14'sd 5668) * $signed(input_fmap_165[7:0]) +
	( 16'sd 31921) * $signed(input_fmap_166[7:0]) +
	( 16'sd 16403) * $signed(input_fmap_167[7:0]) +
	( 16'sd 32695) * $signed(input_fmap_168[7:0]) +
	( 16'sd 31522) * $signed(input_fmap_169[7:0]) +
	( 9'sd 158) * $signed(input_fmap_170[7:0]) +
	( 16'sd 16729) * $signed(input_fmap_171[7:0]) +
	( 16'sd 19873) * $signed(input_fmap_172[7:0]) +
	( 16'sd 23074) * $signed(input_fmap_173[7:0]) +
	( 13'sd 2750) * $signed(input_fmap_174[7:0]) +
	( 16'sd 21960) * $signed(input_fmap_175[7:0]) +
	( 16'sd 30786) * $signed(input_fmap_176[7:0]) +
	( 9'sd 140) * $signed(input_fmap_177[7:0]) +
	( 15'sd 11323) * $signed(input_fmap_178[7:0]) +
	( 16'sd 16529) * $signed(input_fmap_179[7:0]) +
	( 15'sd 9762) * $signed(input_fmap_180[7:0]) +
	( 15'sd 15227) * $signed(input_fmap_181[7:0]) +
	( 16'sd 22390) * $signed(input_fmap_182[7:0]) +
	( 16'sd 17790) * $signed(input_fmap_183[7:0]) +
	( 13'sd 3608) * $signed(input_fmap_184[7:0]) +
	( 16'sd 28826) * $signed(input_fmap_185[7:0]) +
	( 16'sd 22586) * $signed(input_fmap_186[7:0]) +
	( 14'sd 5588) * $signed(input_fmap_187[7:0]) +
	( 15'sd 14382) * $signed(input_fmap_188[7:0]) +
	( 16'sd 29972) * $signed(input_fmap_189[7:0]) +
	( 14'sd 5392) * $signed(input_fmap_190[7:0]) +
	( 13'sd 2436) * $signed(input_fmap_191[7:0]) +
	( 16'sd 19804) * $signed(input_fmap_192[7:0]) +
	( 16'sd 29813) * $signed(input_fmap_193[7:0]) +
	( 13'sd 3290) * $signed(input_fmap_194[7:0]) +
	( 15'sd 15184) * $signed(input_fmap_195[7:0]) +
	( 15'sd 10790) * $signed(input_fmap_196[7:0]) +
	( 16'sd 21870) * $signed(input_fmap_197[7:0]) +
	( 14'sd 8106) * $signed(input_fmap_198[7:0]) +
	( 16'sd 25961) * $signed(input_fmap_199[7:0]) +
	( 15'sd 11498) * $signed(input_fmap_200[7:0]) +
	( 13'sd 3927) * $signed(input_fmap_201[7:0]) +
	( 14'sd 7444) * $signed(input_fmap_202[7:0]) +
	( 16'sd 21105) * $signed(input_fmap_203[7:0]) +
	( 15'sd 14536) * $signed(input_fmap_204[7:0]) +
	( 16'sd 19973) * $signed(input_fmap_205[7:0]) +
	( 16'sd 28728) * $signed(input_fmap_206[7:0]) +
	( 16'sd 19275) * $signed(input_fmap_207[7:0]) +
	( 16'sd 31784) * $signed(input_fmap_208[7:0]) +
	( 13'sd 3734) * $signed(input_fmap_209[7:0]) +
	( 16'sd 20219) * $signed(input_fmap_210[7:0]) +
	( 16'sd 28937) * $signed(input_fmap_211[7:0]) +
	( 15'sd 10399) * $signed(input_fmap_212[7:0]) +
	( 12'sd 2016) * $signed(input_fmap_213[7:0]) +
	( 16'sd 31183) * $signed(input_fmap_214[7:0]) +
	( 14'sd 6347) * $signed(input_fmap_215[7:0]) +
	( 13'sd 2467) * $signed(input_fmap_216[7:0]) +
	( 15'sd 9646) * $signed(input_fmap_217[7:0]) +
	( 13'sd 2957) * $signed(input_fmap_218[7:0]) +
	( 16'sd 21377) * $signed(input_fmap_219[7:0]) +
	( 5'sd 9) * $signed(input_fmap_220[7:0]) +
	( 16'sd 16849) * $signed(input_fmap_221[7:0]) +
	( 16'sd 32739) * $signed(input_fmap_222[7:0]) +
	( 15'sd 12113) * $signed(input_fmap_223[7:0]) +
	( 14'sd 4526) * $signed(input_fmap_224[7:0]) +
	( 15'sd 15038) * $signed(input_fmap_225[7:0]) +
	( 14'sd 5076) * $signed(input_fmap_226[7:0]) +
	( 14'sd 5340) * $signed(input_fmap_227[7:0]) +
	( 14'sd 8188) * $signed(input_fmap_228[7:0]) +
	( 13'sd 3724) * $signed(input_fmap_229[7:0]) +
	( 16'sd 21825) * $signed(input_fmap_230[7:0]) +
	( 16'sd 17286) * $signed(input_fmap_231[7:0]) +
	( 16'sd 21119) * $signed(input_fmap_232[7:0]) +
	( 13'sd 3459) * $signed(input_fmap_233[7:0]) +
	( 15'sd 13524) * $signed(input_fmap_234[7:0]) +
	( 16'sd 29477) * $signed(input_fmap_235[7:0]) +
	( 14'sd 7208) * $signed(input_fmap_236[7:0]) +
	( 15'sd 11467) * $signed(input_fmap_237[7:0]) +
	( 15'sd 12472) * $signed(input_fmap_238[7:0]) +
	( 16'sd 23869) * $signed(input_fmap_239[7:0]) +
	( 11'sd 628) * $signed(input_fmap_240[7:0]) +
	( 16'sd 16471) * $signed(input_fmap_241[7:0]) +
	( 15'sd 15903) * $signed(input_fmap_242[7:0]) +
	( 16'sd 22029) * $signed(input_fmap_243[7:0]) +
	( 16'sd 30744) * $signed(input_fmap_244[7:0]) +
	( 16'sd 24081) * $signed(input_fmap_245[7:0]) +
	( 15'sd 9589) * $signed(input_fmap_246[7:0]) +
	( 16'sd 16688) * $signed(input_fmap_247[7:0]) +
	( 14'sd 6003) * $signed(input_fmap_248[7:0]) +
	( 16'sd 30328) * $signed(input_fmap_249[7:0]) +
	( 13'sd 2662) * $signed(input_fmap_250[7:0]) +
	( 14'sd 7282) * $signed(input_fmap_251[7:0]) +
	( 16'sd 26611) * $signed(input_fmap_252[7:0]) +
	( 16'sd 31923) * $signed(input_fmap_253[7:0]) +
	( 13'sd 4059) * $signed(input_fmap_254[7:0]) +
	( 14'sd 7988) * $signed(input_fmap_255[7:0]);

logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 16'd31567;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 12'd1907;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 11'd801;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 15'd12726;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 13'd2262;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 12'd1913;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 15'd11330;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 15'd8554;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 13'd2338;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 14'd7894;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 16'd24377;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 16'd27062;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 16'd22535;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 15'd14653;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 12'd1962;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 15'd14695;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 13'd2964;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 15'd13785;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 16'd30327;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 16'd22090;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 13'd2424;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 16'd30449;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 15'd9586;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 16'd24046;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 16'd17621;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 16'd22679;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 16'd23447;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 15'd10062;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 15'd10482;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 15'd8855;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 16'd29371;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 16'd32033;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 15'd13513;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 13'd3890;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 15'd10908;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 14'd5411;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 16'd25570;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 15'd10231;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 16'd29395;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 16'd21161;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 15'd15163;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 14'd7259;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 14'd4137;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 14'd4435;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 15'd11925;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 14'd5233;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 16'd31907;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 16'd24215;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 16'd26424;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 16'd19671;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 16'd21670;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 16'd32541;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 16'd30236;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 14'd4842;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 13'd3381;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 16'd23693;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 15'd11793;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 16'd30308;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 15'd15158;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 16'd29569;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 16'd27576;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 15'd15078;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 14'd5423;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 15'd14742;
logic [31:0] bias_add_64;
assign bias_add_64 = conv_mac_64 + 14'd4529;
logic [31:0] bias_add_65;
assign bias_add_65 = conv_mac_65 + 15'd8375;
logic [31:0] bias_add_66;
assign bias_add_66 = conv_mac_66 + 16'd21419;
logic [31:0] bias_add_67;
assign bias_add_67 = conv_mac_67 + 14'd7582;
logic [31:0] bias_add_68;
assign bias_add_68 = conv_mac_68 + 15'd10605;
logic [31:0] bias_add_69;
assign bias_add_69 = conv_mac_69 + 15'd11166;
logic [31:0] bias_add_70;
assign bias_add_70 = conv_mac_70 + 15'd10329;
logic [31:0] bias_add_71;
assign bias_add_71 = conv_mac_71 + 16'd18913;
logic [31:0] bias_add_72;
assign bias_add_72 = conv_mac_72 + 16'd19779;
logic [31:0] bias_add_73;
assign bias_add_73 = conv_mac_73 + 16'd24588;
logic [31:0] bias_add_74;
assign bias_add_74 = conv_mac_74 + 10'd485;
logic [31:0] bias_add_75;
assign bias_add_75 = conv_mac_75 + 16'd29266;
logic [31:0] bias_add_76;
assign bias_add_76 = conv_mac_76 + 16'd31766;
logic [31:0] bias_add_77;
assign bias_add_77 = conv_mac_77 + 16'd18963;
logic [31:0] bias_add_78;
assign bias_add_78 = conv_mac_78 + 16'd22140;
logic [31:0] bias_add_79;
assign bias_add_79 = conv_mac_79 + 9'd133;
logic [31:0] bias_add_80;
assign bias_add_80 = conv_mac_80 + 13'd3675;
logic [31:0] bias_add_81;
assign bias_add_81 = conv_mac_81 + 14'd6947;
logic [31:0] bias_add_82;
assign bias_add_82 = conv_mac_82 + 16'd20170;
logic [31:0] bias_add_83;
assign bias_add_83 = conv_mac_83 + 15'd8256;
logic [31:0] bias_add_84;
assign bias_add_84 = conv_mac_84 + 16'd24342;
logic [31:0] bias_add_85;
assign bias_add_85 = conv_mac_85 + 15'd8488;
logic [31:0] bias_add_86;
assign bias_add_86 = conv_mac_86 + 15'd14953;
logic [31:0] bias_add_87;
assign bias_add_87 = conv_mac_87 + 15'd12642;
logic [31:0] bias_add_88;
assign bias_add_88 = conv_mac_88 + 15'd9972;
logic [31:0] bias_add_89;
assign bias_add_89 = conv_mac_89 + 15'd9010;
logic [31:0] bias_add_90;
assign bias_add_90 = conv_mac_90 + 15'd9616;
logic [31:0] bias_add_91;
assign bias_add_91 = conv_mac_91 + 14'd4549;
logic [31:0] bias_add_92;
assign bias_add_92 = conv_mac_92 + 15'd10409;
logic [31:0] bias_add_93;
assign bias_add_93 = conv_mac_93 + 16'd31986;
logic [31:0] bias_add_94;
assign bias_add_94 = conv_mac_94 + 16'd18830;
logic [31:0] bias_add_95;
assign bias_add_95 = conv_mac_95 + 16'd18613;
logic [31:0] bias_add_96;
assign bias_add_96 = conv_mac_96 + 16'd19058;
logic [31:0] bias_add_97;
assign bias_add_97 = conv_mac_97 + 14'd6978;
logic [31:0] bias_add_98;
assign bias_add_98 = conv_mac_98 + 16'd21915;
logic [31:0] bias_add_99;
assign bias_add_99 = conv_mac_99 + 16'd23132;
logic [31:0] bias_add_100;
assign bias_add_100 = conv_mac_100 + 16'd18384;
logic [31:0] bias_add_101;
assign bias_add_101 = conv_mac_101 + 15'd13636;
logic [31:0] bias_add_102;
assign bias_add_102 = conv_mac_102 + 12'd1373;
logic [31:0] bias_add_103;
assign bias_add_103 = conv_mac_103 + 15'd13904;
logic [31:0] bias_add_104;
assign bias_add_104 = conv_mac_104 + 16'd18861;
logic [31:0] bias_add_105;
assign bias_add_105 = conv_mac_105 + 16'd28669;
logic [31:0] bias_add_106;
assign bias_add_106 = conv_mac_106 + 15'd16363;
logic [31:0] bias_add_107;
assign bias_add_107 = conv_mac_107 + 16'd26130;
logic [31:0] bias_add_108;
assign bias_add_108 = conv_mac_108 + 14'd5604;
logic [31:0] bias_add_109;
assign bias_add_109 = conv_mac_109 + 16'd29476;
logic [31:0] bias_add_110;
assign bias_add_110 = conv_mac_110 + 16'd17671;
logic [31:0] bias_add_111;
assign bias_add_111 = conv_mac_111 + 15'd9918;
logic [31:0] bias_add_112;
assign bias_add_112 = conv_mac_112 + 16'd17555;
logic [31:0] bias_add_113;
assign bias_add_113 = conv_mac_113 + 11'd870;
logic [31:0] bias_add_114;
assign bias_add_114 = conv_mac_114 + 15'd14412;
logic [31:0] bias_add_115;
assign bias_add_115 = conv_mac_115 + 16'd31179;
logic [31:0] bias_add_116;
assign bias_add_116 = conv_mac_116 + 13'd4062;
logic [31:0] bias_add_117;
assign bias_add_117 = conv_mac_117 + 13'd3679;
logic [31:0] bias_add_118;
assign bias_add_118 = conv_mac_118 + 16'd26464;
logic [31:0] bias_add_119;
assign bias_add_119 = conv_mac_119 + 16'd19404;
logic [31:0] bias_add_120;
assign bias_add_120 = conv_mac_120 + 16'd19459;
logic [31:0] bias_add_121;
assign bias_add_121 = conv_mac_121 + 16'd19093;
logic [31:0] bias_add_122;
assign bias_add_122 = conv_mac_122 + 16'd17391;
logic [31:0] bias_add_123;
assign bias_add_123 = conv_mac_123 + 16'd20253;
logic [31:0] bias_add_124;
assign bias_add_124 = conv_mac_124 + 14'd7705;
logic [31:0] bias_add_125;
assign bias_add_125 = conv_mac_125 + 16'd30661;
logic [31:0] bias_add_126;
assign bias_add_126 = conv_mac_126 + 16'd22795;
logic [31:0] bias_add_127;
assign bias_add_127 = conv_mac_127 + 16'd19114;
logic [31:0] bias_add_128;
assign bias_add_128 = conv_mac_128 + 15'd11097;
logic [31:0] bias_add_129;
assign bias_add_129 = conv_mac_129 + 15'd9037;
logic [31:0] bias_add_130;
assign bias_add_130 = conv_mac_130 + 14'd5001;
logic [31:0] bias_add_131;
assign bias_add_131 = conv_mac_131 + 15'd12623;
logic [31:0] bias_add_132;
assign bias_add_132 = conv_mac_132 + 16'd27310;
logic [31:0] bias_add_133;
assign bias_add_133 = conv_mac_133 + 16'd18246;
logic [31:0] bias_add_134;
assign bias_add_134 = conv_mac_134 + 16'd16615;
logic [31:0] bias_add_135;
assign bias_add_135 = conv_mac_135 + 16'd30107;
logic [31:0] bias_add_136;
assign bias_add_136 = conv_mac_136 + 16'd27158;
logic [31:0] bias_add_137;
assign bias_add_137 = conv_mac_137 + 16'd31955;
logic [31:0] bias_add_138;
assign bias_add_138 = conv_mac_138 + 16'd21800;
logic [31:0] bias_add_139;
assign bias_add_139 = conv_mac_139 + 10'd384;
logic [31:0] bias_add_140;
assign bias_add_140 = conv_mac_140 + 15'd8821;
logic [31:0] bias_add_141;
assign bias_add_141 = conv_mac_141 + 14'd6768;
logic [31:0] bias_add_142;
assign bias_add_142 = conv_mac_142 + 9'd179;
logic [31:0] bias_add_143;
assign bias_add_143 = conv_mac_143 + 16'd32362;
logic [31:0] bias_add_144;
assign bias_add_144 = conv_mac_144 + 16'd17393;
logic [31:0] bias_add_145;
assign bias_add_145 = conv_mac_145 + 15'd12336;
logic [31:0] bias_add_146;
assign bias_add_146 = conv_mac_146 + 14'd4971;
logic [31:0] bias_add_147;
assign bias_add_147 = conv_mac_147 + 16'd28531;
logic [31:0] bias_add_148;
assign bias_add_148 = conv_mac_148 + 16'd19618;
logic [31:0] bias_add_149;
assign bias_add_149 = conv_mac_149 + 16'd27649;
logic [31:0] bias_add_150;
assign bias_add_150 = conv_mac_150 + 13'd3695;
logic [31:0] bias_add_151;
assign bias_add_151 = conv_mac_151 + 16'd17256;
logic [31:0] bias_add_152;
assign bias_add_152 = conv_mac_152 + 15'd16237;
logic [31:0] bias_add_153;
assign bias_add_153 = conv_mac_153 + 16'd29298;
logic [31:0] bias_add_154;
assign bias_add_154 = conv_mac_154 + 15'd12133;
logic [31:0] bias_add_155;
assign bias_add_155 = conv_mac_155 + 15'd9467;
logic [31:0] bias_add_156;
assign bias_add_156 = conv_mac_156 + 16'd31874;
logic [31:0] bias_add_157;
assign bias_add_157 = conv_mac_157 + 10'd482;
logic [31:0] bias_add_158;
assign bias_add_158 = conv_mac_158 + 15'd11942;
logic [31:0] bias_add_159;
assign bias_add_159 = conv_mac_159 + 16'd20749;
logic [31:0] bias_add_160;
assign bias_add_160 = conv_mac_160 + 16'd26541;
logic [31:0] bias_add_161;
assign bias_add_161 = conv_mac_161 + 16'd16870;
logic [31:0] bias_add_162;
assign bias_add_162 = conv_mac_162 + 16'd17767;
logic [31:0] bias_add_163;
assign bias_add_163 = conv_mac_163 + 16'd30739;
logic [31:0] bias_add_164;
assign bias_add_164 = conv_mac_164 + 16'd26038;
logic [31:0] bias_add_165;
assign bias_add_165 = conv_mac_165 + 16'd27217;
logic [31:0] bias_add_166;
assign bias_add_166 = conv_mac_166 + 13'd2698;
logic [31:0] bias_add_167;
assign bias_add_167 = conv_mac_167 + 16'd22569;
logic [31:0] bias_add_168;
assign bias_add_168 = conv_mac_168 + 16'd17976;
logic [31:0] bias_add_169;
assign bias_add_169 = conv_mac_169 + 16'd24612;
logic [31:0] bias_add_170;
assign bias_add_170 = conv_mac_170 + 16'd23987;
logic [31:0] bias_add_171;
assign bias_add_171 = conv_mac_171 + 16'd19199;
logic [31:0] bias_add_172;
assign bias_add_172 = conv_mac_172 + 16'd29596;
logic [31:0] bias_add_173;
assign bias_add_173 = conv_mac_173 + 16'd25265;
logic [31:0] bias_add_174;
assign bias_add_174 = conv_mac_174 + 12'd1337;
logic [31:0] bias_add_175;
assign bias_add_175 = conv_mac_175 + 16'd26882;
logic [31:0] bias_add_176;
assign bias_add_176 = conv_mac_176 + 16'd23448;
logic [31:0] bias_add_177;
assign bias_add_177 = conv_mac_177 + 13'd3937;
logic [31:0] bias_add_178;
assign bias_add_178 = conv_mac_178 + 16'd23933;
logic [31:0] bias_add_179;
assign bias_add_179 = conv_mac_179 + 16'd24352;
logic [31:0] bias_add_180;
assign bias_add_180 = conv_mac_180 + 16'd22556;
logic [31:0] bias_add_181;
assign bias_add_181 = conv_mac_181 + 16'd21436;
logic [31:0] bias_add_182;
assign bias_add_182 = conv_mac_182 + 16'd17577;
logic [31:0] bias_add_183;
assign bias_add_183 = conv_mac_183 + 16'd32456;
logic [31:0] bias_add_184;
assign bias_add_184 = conv_mac_184 + 15'd14956;
logic [31:0] bias_add_185;
assign bias_add_185 = conv_mac_185 + 15'd14634;
logic [31:0] bias_add_186;
assign bias_add_186 = conv_mac_186 + 15'd10826;
logic [31:0] bias_add_187;
assign bias_add_187 = conv_mac_187 + 15'd14925;
logic [31:0] bias_add_188;
assign bias_add_188 = conv_mac_188 + 16'd27059;
logic [31:0] bias_add_189;
assign bias_add_189 = conv_mac_189 + 14'd7046;
logic [31:0] bias_add_190;
assign bias_add_190 = conv_mac_190 + 9'd248;
logic [31:0] bias_add_191;
assign bias_add_191 = conv_mac_191 + 12'd1810;
logic [31:0] bias_add_192;
assign bias_add_192 = conv_mac_192 + 16'd21379;
logic [31:0] bias_add_193;
assign bias_add_193 = conv_mac_193 + 16'd20301;
logic [31:0] bias_add_194;
assign bias_add_194 = conv_mac_194 + 16'd19852;
logic [31:0] bias_add_195;
assign bias_add_195 = conv_mac_195 + 14'd5090;
logic [31:0] bias_add_196;
assign bias_add_196 = conv_mac_196 + 14'd4816;
logic [31:0] bias_add_197;
assign bias_add_197 = conv_mac_197 + 16'd30945;
logic [31:0] bias_add_198;
assign bias_add_198 = conv_mac_198 + 16'd17298;
logic [31:0] bias_add_199;
assign bias_add_199 = conv_mac_199 + 14'd6839;
logic [31:0] bias_add_200;
assign bias_add_200 = conv_mac_200 + 13'd2198;
logic [31:0] bias_add_201;
assign bias_add_201 = conv_mac_201 + 14'd5477;
logic [31:0] bias_add_202;
assign bias_add_202 = conv_mac_202 + 16'd26485;
logic [31:0] bias_add_203;
assign bias_add_203 = conv_mac_203 + 13'd2200;
logic [31:0] bias_add_204;
assign bias_add_204 = conv_mac_204 + 16'd26974;
logic [31:0] bias_add_205;
assign bias_add_205 = conv_mac_205 + 16'd23427;
logic [31:0] bias_add_206;
assign bias_add_206 = conv_mac_206 + 15'd12721;
logic [31:0] bias_add_207;
assign bias_add_207 = conv_mac_207 + 15'd13007;
logic [31:0] bias_add_208;
assign bias_add_208 = conv_mac_208 + 16'd26948;
logic [31:0] bias_add_209;
assign bias_add_209 = conv_mac_209 + 16'd21295;
logic [31:0] bias_add_210;
assign bias_add_210 = conv_mac_210 + 16'd24066;
logic [31:0] bias_add_211;
assign bias_add_211 = conv_mac_211 + 16'd24630;
logic [31:0] bias_add_212;
assign bias_add_212 = conv_mac_212 + 11'd636;
logic [31:0] bias_add_213;
assign bias_add_213 = conv_mac_213 + 16'd19922;
logic [31:0] bias_add_214;
assign bias_add_214 = conv_mac_214 + 16'd23880;
logic [31:0] bias_add_215;
assign bias_add_215 = conv_mac_215 + 16'd22037;
logic [31:0] bias_add_216;
assign bias_add_216 = conv_mac_216 + 16'd25294;
logic [31:0] bias_add_217;
assign bias_add_217 = conv_mac_217 + 13'd2602;
logic [31:0] bias_add_218;
assign bias_add_218 = conv_mac_218 + 16'd32711;
logic [31:0] bias_add_219;
assign bias_add_219 = conv_mac_219 + 13'd3700;
logic [31:0] bias_add_220;
assign bias_add_220 = conv_mac_220 + 14'd4731;
logic [31:0] bias_add_221;
assign bias_add_221 = conv_mac_221 + 14'd7313;
logic [31:0] bias_add_222;
assign bias_add_222 = conv_mac_222 + 16'd16456;
logic [31:0] bias_add_223;
assign bias_add_223 = conv_mac_223 + 14'd4950;
logic [31:0] bias_add_224;
assign bias_add_224 = conv_mac_224 + 16'd28724;
logic [31:0] bias_add_225;
assign bias_add_225 = conv_mac_225 + 16'd25548;
logic [31:0] bias_add_226;
assign bias_add_226 = conv_mac_226 + 15'd14135;
logic [31:0] bias_add_227;
assign bias_add_227 = conv_mac_227 + 13'd3666;
logic [31:0] bias_add_228;
assign bias_add_228 = conv_mac_228 + 15'd12235;
logic [31:0] bias_add_229;
assign bias_add_229 = conv_mac_229 + 13'd2185;
logic [31:0] bias_add_230;
assign bias_add_230 = conv_mac_230 + 15'd11702;
logic [31:0] bias_add_231;
assign bias_add_231 = conv_mac_231 + 16'd29372;
logic [31:0] bias_add_232;
assign bias_add_232 = conv_mac_232 + 15'd11569;
logic [31:0] bias_add_233;
assign bias_add_233 = conv_mac_233 + 16'd24953;
logic [31:0] bias_add_234;
assign bias_add_234 = conv_mac_234 + 14'd5935;
logic [31:0] bias_add_235;
assign bias_add_235 = conv_mac_235 + 16'd26787;
logic [31:0] bias_add_236;
assign bias_add_236 = conv_mac_236 + 12'd1174;
logic [31:0] bias_add_237;
assign bias_add_237 = conv_mac_237 + 16'd30800;
logic [31:0] bias_add_238;
assign bias_add_238 = conv_mac_238 + 14'd5956;
logic [31:0] bias_add_239;
assign bias_add_239 = conv_mac_239 + 15'd14848;
logic [31:0] bias_add_240;
assign bias_add_240 = conv_mac_240 + 16'd25162;
logic [31:0] bias_add_241;
assign bias_add_241 = conv_mac_241 + 13'd3054;
logic [31:0] bias_add_242;
assign bias_add_242 = conv_mac_242 + 15'd12989;
logic [31:0] bias_add_243;
assign bias_add_243 = conv_mac_243 + 14'd5057;
logic [31:0] bias_add_244;
assign bias_add_244 = conv_mac_244 + 16'd30973;
logic [31:0] bias_add_245;
assign bias_add_245 = conv_mac_245 + 16'd26726;
logic [31:0] bias_add_246;
assign bias_add_246 = conv_mac_246 + 16'd16980;
logic [31:0] bias_add_247;
assign bias_add_247 = conv_mac_247 + 16'd31724;
logic [31:0] bias_add_248;
assign bias_add_248 = conv_mac_248 + 16'd18228;
logic [31:0] bias_add_249;
assign bias_add_249 = conv_mac_249 + 16'd28461;
logic [31:0] bias_add_250;
assign bias_add_250 = conv_mac_250 + 13'd3476;
logic [31:0] bias_add_251;
assign bias_add_251 = conv_mac_251 + 16'd26105;
logic [31:0] bias_add_252;
assign bias_add_252 = conv_mac_252 + 16'd25605;
logic [31:0] bias_add_253;
assign bias_add_253 = conv_mac_253 + 12'd1819;
logic [31:0] bias_add_254;
assign bias_add_254 = conv_mac_254 + 15'd11908;
logic [31:0] bias_add_255;
assign bias_add_255 = conv_mac_255 + 14'd5487;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[21:15]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[21:15]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[21:15]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[21:15]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[21:15]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[21:15]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[21:15]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[21:15]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[21:15]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[21:15]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[21:15]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[21:15]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[21:15]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[21:15]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[21:15]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[21:15]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[21:15]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[21:15]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[21:15]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[21:15]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[21:15]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[21:15]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[21:15]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[21:15]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[21:15]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[21:15]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[21:15]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[21:15]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[21:15]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[21:15]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[21:15]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[21:15]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[21:15]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[21:15]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[21:15]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[21:15]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[21:15]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[21:15]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[21:15]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[21:15]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[21:15]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[21:15]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[21:15]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[21:15]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[21:15]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[21:15]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[21:15]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[21:15]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[21:15]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[21:15]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[21:15]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[21:15]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[21:15]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[21:15]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[21:15]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[21:15]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[21:15]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[21:15]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[21:15]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[21:15]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[21:15]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[21:15]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[21:15]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[21:15]}} :'d6) : '0;
logic [7:0] relu_64;
assign relu_64[7:0] = (bias_add_64[31]==0) ? ((bias_add_64<3'd6) ? {{bias_add_64[31],bias_add_64[21:15]}} :'d6) : '0;
logic [7:0] relu_65;
assign relu_65[7:0] = (bias_add_65[31]==0) ? ((bias_add_65<3'd6) ? {{bias_add_65[31],bias_add_65[21:15]}} :'d6) : '0;
logic [7:0] relu_66;
assign relu_66[7:0] = (bias_add_66[31]==0) ? ((bias_add_66<3'd6) ? {{bias_add_66[31],bias_add_66[21:15]}} :'d6) : '0;
logic [7:0] relu_67;
assign relu_67[7:0] = (bias_add_67[31]==0) ? ((bias_add_67<3'd6) ? {{bias_add_67[31],bias_add_67[21:15]}} :'d6) : '0;
logic [7:0] relu_68;
assign relu_68[7:0] = (bias_add_68[31]==0) ? ((bias_add_68<3'd6) ? {{bias_add_68[31],bias_add_68[21:15]}} :'d6) : '0;
logic [7:0] relu_69;
assign relu_69[7:0] = (bias_add_69[31]==0) ? ((bias_add_69<3'd6) ? {{bias_add_69[31],bias_add_69[21:15]}} :'d6) : '0;
logic [7:0] relu_70;
assign relu_70[7:0] = (bias_add_70[31]==0) ? ((bias_add_70<3'd6) ? {{bias_add_70[31],bias_add_70[21:15]}} :'d6) : '0;
logic [7:0] relu_71;
assign relu_71[7:0] = (bias_add_71[31]==0) ? ((bias_add_71<3'd6) ? {{bias_add_71[31],bias_add_71[21:15]}} :'d6) : '0;
logic [7:0] relu_72;
assign relu_72[7:0] = (bias_add_72[31]==0) ? ((bias_add_72<3'd6) ? {{bias_add_72[31],bias_add_72[21:15]}} :'d6) : '0;
logic [7:0] relu_73;
assign relu_73[7:0] = (bias_add_73[31]==0) ? ((bias_add_73<3'd6) ? {{bias_add_73[31],bias_add_73[21:15]}} :'d6) : '0;
logic [7:0] relu_74;
assign relu_74[7:0] = (bias_add_74[31]==0) ? ((bias_add_74<3'd6) ? {{bias_add_74[31],bias_add_74[21:15]}} :'d6) : '0;
logic [7:0] relu_75;
assign relu_75[7:0] = (bias_add_75[31]==0) ? ((bias_add_75<3'd6) ? {{bias_add_75[31],bias_add_75[21:15]}} :'d6) : '0;
logic [7:0] relu_76;
assign relu_76[7:0] = (bias_add_76[31]==0) ? ((bias_add_76<3'd6) ? {{bias_add_76[31],bias_add_76[21:15]}} :'d6) : '0;
logic [7:0] relu_77;
assign relu_77[7:0] = (bias_add_77[31]==0) ? ((bias_add_77<3'd6) ? {{bias_add_77[31],bias_add_77[21:15]}} :'d6) : '0;
logic [7:0] relu_78;
assign relu_78[7:0] = (bias_add_78[31]==0) ? ((bias_add_78<3'd6) ? {{bias_add_78[31],bias_add_78[21:15]}} :'d6) : '0;
logic [7:0] relu_79;
assign relu_79[7:0] = (bias_add_79[31]==0) ? ((bias_add_79<3'd6) ? {{bias_add_79[31],bias_add_79[21:15]}} :'d6) : '0;
logic [7:0] relu_80;
assign relu_80[7:0] = (bias_add_80[31]==0) ? ((bias_add_80<3'd6) ? {{bias_add_80[31],bias_add_80[21:15]}} :'d6) : '0;
logic [7:0] relu_81;
assign relu_81[7:0] = (bias_add_81[31]==0) ? ((bias_add_81<3'd6) ? {{bias_add_81[31],bias_add_81[21:15]}} :'d6) : '0;
logic [7:0] relu_82;
assign relu_82[7:0] = (bias_add_82[31]==0) ? ((bias_add_82<3'd6) ? {{bias_add_82[31],bias_add_82[21:15]}} :'d6) : '0;
logic [7:0] relu_83;
assign relu_83[7:0] = (bias_add_83[31]==0) ? ((bias_add_83<3'd6) ? {{bias_add_83[31],bias_add_83[21:15]}} :'d6) : '0;
logic [7:0] relu_84;
assign relu_84[7:0] = (bias_add_84[31]==0) ? ((bias_add_84<3'd6) ? {{bias_add_84[31],bias_add_84[21:15]}} :'d6) : '0;
logic [7:0] relu_85;
assign relu_85[7:0] = (bias_add_85[31]==0) ? ((bias_add_85<3'd6) ? {{bias_add_85[31],bias_add_85[21:15]}} :'d6) : '0;
logic [7:0] relu_86;
assign relu_86[7:0] = (bias_add_86[31]==0) ? ((bias_add_86<3'd6) ? {{bias_add_86[31],bias_add_86[21:15]}} :'d6) : '0;
logic [7:0] relu_87;
assign relu_87[7:0] = (bias_add_87[31]==0) ? ((bias_add_87<3'd6) ? {{bias_add_87[31],bias_add_87[21:15]}} :'d6) : '0;
logic [7:0] relu_88;
assign relu_88[7:0] = (bias_add_88[31]==0) ? ((bias_add_88<3'd6) ? {{bias_add_88[31],bias_add_88[21:15]}} :'d6) : '0;
logic [7:0] relu_89;
assign relu_89[7:0] = (bias_add_89[31]==0) ? ((bias_add_89<3'd6) ? {{bias_add_89[31],bias_add_89[21:15]}} :'d6) : '0;
logic [7:0] relu_90;
assign relu_90[7:0] = (bias_add_90[31]==0) ? ((bias_add_90<3'd6) ? {{bias_add_90[31],bias_add_90[21:15]}} :'d6) : '0;
logic [7:0] relu_91;
assign relu_91[7:0] = (bias_add_91[31]==0) ? ((bias_add_91<3'd6) ? {{bias_add_91[31],bias_add_91[21:15]}} :'d6) : '0;
logic [7:0] relu_92;
assign relu_92[7:0] = (bias_add_92[31]==0) ? ((bias_add_92<3'd6) ? {{bias_add_92[31],bias_add_92[21:15]}} :'d6) : '0;
logic [7:0] relu_93;
assign relu_93[7:0] = (bias_add_93[31]==0) ? ((bias_add_93<3'd6) ? {{bias_add_93[31],bias_add_93[21:15]}} :'d6) : '0;
logic [7:0] relu_94;
assign relu_94[7:0] = (bias_add_94[31]==0) ? ((bias_add_94<3'd6) ? {{bias_add_94[31],bias_add_94[21:15]}} :'d6) : '0;
logic [7:0] relu_95;
assign relu_95[7:0] = (bias_add_95[31]==0) ? ((bias_add_95<3'd6) ? {{bias_add_95[31],bias_add_95[21:15]}} :'d6) : '0;
logic [7:0] relu_96;
assign relu_96[7:0] = (bias_add_96[31]==0) ? ((bias_add_96<3'd6) ? {{bias_add_96[31],bias_add_96[21:15]}} :'d6) : '0;
logic [7:0] relu_97;
assign relu_97[7:0] = (bias_add_97[31]==0) ? ((bias_add_97<3'd6) ? {{bias_add_97[31],bias_add_97[21:15]}} :'d6) : '0;
logic [7:0] relu_98;
assign relu_98[7:0] = (bias_add_98[31]==0) ? ((bias_add_98<3'd6) ? {{bias_add_98[31],bias_add_98[21:15]}} :'d6) : '0;
logic [7:0] relu_99;
assign relu_99[7:0] = (bias_add_99[31]==0) ? ((bias_add_99<3'd6) ? {{bias_add_99[31],bias_add_99[21:15]}} :'d6) : '0;
logic [7:0] relu_100;
assign relu_100[7:0] = (bias_add_100[31]==0) ? ((bias_add_100<3'd6) ? {{bias_add_100[31],bias_add_100[21:15]}} :'d6) : '0;
logic [7:0] relu_101;
assign relu_101[7:0] = (bias_add_101[31]==0) ? ((bias_add_101<3'd6) ? {{bias_add_101[31],bias_add_101[21:15]}} :'d6) : '0;
logic [7:0] relu_102;
assign relu_102[7:0] = (bias_add_102[31]==0) ? ((bias_add_102<3'd6) ? {{bias_add_102[31],bias_add_102[21:15]}} :'d6) : '0;
logic [7:0] relu_103;
assign relu_103[7:0] = (bias_add_103[31]==0) ? ((bias_add_103<3'd6) ? {{bias_add_103[31],bias_add_103[21:15]}} :'d6) : '0;
logic [7:0] relu_104;
assign relu_104[7:0] = (bias_add_104[31]==0) ? ((bias_add_104<3'd6) ? {{bias_add_104[31],bias_add_104[21:15]}} :'d6) : '0;
logic [7:0] relu_105;
assign relu_105[7:0] = (bias_add_105[31]==0) ? ((bias_add_105<3'd6) ? {{bias_add_105[31],bias_add_105[21:15]}} :'d6) : '0;
logic [7:0] relu_106;
assign relu_106[7:0] = (bias_add_106[31]==0) ? ((bias_add_106<3'd6) ? {{bias_add_106[31],bias_add_106[21:15]}} :'d6) : '0;
logic [7:0] relu_107;
assign relu_107[7:0] = (bias_add_107[31]==0) ? ((bias_add_107<3'd6) ? {{bias_add_107[31],bias_add_107[21:15]}} :'d6) : '0;
logic [7:0] relu_108;
assign relu_108[7:0] = (bias_add_108[31]==0) ? ((bias_add_108<3'd6) ? {{bias_add_108[31],bias_add_108[21:15]}} :'d6) : '0;
logic [7:0] relu_109;
assign relu_109[7:0] = (bias_add_109[31]==0) ? ((bias_add_109<3'd6) ? {{bias_add_109[31],bias_add_109[21:15]}} :'d6) : '0;
logic [7:0] relu_110;
assign relu_110[7:0] = (bias_add_110[31]==0) ? ((bias_add_110<3'd6) ? {{bias_add_110[31],bias_add_110[21:15]}} :'d6) : '0;
logic [7:0] relu_111;
assign relu_111[7:0] = (bias_add_111[31]==0) ? ((bias_add_111<3'd6) ? {{bias_add_111[31],bias_add_111[21:15]}} :'d6) : '0;
logic [7:0] relu_112;
assign relu_112[7:0] = (bias_add_112[31]==0) ? ((bias_add_112<3'd6) ? {{bias_add_112[31],bias_add_112[21:15]}} :'d6) : '0;
logic [7:0] relu_113;
assign relu_113[7:0] = (bias_add_113[31]==0) ? ((bias_add_113<3'd6) ? {{bias_add_113[31],bias_add_113[21:15]}} :'d6) : '0;
logic [7:0] relu_114;
assign relu_114[7:0] = (bias_add_114[31]==0) ? ((bias_add_114<3'd6) ? {{bias_add_114[31],bias_add_114[21:15]}} :'d6) : '0;
logic [7:0] relu_115;
assign relu_115[7:0] = (bias_add_115[31]==0) ? ((bias_add_115<3'd6) ? {{bias_add_115[31],bias_add_115[21:15]}} :'d6) : '0;
logic [7:0] relu_116;
assign relu_116[7:0] = (bias_add_116[31]==0) ? ((bias_add_116<3'd6) ? {{bias_add_116[31],bias_add_116[21:15]}} :'d6) : '0;
logic [7:0] relu_117;
assign relu_117[7:0] = (bias_add_117[31]==0) ? ((bias_add_117<3'd6) ? {{bias_add_117[31],bias_add_117[21:15]}} :'d6) : '0;
logic [7:0] relu_118;
assign relu_118[7:0] = (bias_add_118[31]==0) ? ((bias_add_118<3'd6) ? {{bias_add_118[31],bias_add_118[21:15]}} :'d6) : '0;
logic [7:0] relu_119;
assign relu_119[7:0] = (bias_add_119[31]==0) ? ((bias_add_119<3'd6) ? {{bias_add_119[31],bias_add_119[21:15]}} :'d6) : '0;
logic [7:0] relu_120;
assign relu_120[7:0] = (bias_add_120[31]==0) ? ((bias_add_120<3'd6) ? {{bias_add_120[31],bias_add_120[21:15]}} :'d6) : '0;
logic [7:0] relu_121;
assign relu_121[7:0] = (bias_add_121[31]==0) ? ((bias_add_121<3'd6) ? {{bias_add_121[31],bias_add_121[21:15]}} :'d6) : '0;
logic [7:0] relu_122;
assign relu_122[7:0] = (bias_add_122[31]==0) ? ((bias_add_122<3'd6) ? {{bias_add_122[31],bias_add_122[21:15]}} :'d6) : '0;
logic [7:0] relu_123;
assign relu_123[7:0] = (bias_add_123[31]==0) ? ((bias_add_123<3'd6) ? {{bias_add_123[31],bias_add_123[21:15]}} :'d6) : '0;
logic [7:0] relu_124;
assign relu_124[7:0] = (bias_add_124[31]==0) ? ((bias_add_124<3'd6) ? {{bias_add_124[31],bias_add_124[21:15]}} :'d6) : '0;
logic [7:0] relu_125;
assign relu_125[7:0] = (bias_add_125[31]==0) ? ((bias_add_125<3'd6) ? {{bias_add_125[31],bias_add_125[21:15]}} :'d6) : '0;
logic [7:0] relu_126;
assign relu_126[7:0] = (bias_add_126[31]==0) ? ((bias_add_126<3'd6) ? {{bias_add_126[31],bias_add_126[21:15]}} :'d6) : '0;
logic [7:0] relu_127;
assign relu_127[7:0] = (bias_add_127[31]==0) ? ((bias_add_127<3'd6) ? {{bias_add_127[31],bias_add_127[21:15]}} :'d6) : '0;
logic [7:0] relu_128;
assign relu_128[7:0] = (bias_add_128[31]==0) ? ((bias_add_128<3'd6) ? {{bias_add_128[31],bias_add_128[21:15]}} :'d6) : '0;
logic [7:0] relu_129;
assign relu_129[7:0] = (bias_add_129[31]==0) ? ((bias_add_129<3'd6) ? {{bias_add_129[31],bias_add_129[21:15]}} :'d6) : '0;
logic [7:0] relu_130;
assign relu_130[7:0] = (bias_add_130[31]==0) ? ((bias_add_130<3'd6) ? {{bias_add_130[31],bias_add_130[21:15]}} :'d6) : '0;
logic [7:0] relu_131;
assign relu_131[7:0] = (bias_add_131[31]==0) ? ((bias_add_131<3'd6) ? {{bias_add_131[31],bias_add_131[21:15]}} :'d6) : '0;
logic [7:0] relu_132;
assign relu_132[7:0] = (bias_add_132[31]==0) ? ((bias_add_132<3'd6) ? {{bias_add_132[31],bias_add_132[21:15]}} :'d6) : '0;
logic [7:0] relu_133;
assign relu_133[7:0] = (bias_add_133[31]==0) ? ((bias_add_133<3'd6) ? {{bias_add_133[31],bias_add_133[21:15]}} :'d6) : '0;
logic [7:0] relu_134;
assign relu_134[7:0] = (bias_add_134[31]==0) ? ((bias_add_134<3'd6) ? {{bias_add_134[31],bias_add_134[21:15]}} :'d6) : '0;
logic [7:0] relu_135;
assign relu_135[7:0] = (bias_add_135[31]==0) ? ((bias_add_135<3'd6) ? {{bias_add_135[31],bias_add_135[21:15]}} :'d6) : '0;
logic [7:0] relu_136;
assign relu_136[7:0] = (bias_add_136[31]==0) ? ((bias_add_136<3'd6) ? {{bias_add_136[31],bias_add_136[21:15]}} :'d6) : '0;
logic [7:0] relu_137;
assign relu_137[7:0] = (bias_add_137[31]==0) ? ((bias_add_137<3'd6) ? {{bias_add_137[31],bias_add_137[21:15]}} :'d6) : '0;
logic [7:0] relu_138;
assign relu_138[7:0] = (bias_add_138[31]==0) ? ((bias_add_138<3'd6) ? {{bias_add_138[31],bias_add_138[21:15]}} :'d6) : '0;
logic [7:0] relu_139;
assign relu_139[7:0] = (bias_add_139[31]==0) ? ((bias_add_139<3'd6) ? {{bias_add_139[31],bias_add_139[21:15]}} :'d6) : '0;
logic [7:0] relu_140;
assign relu_140[7:0] = (bias_add_140[31]==0) ? ((bias_add_140<3'd6) ? {{bias_add_140[31],bias_add_140[21:15]}} :'d6) : '0;
logic [7:0] relu_141;
assign relu_141[7:0] = (bias_add_141[31]==0) ? ((bias_add_141<3'd6) ? {{bias_add_141[31],bias_add_141[21:15]}} :'d6) : '0;
logic [7:0] relu_142;
assign relu_142[7:0] = (bias_add_142[31]==0) ? ((bias_add_142<3'd6) ? {{bias_add_142[31],bias_add_142[21:15]}} :'d6) : '0;
logic [7:0] relu_143;
assign relu_143[7:0] = (bias_add_143[31]==0) ? ((bias_add_143<3'd6) ? {{bias_add_143[31],bias_add_143[21:15]}} :'d6) : '0;
logic [7:0] relu_144;
assign relu_144[7:0] = (bias_add_144[31]==0) ? ((bias_add_144<3'd6) ? {{bias_add_144[31],bias_add_144[21:15]}} :'d6) : '0;
logic [7:0] relu_145;
assign relu_145[7:0] = (bias_add_145[31]==0) ? ((bias_add_145<3'd6) ? {{bias_add_145[31],bias_add_145[21:15]}} :'d6) : '0;
logic [7:0] relu_146;
assign relu_146[7:0] = (bias_add_146[31]==0) ? ((bias_add_146<3'd6) ? {{bias_add_146[31],bias_add_146[21:15]}} :'d6) : '0;
logic [7:0] relu_147;
assign relu_147[7:0] = (bias_add_147[31]==0) ? ((bias_add_147<3'd6) ? {{bias_add_147[31],bias_add_147[21:15]}} :'d6) : '0;
logic [7:0] relu_148;
assign relu_148[7:0] = (bias_add_148[31]==0) ? ((bias_add_148<3'd6) ? {{bias_add_148[31],bias_add_148[21:15]}} :'d6) : '0;
logic [7:0] relu_149;
assign relu_149[7:0] = (bias_add_149[31]==0) ? ((bias_add_149<3'd6) ? {{bias_add_149[31],bias_add_149[21:15]}} :'d6) : '0;
logic [7:0] relu_150;
assign relu_150[7:0] = (bias_add_150[31]==0) ? ((bias_add_150<3'd6) ? {{bias_add_150[31],bias_add_150[21:15]}} :'d6) : '0;
logic [7:0] relu_151;
assign relu_151[7:0] = (bias_add_151[31]==0) ? ((bias_add_151<3'd6) ? {{bias_add_151[31],bias_add_151[21:15]}} :'d6) : '0;
logic [7:0] relu_152;
assign relu_152[7:0] = (bias_add_152[31]==0) ? ((bias_add_152<3'd6) ? {{bias_add_152[31],bias_add_152[21:15]}} :'d6) : '0;
logic [7:0] relu_153;
assign relu_153[7:0] = (bias_add_153[31]==0) ? ((bias_add_153<3'd6) ? {{bias_add_153[31],bias_add_153[21:15]}} :'d6) : '0;
logic [7:0] relu_154;
assign relu_154[7:0] = (bias_add_154[31]==0) ? ((bias_add_154<3'd6) ? {{bias_add_154[31],bias_add_154[21:15]}} :'d6) : '0;
logic [7:0] relu_155;
assign relu_155[7:0] = (bias_add_155[31]==0) ? ((bias_add_155<3'd6) ? {{bias_add_155[31],bias_add_155[21:15]}} :'d6) : '0;
logic [7:0] relu_156;
assign relu_156[7:0] = (bias_add_156[31]==0) ? ((bias_add_156<3'd6) ? {{bias_add_156[31],bias_add_156[21:15]}} :'d6) : '0;
logic [7:0] relu_157;
assign relu_157[7:0] = (bias_add_157[31]==0) ? ((bias_add_157<3'd6) ? {{bias_add_157[31],bias_add_157[21:15]}} :'d6) : '0;
logic [7:0] relu_158;
assign relu_158[7:0] = (bias_add_158[31]==0) ? ((bias_add_158<3'd6) ? {{bias_add_158[31],bias_add_158[21:15]}} :'d6) : '0;
logic [7:0] relu_159;
assign relu_159[7:0] = (bias_add_159[31]==0) ? ((bias_add_159<3'd6) ? {{bias_add_159[31],bias_add_159[21:15]}} :'d6) : '0;
logic [7:0] relu_160;
assign relu_160[7:0] = (bias_add_160[31]==0) ? ((bias_add_160<3'd6) ? {{bias_add_160[31],bias_add_160[21:15]}} :'d6) : '0;
logic [7:0] relu_161;
assign relu_161[7:0] = (bias_add_161[31]==0) ? ((bias_add_161<3'd6) ? {{bias_add_161[31],bias_add_161[21:15]}} :'d6) : '0;
logic [7:0] relu_162;
assign relu_162[7:0] = (bias_add_162[31]==0) ? ((bias_add_162<3'd6) ? {{bias_add_162[31],bias_add_162[21:15]}} :'d6) : '0;
logic [7:0] relu_163;
assign relu_163[7:0] = (bias_add_163[31]==0) ? ((bias_add_163<3'd6) ? {{bias_add_163[31],bias_add_163[21:15]}} :'d6) : '0;
logic [7:0] relu_164;
assign relu_164[7:0] = (bias_add_164[31]==0) ? ((bias_add_164<3'd6) ? {{bias_add_164[31],bias_add_164[21:15]}} :'d6) : '0;
logic [7:0] relu_165;
assign relu_165[7:0] = (bias_add_165[31]==0) ? ((bias_add_165<3'd6) ? {{bias_add_165[31],bias_add_165[21:15]}} :'d6) : '0;
logic [7:0] relu_166;
assign relu_166[7:0] = (bias_add_166[31]==0) ? ((bias_add_166<3'd6) ? {{bias_add_166[31],bias_add_166[21:15]}} :'d6) : '0;
logic [7:0] relu_167;
assign relu_167[7:0] = (bias_add_167[31]==0) ? ((bias_add_167<3'd6) ? {{bias_add_167[31],bias_add_167[21:15]}} :'d6) : '0;
logic [7:0] relu_168;
assign relu_168[7:0] = (bias_add_168[31]==0) ? ((bias_add_168<3'd6) ? {{bias_add_168[31],bias_add_168[21:15]}} :'d6) : '0;
logic [7:0] relu_169;
assign relu_169[7:0] = (bias_add_169[31]==0) ? ((bias_add_169<3'd6) ? {{bias_add_169[31],bias_add_169[21:15]}} :'d6) : '0;
logic [7:0] relu_170;
assign relu_170[7:0] = (bias_add_170[31]==0) ? ((bias_add_170<3'd6) ? {{bias_add_170[31],bias_add_170[21:15]}} :'d6) : '0;
logic [7:0] relu_171;
assign relu_171[7:0] = (bias_add_171[31]==0) ? ((bias_add_171<3'd6) ? {{bias_add_171[31],bias_add_171[21:15]}} :'d6) : '0;
logic [7:0] relu_172;
assign relu_172[7:0] = (bias_add_172[31]==0) ? ((bias_add_172<3'd6) ? {{bias_add_172[31],bias_add_172[21:15]}} :'d6) : '0;
logic [7:0] relu_173;
assign relu_173[7:0] = (bias_add_173[31]==0) ? ((bias_add_173<3'd6) ? {{bias_add_173[31],bias_add_173[21:15]}} :'d6) : '0;
logic [7:0] relu_174;
assign relu_174[7:0] = (bias_add_174[31]==0) ? ((bias_add_174<3'd6) ? {{bias_add_174[31],bias_add_174[21:15]}} :'d6) : '0;
logic [7:0] relu_175;
assign relu_175[7:0] = (bias_add_175[31]==0) ? ((bias_add_175<3'd6) ? {{bias_add_175[31],bias_add_175[21:15]}} :'d6) : '0;
logic [7:0] relu_176;
assign relu_176[7:0] = (bias_add_176[31]==0) ? ((bias_add_176<3'd6) ? {{bias_add_176[31],bias_add_176[21:15]}} :'d6) : '0;
logic [7:0] relu_177;
assign relu_177[7:0] = (bias_add_177[31]==0) ? ((bias_add_177<3'd6) ? {{bias_add_177[31],bias_add_177[21:15]}} :'d6) : '0;
logic [7:0] relu_178;
assign relu_178[7:0] = (bias_add_178[31]==0) ? ((bias_add_178<3'd6) ? {{bias_add_178[31],bias_add_178[21:15]}} :'d6) : '0;
logic [7:0] relu_179;
assign relu_179[7:0] = (bias_add_179[31]==0) ? ((bias_add_179<3'd6) ? {{bias_add_179[31],bias_add_179[21:15]}} :'d6) : '0;
logic [7:0] relu_180;
assign relu_180[7:0] = (bias_add_180[31]==0) ? ((bias_add_180<3'd6) ? {{bias_add_180[31],bias_add_180[21:15]}} :'d6) : '0;
logic [7:0] relu_181;
assign relu_181[7:0] = (bias_add_181[31]==0) ? ((bias_add_181<3'd6) ? {{bias_add_181[31],bias_add_181[21:15]}} :'d6) : '0;
logic [7:0] relu_182;
assign relu_182[7:0] = (bias_add_182[31]==0) ? ((bias_add_182<3'd6) ? {{bias_add_182[31],bias_add_182[21:15]}} :'d6) : '0;
logic [7:0] relu_183;
assign relu_183[7:0] = (bias_add_183[31]==0) ? ((bias_add_183<3'd6) ? {{bias_add_183[31],bias_add_183[21:15]}} :'d6) : '0;
logic [7:0] relu_184;
assign relu_184[7:0] = (bias_add_184[31]==0) ? ((bias_add_184<3'd6) ? {{bias_add_184[31],bias_add_184[21:15]}} :'d6) : '0;
logic [7:0] relu_185;
assign relu_185[7:0] = (bias_add_185[31]==0) ? ((bias_add_185<3'd6) ? {{bias_add_185[31],bias_add_185[21:15]}} :'d6) : '0;
logic [7:0] relu_186;
assign relu_186[7:0] = (bias_add_186[31]==0) ? ((bias_add_186<3'd6) ? {{bias_add_186[31],bias_add_186[21:15]}} :'d6) : '0;
logic [7:0] relu_187;
assign relu_187[7:0] = (bias_add_187[31]==0) ? ((bias_add_187<3'd6) ? {{bias_add_187[31],bias_add_187[21:15]}} :'d6) : '0;
logic [7:0] relu_188;
assign relu_188[7:0] = (bias_add_188[31]==0) ? ((bias_add_188<3'd6) ? {{bias_add_188[31],bias_add_188[21:15]}} :'d6) : '0;
logic [7:0] relu_189;
assign relu_189[7:0] = (bias_add_189[31]==0) ? ((bias_add_189<3'd6) ? {{bias_add_189[31],bias_add_189[21:15]}} :'d6) : '0;
logic [7:0] relu_190;
assign relu_190[7:0] = (bias_add_190[31]==0) ? ((bias_add_190<3'd6) ? {{bias_add_190[31],bias_add_190[21:15]}} :'d6) : '0;
logic [7:0] relu_191;
assign relu_191[7:0] = (bias_add_191[31]==0) ? ((bias_add_191<3'd6) ? {{bias_add_191[31],bias_add_191[21:15]}} :'d6) : '0;
logic [7:0] relu_192;
assign relu_192[7:0] = (bias_add_192[31]==0) ? ((bias_add_192<3'd6) ? {{bias_add_192[31],bias_add_192[21:15]}} :'d6) : '0;
logic [7:0] relu_193;
assign relu_193[7:0] = (bias_add_193[31]==0) ? ((bias_add_193<3'd6) ? {{bias_add_193[31],bias_add_193[21:15]}} :'d6) : '0;
logic [7:0] relu_194;
assign relu_194[7:0] = (bias_add_194[31]==0) ? ((bias_add_194<3'd6) ? {{bias_add_194[31],bias_add_194[21:15]}} :'d6) : '0;
logic [7:0] relu_195;
assign relu_195[7:0] = (bias_add_195[31]==0) ? ((bias_add_195<3'd6) ? {{bias_add_195[31],bias_add_195[21:15]}} :'d6) : '0;
logic [7:0] relu_196;
assign relu_196[7:0] = (bias_add_196[31]==0) ? ((bias_add_196<3'd6) ? {{bias_add_196[31],bias_add_196[21:15]}} :'d6) : '0;
logic [7:0] relu_197;
assign relu_197[7:0] = (bias_add_197[31]==0) ? ((bias_add_197<3'd6) ? {{bias_add_197[31],bias_add_197[21:15]}} :'d6) : '0;
logic [7:0] relu_198;
assign relu_198[7:0] = (bias_add_198[31]==0) ? ((bias_add_198<3'd6) ? {{bias_add_198[31],bias_add_198[21:15]}} :'d6) : '0;
logic [7:0] relu_199;
assign relu_199[7:0] = (bias_add_199[31]==0) ? ((bias_add_199<3'd6) ? {{bias_add_199[31],bias_add_199[21:15]}} :'d6) : '0;
logic [7:0] relu_200;
assign relu_200[7:0] = (bias_add_200[31]==0) ? ((bias_add_200<3'd6) ? {{bias_add_200[31],bias_add_200[21:15]}} :'d6) : '0;
logic [7:0] relu_201;
assign relu_201[7:0] = (bias_add_201[31]==0) ? ((bias_add_201<3'd6) ? {{bias_add_201[31],bias_add_201[21:15]}} :'d6) : '0;
logic [7:0] relu_202;
assign relu_202[7:0] = (bias_add_202[31]==0) ? ((bias_add_202<3'd6) ? {{bias_add_202[31],bias_add_202[21:15]}} :'d6) : '0;
logic [7:0] relu_203;
assign relu_203[7:0] = (bias_add_203[31]==0) ? ((bias_add_203<3'd6) ? {{bias_add_203[31],bias_add_203[21:15]}} :'d6) : '0;
logic [7:0] relu_204;
assign relu_204[7:0] = (bias_add_204[31]==0) ? ((bias_add_204<3'd6) ? {{bias_add_204[31],bias_add_204[21:15]}} :'d6) : '0;
logic [7:0] relu_205;
assign relu_205[7:0] = (bias_add_205[31]==0) ? ((bias_add_205<3'd6) ? {{bias_add_205[31],bias_add_205[21:15]}} :'d6) : '0;
logic [7:0] relu_206;
assign relu_206[7:0] = (bias_add_206[31]==0) ? ((bias_add_206<3'd6) ? {{bias_add_206[31],bias_add_206[21:15]}} :'d6) : '0;
logic [7:0] relu_207;
assign relu_207[7:0] = (bias_add_207[31]==0) ? ((bias_add_207<3'd6) ? {{bias_add_207[31],bias_add_207[21:15]}} :'d6) : '0;
logic [7:0] relu_208;
assign relu_208[7:0] = (bias_add_208[31]==0) ? ((bias_add_208<3'd6) ? {{bias_add_208[31],bias_add_208[21:15]}} :'d6) : '0;
logic [7:0] relu_209;
assign relu_209[7:0] = (bias_add_209[31]==0) ? ((bias_add_209<3'd6) ? {{bias_add_209[31],bias_add_209[21:15]}} :'d6) : '0;
logic [7:0] relu_210;
assign relu_210[7:0] = (bias_add_210[31]==0) ? ((bias_add_210<3'd6) ? {{bias_add_210[31],bias_add_210[21:15]}} :'d6) : '0;
logic [7:0] relu_211;
assign relu_211[7:0] = (bias_add_211[31]==0) ? ((bias_add_211<3'd6) ? {{bias_add_211[31],bias_add_211[21:15]}} :'d6) : '0;
logic [7:0] relu_212;
assign relu_212[7:0] = (bias_add_212[31]==0) ? ((bias_add_212<3'd6) ? {{bias_add_212[31],bias_add_212[21:15]}} :'d6) : '0;
logic [7:0] relu_213;
assign relu_213[7:0] = (bias_add_213[31]==0) ? ((bias_add_213<3'd6) ? {{bias_add_213[31],bias_add_213[21:15]}} :'d6) : '0;
logic [7:0] relu_214;
assign relu_214[7:0] = (bias_add_214[31]==0) ? ((bias_add_214<3'd6) ? {{bias_add_214[31],bias_add_214[21:15]}} :'d6) : '0;
logic [7:0] relu_215;
assign relu_215[7:0] = (bias_add_215[31]==0) ? ((bias_add_215<3'd6) ? {{bias_add_215[31],bias_add_215[21:15]}} :'d6) : '0;
logic [7:0] relu_216;
assign relu_216[7:0] = (bias_add_216[31]==0) ? ((bias_add_216<3'd6) ? {{bias_add_216[31],bias_add_216[21:15]}} :'d6) : '0;
logic [7:0] relu_217;
assign relu_217[7:0] = (bias_add_217[31]==0) ? ((bias_add_217<3'd6) ? {{bias_add_217[31],bias_add_217[21:15]}} :'d6) : '0;
logic [7:0] relu_218;
assign relu_218[7:0] = (bias_add_218[31]==0) ? ((bias_add_218<3'd6) ? {{bias_add_218[31],bias_add_218[21:15]}} :'d6) : '0;
logic [7:0] relu_219;
assign relu_219[7:0] = (bias_add_219[31]==0) ? ((bias_add_219<3'd6) ? {{bias_add_219[31],bias_add_219[21:15]}} :'d6) : '0;
logic [7:0] relu_220;
assign relu_220[7:0] = (bias_add_220[31]==0) ? ((bias_add_220<3'd6) ? {{bias_add_220[31],bias_add_220[21:15]}} :'d6) : '0;
logic [7:0] relu_221;
assign relu_221[7:0] = (bias_add_221[31]==0) ? ((bias_add_221<3'd6) ? {{bias_add_221[31],bias_add_221[21:15]}} :'d6) : '0;
logic [7:0] relu_222;
assign relu_222[7:0] = (bias_add_222[31]==0) ? ((bias_add_222<3'd6) ? {{bias_add_222[31],bias_add_222[21:15]}} :'d6) : '0;
logic [7:0] relu_223;
assign relu_223[7:0] = (bias_add_223[31]==0) ? ((bias_add_223<3'd6) ? {{bias_add_223[31],bias_add_223[21:15]}} :'d6) : '0;
logic [7:0] relu_224;
assign relu_224[7:0] = (bias_add_224[31]==0) ? ((bias_add_224<3'd6) ? {{bias_add_224[31],bias_add_224[21:15]}} :'d6) : '0;
logic [7:0] relu_225;
assign relu_225[7:0] = (bias_add_225[31]==0) ? ((bias_add_225<3'd6) ? {{bias_add_225[31],bias_add_225[21:15]}} :'d6) : '0;
logic [7:0] relu_226;
assign relu_226[7:0] = (bias_add_226[31]==0) ? ((bias_add_226<3'd6) ? {{bias_add_226[31],bias_add_226[21:15]}} :'d6) : '0;
logic [7:0] relu_227;
assign relu_227[7:0] = (bias_add_227[31]==0) ? ((bias_add_227<3'd6) ? {{bias_add_227[31],bias_add_227[21:15]}} :'d6) : '0;
logic [7:0] relu_228;
assign relu_228[7:0] = (bias_add_228[31]==0) ? ((bias_add_228<3'd6) ? {{bias_add_228[31],bias_add_228[21:15]}} :'d6) : '0;
logic [7:0] relu_229;
assign relu_229[7:0] = (bias_add_229[31]==0) ? ((bias_add_229<3'd6) ? {{bias_add_229[31],bias_add_229[21:15]}} :'d6) : '0;
logic [7:0] relu_230;
assign relu_230[7:0] = (bias_add_230[31]==0) ? ((bias_add_230<3'd6) ? {{bias_add_230[31],bias_add_230[21:15]}} :'d6) : '0;
logic [7:0] relu_231;
assign relu_231[7:0] = (bias_add_231[31]==0) ? ((bias_add_231<3'd6) ? {{bias_add_231[31],bias_add_231[21:15]}} :'d6) : '0;
logic [7:0] relu_232;
assign relu_232[7:0] = (bias_add_232[31]==0) ? ((bias_add_232<3'd6) ? {{bias_add_232[31],bias_add_232[21:15]}} :'d6) : '0;
logic [7:0] relu_233;
assign relu_233[7:0] = (bias_add_233[31]==0) ? ((bias_add_233<3'd6) ? {{bias_add_233[31],bias_add_233[21:15]}} :'d6) : '0;
logic [7:0] relu_234;
assign relu_234[7:0] = (bias_add_234[31]==0) ? ((bias_add_234<3'd6) ? {{bias_add_234[31],bias_add_234[21:15]}} :'d6) : '0;
logic [7:0] relu_235;
assign relu_235[7:0] = (bias_add_235[31]==0) ? ((bias_add_235<3'd6) ? {{bias_add_235[31],bias_add_235[21:15]}} :'d6) : '0;
logic [7:0] relu_236;
assign relu_236[7:0] = (bias_add_236[31]==0) ? ((bias_add_236<3'd6) ? {{bias_add_236[31],bias_add_236[21:15]}} :'d6) : '0;
logic [7:0] relu_237;
assign relu_237[7:0] = (bias_add_237[31]==0) ? ((bias_add_237<3'd6) ? {{bias_add_237[31],bias_add_237[21:15]}} :'d6) : '0;
logic [7:0] relu_238;
assign relu_238[7:0] = (bias_add_238[31]==0) ? ((bias_add_238<3'd6) ? {{bias_add_238[31],bias_add_238[21:15]}} :'d6) : '0;
logic [7:0] relu_239;
assign relu_239[7:0] = (bias_add_239[31]==0) ? ((bias_add_239<3'd6) ? {{bias_add_239[31],bias_add_239[21:15]}} :'d6) : '0;
logic [7:0] relu_240;
assign relu_240[7:0] = (bias_add_240[31]==0) ? ((bias_add_240<3'd6) ? {{bias_add_240[31],bias_add_240[21:15]}} :'d6) : '0;
logic [7:0] relu_241;
assign relu_241[7:0] = (bias_add_241[31]==0) ? ((bias_add_241<3'd6) ? {{bias_add_241[31],bias_add_241[21:15]}} :'d6) : '0;
logic [7:0] relu_242;
assign relu_242[7:0] = (bias_add_242[31]==0) ? ((bias_add_242<3'd6) ? {{bias_add_242[31],bias_add_242[21:15]}} :'d6) : '0;
logic [7:0] relu_243;
assign relu_243[7:0] = (bias_add_243[31]==0) ? ((bias_add_243<3'd6) ? {{bias_add_243[31],bias_add_243[21:15]}} :'d6) : '0;
logic [7:0] relu_244;
assign relu_244[7:0] = (bias_add_244[31]==0) ? ((bias_add_244<3'd6) ? {{bias_add_244[31],bias_add_244[21:15]}} :'d6) : '0;
logic [7:0] relu_245;
assign relu_245[7:0] = (bias_add_245[31]==0) ? ((bias_add_245<3'd6) ? {{bias_add_245[31],bias_add_245[21:15]}} :'d6) : '0;
logic [7:0] relu_246;
assign relu_246[7:0] = (bias_add_246[31]==0) ? ((bias_add_246<3'd6) ? {{bias_add_246[31],bias_add_246[21:15]}} :'d6) : '0;
logic [7:0] relu_247;
assign relu_247[7:0] = (bias_add_247[31]==0) ? ((bias_add_247<3'd6) ? {{bias_add_247[31],bias_add_247[21:15]}} :'d6) : '0;
logic [7:0] relu_248;
assign relu_248[7:0] = (bias_add_248[31]==0) ? ((bias_add_248<3'd6) ? {{bias_add_248[31],bias_add_248[21:15]}} :'d6) : '0;
logic [7:0] relu_249;
assign relu_249[7:0] = (bias_add_249[31]==0) ? ((bias_add_249<3'd6) ? {{bias_add_249[31],bias_add_249[21:15]}} :'d6) : '0;
logic [7:0] relu_250;
assign relu_250[7:0] = (bias_add_250[31]==0) ? ((bias_add_250<3'd6) ? {{bias_add_250[31],bias_add_250[21:15]}} :'d6) : '0;
logic [7:0] relu_251;
assign relu_251[7:0] = (bias_add_251[31]==0) ? ((bias_add_251<3'd6) ? {{bias_add_251[31],bias_add_251[21:15]}} :'d6) : '0;
logic [7:0] relu_252;
assign relu_252[7:0] = (bias_add_252[31]==0) ? ((bias_add_252<3'd6) ? {{bias_add_252[31],bias_add_252[21:15]}} :'d6) : '0;
logic [7:0] relu_253;
assign relu_253[7:0] = (bias_add_253[31]==0) ? ((bias_add_253<3'd6) ? {{bias_add_253[31],bias_add_253[21:15]}} :'d6) : '0;
logic [7:0] relu_254;
assign relu_254[7:0] = (bias_add_254[31]==0) ? ((bias_add_254<3'd6) ? {{bias_add_254[31],bias_add_254[21:15]}} :'d6) : '0;
logic [7:0] relu_255;
assign relu_255[7:0] = (bias_add_255[31]==0) ? ((bias_add_255<3'd6) ? {{bias_add_255[31],bias_add_255[21:15]}} :'d6) : '0;

assign output_act = {
	relu_255,
	relu_254,
	relu_253,
	relu_252,
	relu_251,
	relu_250,
	relu_249,
	relu_248,
	relu_247,
	relu_246,
	relu_245,
	relu_244,
	relu_243,
	relu_242,
	relu_241,
	relu_240,
	relu_239,
	relu_238,
	relu_237,
	relu_236,
	relu_235,
	relu_234,
	relu_233,
	relu_232,
	relu_231,
	relu_230,
	relu_229,
	relu_228,
	relu_227,
	relu_226,
	relu_225,
	relu_224,
	relu_223,
	relu_222,
	relu_221,
	relu_220,
	relu_219,
	relu_218,
	relu_217,
	relu_216,
	relu_215,
	relu_214,
	relu_213,
	relu_212,
	relu_211,
	relu_210,
	relu_209,
	relu_208,
	relu_207,
	relu_206,
	relu_205,
	relu_204,
	relu_203,
	relu_202,
	relu_201,
	relu_200,
	relu_199,
	relu_198,
	relu_197,
	relu_196,
	relu_195,
	relu_194,
	relu_193,
	relu_192,
	relu_191,
	relu_190,
	relu_189,
	relu_188,
	relu_187,
	relu_186,
	relu_185,
	relu_184,
	relu_183,
	relu_182,
	relu_181,
	relu_180,
	relu_179,
	relu_178,
	relu_177,
	relu_176,
	relu_175,
	relu_174,
	relu_173,
	relu_172,
	relu_171,
	relu_170,
	relu_169,
	relu_168,
	relu_167,
	relu_166,
	relu_165,
	relu_164,
	relu_163,
	relu_162,
	relu_161,
	relu_160,
	relu_159,
	relu_158,
	relu_157,
	relu_156,
	relu_155,
	relu_154,
	relu_153,
	relu_152,
	relu_151,
	relu_150,
	relu_149,
	relu_148,
	relu_147,
	relu_146,
	relu_145,
	relu_144,
	relu_143,
	relu_142,
	relu_141,
	relu_140,
	relu_139,
	relu_138,
	relu_137,
	relu_136,
	relu_135,
	relu_134,
	relu_133,
	relu_132,
	relu_131,
	relu_130,
	relu_129,
	relu_128,
	relu_127,
	relu_126,
	relu_125,
	relu_124,
	relu_123,
	relu_122,
	relu_121,
	relu_120,
	relu_119,
	relu_118,
	relu_117,
	relu_116,
	relu_115,
	relu_114,
	relu_113,
	relu_112,
	relu_111,
	relu_110,
	relu_109,
	relu_108,
	relu_107,
	relu_106,
	relu_105,
	relu_104,
	relu_103,
	relu_102,
	relu_101,
	relu_100,
	relu_99,
	relu_98,
	relu_97,
	relu_96,
	relu_95,
	relu_94,
	relu_93,
	relu_92,
	relu_91,
	relu_90,
	relu_89,
	relu_88,
	relu_87,
	relu_86,
	relu_85,
	relu_84,
	relu_83,
	relu_82,
	relu_81,
	relu_80,
	relu_79,
	relu_78,
	relu_77,
	relu_76,
	relu_75,
	relu_74,
	relu_73,
	relu_72,
	relu_71,
	relu_70,
	relu_69,
	relu_68,
	relu_67,
	relu_66,
	relu_65,
	relu_64,
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
